		9225 => x"FF",
		9226 => x"FF",
		9227 => x"FF",
		9228 => x"FF",
		9229 => x"FF",
		9230 => x"FF",
		9231 => x"FF",
		9232 => x"FF",
		9233 => x"FF",
		9234 => x"FF",
		9235 => x"FF",
		9236 => x"FF",
		9237 => x"FF",
		9238 => x"FF",
		9239 => x"FF",
		9240 => x"FF",
		9241 => x"FF",
		9242 => x"FF",
		9243 => x"FF",
		9244 => x"FF",
		9245 => x"FF",
		9246 => x"FF",
		9247 => x"FF",
		9248 => x"FF",
		9249 => x"FF",
		9250 => x"FF",
		9251 => x"FF",
		9252 => x"FF",
		9253 => x"FF",
		9254 => x"FF",
		9255 => x"FF",
		9256 => x"FF",
		9257 => x"FF",
		9258 => x"FF",
		9259 => x"FF",
		9260 => x"FF",
		9261 => x"FF",
		9262 => x"FF",
		9263 => x"FF",
		9264 => x"FF",
		9265 => x"FF",
		9266 => x"FF",
		9267 => x"FF",
		9268 => x"FF",
		9269 => x"FF",
		9270 => x"FF",
		9271 => x"FF",
		9272 => x"FF",
		9273 => x"FF",
		9274 => x"FF",
		10249 => x"FF",
		10250 => x"FF",
		10251 => x"FF",
		10252 => x"FF",
		10253 => x"FF",
		10254 => x"FF",
		10255 => x"FF",
		10256 => x"FF",
		10257 => x"FF",
		10258 => x"FF",
		10259 => x"FF",
		10260 => x"FF",
		10261 => x"FF",
		10262 => x"FF",
		10263 => x"FF",
		10264 => x"FF",
		10265 => x"FF",
		10266 => x"FF",
		10267 => x"FF",
		10268 => x"FF",
		10269 => x"FF",
		10270 => x"FF",
		10271 => x"FF",
		10272 => x"FF",
		10273 => x"FF",
		10274 => x"FF",
		10275 => x"FF",
		10276 => x"FF",
		10277 => x"FF",
		10278 => x"FF",
		10279 => x"FF",
		10280 => x"FF",
		10281 => x"FF",
		10282 => x"FF",
		10283 => x"FF",
		10284 => x"FF",
		10285 => x"FF",
		10286 => x"FF",
		10287 => x"FF",
		10288 => x"FF",
		10289 => x"FF",
		10290 => x"FF",
		10291 => x"FF",
		10292 => x"FF",
		10293 => x"FF",
		10294 => x"FF",
		10295 => x"FF",
		10296 => x"FF",
		10297 => x"FF",
		10298 => x"FF",
		11273 => x"FF",
		11274 => x"FF",
		11275 => x"FF",
		11276 => x"FF",
		11277 => x"FF",
		11278 => x"FF",
		11279 => x"FF",
		11280 => x"FF",
		11281 => x"FF",
		11282 => x"FF",
		11283 => x"FF",
		11284 => x"FF",
		11285 => x"FF",
		11286 => x"FF",
		11287 => x"FF",
		11288 => x"FF",
		11289 => x"FF",
		11290 => x"FF",
		11291 => x"FF",
		11292 => x"FF",
		11293 => x"FF",
		11294 => x"FF",
		11295 => x"FF",
		11296 => x"FF",
		11297 => x"FF",
		11298 => x"FF",
		11299 => x"FF",
		11300 => x"FF",
		11301 => x"FF",
		11302 => x"FF",
		11303 => x"FF",
		11304 => x"FF",
		11305 => x"FF",
		11306 => x"FF",
		11307 => x"FF",
		11308 => x"FF",
		11309 => x"FF",
		11310 => x"FF",
		11311 => x"FF",
		11312 => x"FF",
		11313 => x"FF",
		11314 => x"FF",
		11315 => x"FF",
		11316 => x"FF",
		11317 => x"FF",
		11318 => x"FF",
		11319 => x"FF",
		11320 => x"FF",
		11321 => x"FF",
		11322 => x"FF",
		12297 => x"FF",
		12298 => x"FF",
		12299 => x"FF",
		12300 => x"FF",
		12301 => x"FF",
		12302 => x"FF",
		12303 => x"FF",
		12304 => x"FF",
		12305 => x"FF",
		12306 => x"FF",
		12307 => x"FF",
		12308 => x"FF",
		12309 => x"FF",
		12310 => x"FF",
		12311 => x"FF",
		12312 => x"FF",
		12313 => x"FF",
		12314 => x"FF",
		12315 => x"FF",
		12316 => x"FF",
		12317 => x"FF",
		12318 => x"FF",
		12319 => x"FF",
		12320 => x"FF",
		12321 => x"FF",
		12322 => x"FF",
		12323 => x"FF",
		12324 => x"FF",
		12325 => x"FF",
		12326 => x"FF",
		12327 => x"FF",
		12328 => x"FF",
		12329 => x"FF",
		12330 => x"FF",
		12331 => x"FF",
		12332 => x"FF",
		12333 => x"FF",
		12334 => x"FF",
		12335 => x"FF",
		12336 => x"FF",
		12337 => x"FF",
		12338 => x"FF",
		12339 => x"FF",
		12340 => x"FF",
		12341 => x"FF",
		12342 => x"FF",
		12343 => x"FF",
		12344 => x"FF",
		12345 => x"FF",
		12346 => x"FF",
		13321 => x"FF",
		13322 => x"FF",
		13323 => x"FF",
		13324 => x"FF",
		13325 => x"FF",
		13326 => x"FF",
		13327 => x"FF",
		13328 => x"FF",
		13329 => x"FF",
		13330 => x"FF",
		13331 => x"FF",
		13332 => x"FF",
		13333 => x"FF",
		13334 => x"FF",
		13335 => x"FF",
		13336 => x"FF",
		13337 => x"FF",
		13338 => x"FF",
		13339 => x"FF",
		13340 => x"FF",
		13341 => x"FF",
		13342 => x"FF",
		13343 => x"FF",
		13344 => x"FF",
		13345 => x"FF",
		13346 => x"FF",
		13347 => x"FF",
		13348 => x"FF",
		13349 => x"FF",
		13350 => x"FF",
		13351 => x"FF",
		13352 => x"FF",
		13353 => x"FF",
		13354 => x"FF",
		13355 => x"FF",
		13356 => x"FF",
		13357 => x"FF",
		13358 => x"FF",
		13359 => x"FF",
		13360 => x"FF",
		13361 => x"FF",
		13362 => x"FF",
		13363 => x"FF",
		13364 => x"FF",
		13365 => x"FF",
		13366 => x"FF",
		13367 => x"FF",
		13368 => x"FF",
		13369 => x"FF",
		13370 => x"FF",
		14345 => x"FF",
		14346 => x"FF",
		14347 => x"FF",
		14348 => x"FF",
		14349 => x"FF",
		14360 => x"FF",
		14361 => x"FF",
		14362 => x"FF",
		14363 => x"FF",
		14364 => x"FF",
		14375 => x"FF",
		14376 => x"FF",
		14377 => x"FF",
		14378 => x"FF",
		14379 => x"FF",
		14390 => x"FF",
		14391 => x"FF",
		14392 => x"FF",
		14393 => x"FF",
		14394 => x"FF",
		15369 => x"FF",
		15370 => x"FF",
		15371 => x"FF",
		15372 => x"FF",
		15373 => x"FF",
		15384 => x"FF",
		15385 => x"FF",
		15386 => x"FF",
		15387 => x"FF",
		15388 => x"FF",
		15399 => x"FF",
		15400 => x"FF",
		15401 => x"FF",
		15402 => x"FF",
		15403 => x"FF",
		15414 => x"FF",
		15415 => x"FF",
		15416 => x"FF",
		15417 => x"FF",
		15418 => x"FF",
		16393 => x"FF",
		16394 => x"FF",
		16395 => x"FF",
		16396 => x"FF",
		16397 => x"FF",
		16408 => x"FF",
		16409 => x"FF",
		16410 => x"FF",
		16411 => x"FF",
		16412 => x"FF",
		16423 => x"FF",
		16424 => x"FF",
		16425 => x"FF",
		16426 => x"FF",
		16427 => x"FF",
		16438 => x"FF",
		16439 => x"FF",
		16440 => x"FF",
		16441 => x"FF",
		16442 => x"FF",
		17417 => x"FF",
		17418 => x"FF",
		17419 => x"FF",
		17420 => x"FF",
		17421 => x"FF",
		17432 => x"FF",
		17433 => x"FF",
		17434 => x"FF",
		17435 => x"FF",
		17436 => x"FF",
		17447 => x"FF",
		17448 => x"FF",
		17449 => x"FF",
		17450 => x"FF",
		17451 => x"FF",
		17462 => x"FF",
		17463 => x"FF",
		17464 => x"FF",
		17465 => x"FF",
		17466 => x"FF",
		18441 => x"FF",
		18442 => x"FF",
		18443 => x"FF",
		18444 => x"FF",
		18445 => x"FF",
		18456 => x"FF",
		18457 => x"FF",
		18458 => x"FF",
		18459 => x"FF",
		18460 => x"FF",
		18471 => x"FF",
		18472 => x"FF",
		18473 => x"FF",
		18474 => x"FF",
		18475 => x"FF",
		18486 => x"FF",
		18487 => x"FF",
		18488 => x"FF",
		18489 => x"FF",
		18490 => x"FF",
		19465 => x"FF",
		19466 => x"FF",
		19467 => x"FF",
		19468 => x"FF",
		19469 => x"FF",
		19480 => x"FF",
		19481 => x"FF",
		19482 => x"FF",
		19483 => x"FF",
		19484 => x"FF",
		19495 => x"FF",
		19496 => x"FF",
		19497 => x"FF",
		19498 => x"FF",
		19499 => x"FF",
		19510 => x"FF",
		19511 => x"FF",
		19512 => x"FF",
		19513 => x"FF",
		19514 => x"FF",
		20489 => x"FF",
		20490 => x"FF",
		20491 => x"FF",
		20492 => x"FF",
		20493 => x"FF",
		20504 => x"FF",
		20505 => x"FF",
		20506 => x"FF",
		20507 => x"FF",
		20508 => x"FF",
		20519 => x"FF",
		20520 => x"FF",
		20521 => x"FF",
		20522 => x"FF",
		20523 => x"FF",
		20534 => x"FF",
		20535 => x"FF",
		20536 => x"FF",
		20537 => x"FF",
		20538 => x"FF",
		21513 => x"FF",
		21514 => x"FF",
		21515 => x"FF",
		21516 => x"FF",
		21517 => x"FF",
		21528 => x"FF",
		21529 => x"FF",
		21530 => x"FF",
		21531 => x"FF",
		21532 => x"FF",
		21543 => x"FF",
		21544 => x"FF",
		21545 => x"FF",
		21546 => x"FF",
		21547 => x"FF",
		21558 => x"FF",
		21559 => x"FF",
		21560 => x"FF",
		21561 => x"FF",
		21562 => x"FF",
		22537 => x"FF",
		22538 => x"FF",
		22539 => x"FF",
		22540 => x"FF",
		22541 => x"FF",
		22552 => x"FF",
		22553 => x"FF",
		22554 => x"FF",
		22555 => x"FF",
		22556 => x"FF",
		22567 => x"FF",
		22568 => x"FF",
		22569 => x"FF",
		22570 => x"FF",
		22571 => x"FF",
		22582 => x"FF",
		22583 => x"FF",
		22584 => x"FF",
		22585 => x"FF",
		22586 => x"FF",
		23561 => x"FF",
		23562 => x"FF",
		23563 => x"FF",
		23564 => x"FF",
		23565 => x"FF",
		23576 => x"FF",
		23577 => x"FF",
		23578 => x"FF",
		23579 => x"FF",
		23580 => x"FF",
		23591 => x"FF",
		23592 => x"FF",
		23593 => x"FF",
		23594 => x"FF",
		23595 => x"FF",
		23606 => x"FF",
		23607 => x"FF",
		23608 => x"FF",
		23609 => x"FF",
		23610 => x"FF",
		24585 => x"FF",
		24586 => x"FF",
		24587 => x"FF",
		24588 => x"FF",
		24589 => x"FF",
		24590 => x"FF",
		24591 => x"FF",
		24592 => x"FF",
		24593 => x"FF",
		24594 => x"FF",
		24595 => x"FF",
		24596 => x"FF",
		24597 => x"FF",
		24598 => x"FF",
		24599 => x"FF",
		24600 => x"FF",
		24601 => x"FF",
		24602 => x"FF",
		24603 => x"FF",
		24604 => x"FF",
		24605 => x"FF",
		24606 => x"FF",
		24607 => x"FF",
		24608 => x"FF",
		24609 => x"FF",
		24610 => x"FF",
		24611 => x"FF",
		24612 => x"FF",
		24613 => x"FF",
		24614 => x"FF",
		24615 => x"FF",
		24616 => x"FF",
		24617 => x"FF",
		24618 => x"FF",
		24619 => x"FF",
		24620 => x"FF",
		24621 => x"FF",
		24622 => x"FF",
		24623 => x"FF",
		24624 => x"FF",
		24625 => x"FF",
		24626 => x"FF",
		24627 => x"FF",
		24628 => x"FF",
		24629 => x"FF",
		24630 => x"FF",
		24631 => x"FF",
		24632 => x"FF",
		24633 => x"FF",
		24634 => x"FF",
		25609 => x"FF",
		25610 => x"FF",
		25611 => x"FF",
		25612 => x"FF",
		25613 => x"FF",
		25614 => x"FF",
		25615 => x"FF",
		25616 => x"FF",
		25617 => x"FF",
		25618 => x"FF",
		25619 => x"FF",
		25620 => x"FF",
		25621 => x"FF",
		25622 => x"FF",
		25623 => x"FF",
		25624 => x"FF",
		25625 => x"FF",
		25626 => x"FF",
		25627 => x"FF",
		25628 => x"FF",
		25629 => x"FF",
		25630 => x"FF",
		25631 => x"FF",
		25632 => x"FF",
		25633 => x"FF",
		25634 => x"FF",
		25635 => x"FF",
		25636 => x"FF",
		25637 => x"FF",
		25638 => x"FF",
		25639 => x"FF",
		25640 => x"FF",
		25641 => x"FF",
		25642 => x"FF",
		25643 => x"FF",
		25644 => x"FF",
		25645 => x"FF",
		25646 => x"FF",
		25647 => x"FF",
		25648 => x"FF",
		25649 => x"FF",
		25650 => x"FF",
		25651 => x"FF",
		25652 => x"FF",
		25653 => x"FF",
		25654 => x"FF",
		25655 => x"FF",
		25656 => x"FF",
		25657 => x"FF",
		25658 => x"FF",
		26633 => x"FF",
		26634 => x"FF",
		26635 => x"FF",
		26636 => x"FF",
		26637 => x"FF",
		26638 => x"FF",
		26639 => x"FF",
		26640 => x"FF",
		26641 => x"FF",
		26642 => x"FF",
		26643 => x"FF",
		26644 => x"FF",
		26645 => x"FF",
		26646 => x"FF",
		26647 => x"FF",
		26648 => x"FF",
		26649 => x"FF",
		26650 => x"FF",
		26651 => x"FF",
		26652 => x"FF",
		26653 => x"FF",
		26654 => x"FF",
		26655 => x"FF",
		26656 => x"FF",
		26657 => x"FF",
		26658 => x"FF",
		26659 => x"FF",
		26660 => x"FF",
		26661 => x"FF",
		26662 => x"FF",
		26663 => x"FF",
		26664 => x"FF",
		26665 => x"FF",
		26666 => x"FF",
		26667 => x"FF",
		26668 => x"FF",
		26669 => x"FF",
		26670 => x"FF",
		26671 => x"FF",
		26672 => x"FF",
		26673 => x"FF",
		26674 => x"FF",
		26675 => x"FF",
		26676 => x"FF",
		26677 => x"FF",
		26678 => x"FF",
		26679 => x"FF",
		26680 => x"FF",
		26681 => x"FF",
		26682 => x"FF",
		27657 => x"FF",
		27658 => x"FF",
		27659 => x"FF",
		27660 => x"FF",
		27661 => x"FF",
		27662 => x"FF",
		27663 => x"FF",
		27664 => x"FF",
		27665 => x"FF",
		27666 => x"FF",
		27667 => x"FF",
		27668 => x"FF",
		27669 => x"FF",
		27670 => x"FF",
		27671 => x"FF",
		27672 => x"FF",
		27673 => x"FF",
		27674 => x"FF",
		27675 => x"FF",
		27676 => x"FF",
		27677 => x"FF",
		27678 => x"FF",
		27679 => x"FF",
		27680 => x"FF",
		27681 => x"FF",
		27682 => x"FF",
		27683 => x"FF",
		27684 => x"FF",
		27685 => x"FF",
		27686 => x"FF",
		27687 => x"FF",
		27688 => x"FF",
		27689 => x"FF",
		27690 => x"FF",
		27691 => x"FF",
		27692 => x"FF",
		27693 => x"FF",
		27694 => x"FF",
		27695 => x"FF",
		27696 => x"FF",
		27697 => x"FF",
		27698 => x"FF",
		27699 => x"FF",
		27700 => x"FF",
		27701 => x"FF",
		27702 => x"FF",
		27703 => x"FF",
		27704 => x"FF",
		27705 => x"FF",
		27706 => x"FF",
		28681 => x"FF",
		28682 => x"FF",
		28683 => x"FF",
		28684 => x"FF",
		28685 => x"FF",
		28686 => x"FF",
		28687 => x"FF",
		28688 => x"FF",
		28689 => x"FF",
		28690 => x"FF",
		28691 => x"FF",
		28692 => x"FF",
		28693 => x"FF",
		28694 => x"FF",
		28695 => x"FF",
		28696 => x"FF",
		28697 => x"FF",
		28698 => x"FF",
		28699 => x"FF",
		28700 => x"FF",
		28701 => x"FF",
		28702 => x"FF",
		28703 => x"FF",
		28704 => x"FF",
		28705 => x"FF",
		28706 => x"FF",
		28707 => x"FF",
		28708 => x"FF",
		28709 => x"FF",
		28710 => x"FF",
		28711 => x"FF",
		28712 => x"FF",
		28713 => x"FF",
		28714 => x"FF",
		28715 => x"FF",
		28716 => x"FF",
		28717 => x"FF",
		28718 => x"FF",
		28719 => x"FF",
		28720 => x"FF",
		28721 => x"FF",
		28722 => x"FF",
		28723 => x"FF",
		28724 => x"FF",
		28725 => x"FF",
		28726 => x"FF",
		28727 => x"FF",
		28728 => x"FF",
		28729 => x"FF",
		28730 => x"FF",
		29705 => x"FF",
		29706 => x"FF",
		29707 => x"FF",
		29708 => x"FF",
		29709 => x"FF",
		29720 => x"FF",
		29721 => x"FF",
		29722 => x"FF",
		29723 => x"FF",
		29724 => x"FF",
		29735 => x"FF",
		29736 => x"FF",
		29737 => x"FF",
		29738 => x"FF",
		29739 => x"FF",
		29750 => x"FF",
		29751 => x"FF",
		29752 => x"FF",
		29753 => x"FF",
		29754 => x"FF",
		30729 => x"FF",
		30730 => x"FF",
		30731 => x"FF",
		30732 => x"FF",
		30733 => x"FF",
		30744 => x"FF",
		30745 => x"FF",
		30746 => x"FF",
		30747 => x"FF",
		30748 => x"FF",
		30759 => x"FF",
		30760 => x"FF",
		30761 => x"FF",
		30762 => x"FF",
		30763 => x"FF",
		30774 => x"FF",
		30775 => x"FF",
		30776 => x"FF",
		30777 => x"FF",
		30778 => x"FF",
		31753 => x"FF",
		31754 => x"FF",
		31755 => x"FF",
		31756 => x"FF",
		31757 => x"FF",
		31768 => x"FF",
		31769 => x"FF",
		31770 => x"FF",
		31771 => x"FF",
		31772 => x"FF",
		31783 => x"FF",
		31784 => x"FF",
		31785 => x"FF",
		31786 => x"FF",
		31787 => x"FF",
		31798 => x"FF",
		31799 => x"FF",
		31800 => x"FF",
		31801 => x"FF",
		31802 => x"FF",
		32777 => x"FF",
		32778 => x"FF",
		32779 => x"FF",
		32780 => x"FF",
		32781 => x"FF",
		32792 => x"FF",
		32793 => x"FF",
		32794 => x"FF",
		32795 => x"FF",
		32796 => x"FF",
		32807 => x"FF",
		32808 => x"FF",
		32809 => x"FF",
		32810 => x"FF",
		32811 => x"FF",
		32822 => x"FF",
		32823 => x"FF",
		32824 => x"FF",
		32825 => x"FF",
		32826 => x"FF",
		33801 => x"FF",
		33802 => x"FF",
		33803 => x"FF",
		33804 => x"FF",
		33805 => x"FF",
		33816 => x"FF",
		33817 => x"FF",
		33818 => x"FF",
		33819 => x"FF",
		33820 => x"FF",
		33831 => x"FF",
		33832 => x"FF",
		33833 => x"FF",
		33834 => x"FF",
		33835 => x"FF",
		33846 => x"FF",
		33847 => x"FF",
		33848 => x"FF",
		33849 => x"FF",
		33850 => x"FF",
		34825 => x"FF",
		34826 => x"FF",
		34827 => x"FF",
		34828 => x"FF",
		34829 => x"FF",
		34840 => x"FF",
		34841 => x"FF",
		34842 => x"FF",
		34843 => x"FF",
		34844 => x"FF",
		34855 => x"FF",
		34856 => x"FF",
		34857 => x"FF",
		34858 => x"FF",
		34859 => x"FF",
		34870 => x"FF",
		34871 => x"FF",
		34872 => x"FF",
		34873 => x"FF",
		34874 => x"FF",
		35849 => x"FF",
		35850 => x"FF",
		35851 => x"FF",
		35852 => x"FF",
		35853 => x"FF",
		35864 => x"FF",
		35865 => x"FF",
		35866 => x"FF",
		35867 => x"FF",
		35868 => x"FF",
		35879 => x"FF",
		35880 => x"FF",
		35881 => x"FF",
		35882 => x"FF",
		35883 => x"FF",
		35894 => x"FF",
		35895 => x"FF",
		35896 => x"FF",
		35897 => x"FF",
		35898 => x"FF",
		36873 => x"FF",
		36874 => x"FF",
		36875 => x"FF",
		36876 => x"FF",
		36877 => x"FF",
		36888 => x"FF",
		36889 => x"FF",
		36890 => x"FF",
		36891 => x"FF",
		36892 => x"FF",
		36903 => x"FF",
		36904 => x"FF",
		36905 => x"FF",
		36906 => x"FF",
		36907 => x"FF",
		36918 => x"FF",
		36919 => x"FF",
		36920 => x"FF",
		36921 => x"FF",
		36922 => x"FF",
		37897 => x"FF",
		37898 => x"FF",
		37899 => x"FF",
		37900 => x"FF",
		37901 => x"FF",
		37912 => x"FF",
		37913 => x"FF",
		37914 => x"FF",
		37915 => x"FF",
		37916 => x"FF",
		37927 => x"FF",
		37928 => x"FF",
		37929 => x"FF",
		37930 => x"FF",
		37931 => x"FF",
		37942 => x"FF",
		37943 => x"FF",
		37944 => x"FF",
		37945 => x"FF",
		37946 => x"FF",
		38921 => x"FF",
		38922 => x"FF",
		38923 => x"FF",
		38924 => x"FF",
		38925 => x"FF",
		38936 => x"FF",
		38937 => x"FF",
		38938 => x"FF",
		38939 => x"FF",
		38940 => x"FF",
		38951 => x"FF",
		38952 => x"FF",
		38953 => x"FF",
		38954 => x"FF",
		38955 => x"FF",
		38966 => x"FF",
		38967 => x"FF",
		38968 => x"FF",
		38969 => x"FF",
		38970 => x"FF",
		39945 => x"FF",
		39946 => x"FF",
		39947 => x"FF",
		39948 => x"FF",
		39949 => x"FF",
		39950 => x"FF",
		39951 => x"FF",
		39952 => x"FF",
		39953 => x"FF",
		39954 => x"FF",
		39955 => x"FF",
		39956 => x"FF",
		39957 => x"FF",
		39958 => x"FF",
		39959 => x"FF",
		39960 => x"FF",
		39961 => x"FF",
		39962 => x"FF",
		39963 => x"FF",
		39964 => x"FF",
		39965 => x"FF",
		39966 => x"FF",
		39967 => x"FF",
		39968 => x"FF",
		39969 => x"FF",
		39970 => x"FF",
		39971 => x"FF",
		39972 => x"FF",
		39973 => x"FF",
		39974 => x"FF",
		39975 => x"FF",
		39976 => x"FF",
		39977 => x"FF",
		39978 => x"FF",
		39979 => x"FF",
		39980 => x"FF",
		39981 => x"FF",
		39982 => x"FF",
		39983 => x"FF",
		39984 => x"FF",
		39985 => x"FF",
		39986 => x"FF",
		39987 => x"FF",
		39988 => x"FF",
		39989 => x"FF",
		39990 => x"FF",
		39991 => x"FF",
		39992 => x"FF",
		39993 => x"FF",
		39994 => x"FF",
		40969 => x"FF",
		40970 => x"FF",
		40971 => x"FF",
		40972 => x"FF",
		40973 => x"FF",
		40974 => x"FF",
		40975 => x"FF",
		40976 => x"FF",
		40977 => x"FF",
		40978 => x"FF",
		40979 => x"FF",
		40980 => x"FF",
		40981 => x"FF",
		40982 => x"FF",
		40983 => x"FF",
		40984 => x"FF",
		40985 => x"FF",
		40986 => x"FF",
		40987 => x"FF",
		40988 => x"FF",
		40989 => x"FF",
		40990 => x"FF",
		40991 => x"FF",
		40992 => x"FF",
		40993 => x"FF",
		40994 => x"FF",
		40995 => x"FF",
		40996 => x"FF",
		40997 => x"FF",
		40998 => x"FF",
		40999 => x"FF",
		41000 => x"FF",
		41001 => x"FF",
		41002 => x"FF",
		41003 => x"FF",
		41004 => x"FF",
		41005 => x"FF",
		41006 => x"FF",
		41007 => x"FF",
		41008 => x"FF",
		41009 => x"FF",
		41010 => x"FF",
		41011 => x"FF",
		41012 => x"FF",
		41013 => x"FF",
		41014 => x"FF",
		41015 => x"FF",
		41016 => x"FF",
		41017 => x"FF",
		41018 => x"FF",
		41993 => x"FF",
		41994 => x"FF",
		41995 => x"FF",
		41996 => x"FF",
		41997 => x"FF",
		41998 => x"FF",
		41999 => x"FF",
		42000 => x"FF",
		42001 => x"FF",
		42002 => x"FF",
		42003 => x"FF",
		42004 => x"FF",
		42005 => x"FF",
		42006 => x"FF",
		42007 => x"FF",
		42008 => x"FF",
		42009 => x"FF",
		42010 => x"FF",
		42011 => x"FF",
		42012 => x"FF",
		42013 => x"FF",
		42014 => x"FF",
		42015 => x"FF",
		42016 => x"FF",
		42017 => x"FF",
		42018 => x"FF",
		42019 => x"FF",
		42020 => x"FF",
		42021 => x"FF",
		42022 => x"FF",
		42023 => x"FF",
		42024 => x"FF",
		42025 => x"FF",
		42026 => x"FF",
		42027 => x"FF",
		42028 => x"FF",
		42029 => x"FF",
		42030 => x"FF",
		42031 => x"FF",
		42032 => x"FF",
		42033 => x"FF",
		42034 => x"FF",
		42035 => x"FF",
		42036 => x"FF",
		42037 => x"FF",
		42038 => x"FF",
		42039 => x"FF",
		42040 => x"FF",
		42041 => x"FF",
		42042 => x"FF",
		43017 => x"FF",
		43018 => x"FF",
		43019 => x"FF",
		43020 => x"FF",
		43021 => x"FF",
		43022 => x"FF",
		43023 => x"FF",
		43024 => x"FF",
		43025 => x"FF",
		43026 => x"FF",
		43027 => x"FF",
		43028 => x"FF",
		43029 => x"FF",
		43030 => x"FF",
		43031 => x"FF",
		43032 => x"FF",
		43033 => x"FF",
		43034 => x"FF",
		43035 => x"FF",
		43036 => x"FF",
		43037 => x"FF",
		43038 => x"FF",
		43039 => x"FF",
		43040 => x"FF",
		43041 => x"FF",
		43042 => x"FF",
		43043 => x"FF",
		43044 => x"FF",
		43045 => x"FF",
		43046 => x"FF",
		43047 => x"FF",
		43048 => x"FF",
		43049 => x"FF",
		43050 => x"FF",
		43051 => x"FF",
		43052 => x"FF",
		43053 => x"FF",
		43054 => x"FF",
		43055 => x"FF",
		43056 => x"FF",
		43057 => x"FF",
		43058 => x"FF",
		43059 => x"FF",
		43060 => x"FF",
		43061 => x"FF",
		43062 => x"FF",
		43063 => x"FF",
		43064 => x"FF",
		43065 => x"FF",
		43066 => x"FF",
		44041 => x"FF",
		44042 => x"FF",
		44043 => x"FF",
		44044 => x"FF",
		44045 => x"FF",
		44046 => x"FF",
		44047 => x"FF",
		44048 => x"FF",
		44049 => x"FF",
		44050 => x"FF",
		44051 => x"FF",
		44052 => x"FF",
		44053 => x"FF",
		44054 => x"FF",
		44055 => x"FF",
		44056 => x"FF",
		44057 => x"FF",
		44058 => x"FF",
		44059 => x"FF",
		44060 => x"FF",
		44061 => x"FF",
		44062 => x"FF",
		44063 => x"FF",
		44064 => x"FF",
		44065 => x"FF",
		44066 => x"FF",
		44067 => x"FF",
		44068 => x"FF",
		44069 => x"FF",
		44070 => x"FF",
		44071 => x"FF",
		44072 => x"FF",
		44073 => x"FF",
		44074 => x"FF",
		44075 => x"FF",
		44076 => x"FF",
		44077 => x"FF",
		44078 => x"FF",
		44079 => x"FF",
		44080 => x"FF",
		44081 => x"FF",
		44082 => x"FF",
		44083 => x"FF",
		44084 => x"FF",
		44085 => x"FF",
		44086 => x"FF",
		44087 => x"FF",
		44088 => x"FF",
		44089 => x"FF",
		44090 => x"FF",
		45065 => x"FF",
		45066 => x"FF",
		45067 => x"FF",
		45068 => x"FF",
		45069 => x"FF",
		45080 => x"FF",
		45081 => x"FF",
		45082 => x"FF",
		45083 => x"FF",
		45084 => x"FF",
		45095 => x"FF",
		45096 => x"FF",
		45097 => x"FF",
		45098 => x"FF",
		45099 => x"FF",
		45110 => x"FF",
		45111 => x"FF",
		45112 => x"FF",
		45113 => x"FF",
		45114 => x"FF",
		46089 => x"FF",
		46090 => x"FF",
		46091 => x"FF",
		46092 => x"FF",
		46093 => x"FF",
		46104 => x"FF",
		46105 => x"FF",
		46106 => x"FF",
		46107 => x"FF",
		46108 => x"FF",
		46119 => x"FF",
		46120 => x"FF",
		46121 => x"FF",
		46122 => x"FF",
		46123 => x"FF",
		46134 => x"FF",
		46135 => x"FF",
		46136 => x"FF",
		46137 => x"FF",
		46138 => x"FF",
		47113 => x"FF",
		47114 => x"FF",
		47115 => x"FF",
		47116 => x"FF",
		47117 => x"FF",
		47128 => x"FF",
		47129 => x"FF",
		47130 => x"FF",
		47131 => x"FF",
		47132 => x"FF",
		47143 => x"FF",
		47144 => x"FF",
		47145 => x"FF",
		47146 => x"FF",
		47147 => x"FF",
		47158 => x"FF",
		47159 => x"FF",
		47160 => x"FF",
		47161 => x"FF",
		47162 => x"FF",
		48137 => x"FF",
		48138 => x"FF",
		48139 => x"FF",
		48140 => x"FF",
		48141 => x"FF",
		48152 => x"FF",
		48153 => x"FF",
		48154 => x"FF",
		48155 => x"FF",
		48156 => x"FF",
		48167 => x"FF",
		48168 => x"FF",
		48169 => x"FF",
		48170 => x"FF",
		48171 => x"FF",
		48182 => x"FF",
		48183 => x"FF",
		48184 => x"FF",
		48185 => x"FF",
		48186 => x"FF",
		49161 => x"FF",
		49162 => x"FF",
		49163 => x"FF",
		49164 => x"FF",
		49165 => x"FF",
		49176 => x"FF",
		49177 => x"FF",
		49178 => x"FF",
		49179 => x"FF",
		49180 => x"FF",
		49191 => x"FF",
		49192 => x"FF",
		49193 => x"FF",
		49194 => x"FF",
		49195 => x"FF",
		49206 => x"FF",
		49207 => x"FF",
		49208 => x"FF",
		49209 => x"FF",
		49210 => x"FF",
		50185 => x"FF",
		50186 => x"FF",
		50187 => x"FF",
		50188 => x"FF",
		50189 => x"FF",
		50200 => x"FF",
		50201 => x"FF",
		50202 => x"FF",
		50203 => x"FF",
		50204 => x"FF",
		50215 => x"FF",
		50216 => x"FF",
		50217 => x"FF",
		50218 => x"FF",
		50219 => x"FF",
		50230 => x"FF",
		50231 => x"FF",
		50232 => x"FF",
		50233 => x"FF",
		50234 => x"FF",
		51209 => x"FF",
		51210 => x"FF",
		51211 => x"FF",
		51212 => x"FF",
		51213 => x"FF",
		51224 => x"FF",
		51225 => x"FF",
		51226 => x"FF",
		51227 => x"FF",
		51228 => x"FF",
		51239 => x"FF",
		51240 => x"FF",
		51241 => x"FF",
		51242 => x"FF",
		51243 => x"FF",
		51254 => x"FF",
		51255 => x"FF",
		51256 => x"FF",
		51257 => x"FF",
		51258 => x"FF",
		52233 => x"FF",
		52234 => x"FF",
		52235 => x"FF",
		52236 => x"FF",
		52237 => x"FF",
		52248 => x"FF",
		52249 => x"FF",
		52250 => x"FF",
		52251 => x"FF",
		52252 => x"FF",
		52263 => x"FF",
		52264 => x"FF",
		52265 => x"FF",
		52266 => x"FF",
		52267 => x"FF",
		52278 => x"FF",
		52279 => x"FF",
		52280 => x"FF",
		52281 => x"FF",
		52282 => x"FF",
		53257 => x"FF",
		53258 => x"FF",
		53259 => x"FF",
		53260 => x"FF",
		53261 => x"FF",
		53272 => x"FF",
		53273 => x"FF",
		53274 => x"FF",
		53275 => x"FF",
		53276 => x"FF",
		53287 => x"FF",
		53288 => x"FF",
		53289 => x"FF",
		53290 => x"FF",
		53291 => x"FF",
		53302 => x"FF",
		53303 => x"FF",
		53304 => x"FF",
		53305 => x"FF",
		53306 => x"FF",
		54281 => x"FF",
		54282 => x"FF",
		54283 => x"FF",
		54284 => x"FF",
		54285 => x"FF",
		54296 => x"FF",
		54297 => x"FF",
		54298 => x"FF",
		54299 => x"FF",
		54300 => x"FF",
		54311 => x"FF",
		54312 => x"FF",
		54313 => x"FF",
		54314 => x"FF",
		54315 => x"FF",
		54326 => x"FF",
		54327 => x"FF",
		54328 => x"FF",
		54329 => x"FF",
		54330 => x"FF",
		55305 => x"FF",
		55306 => x"FF",
		55307 => x"FF",
		55308 => x"FF",
		55309 => x"FF",
		55310 => x"FF",
		55311 => x"FF",
		55312 => x"FF",
		55313 => x"FF",
		55314 => x"FF",
		55315 => x"FF",
		55316 => x"FF",
		55317 => x"FF",
		55318 => x"FF",
		55319 => x"FF",
		55320 => x"FF",
		55321 => x"FF",
		55322 => x"FF",
		55323 => x"FF",
		55324 => x"FF",
		55325 => x"FF",
		55326 => x"FF",
		55327 => x"FF",
		55328 => x"FF",
		55329 => x"FF",
		55330 => x"FF",
		55331 => x"FF",
		55332 => x"FF",
		55333 => x"FF",
		55334 => x"FF",
		55335 => x"FF",
		55336 => x"FF",
		55337 => x"FF",
		55338 => x"FF",
		55339 => x"FF",
		55340 => x"FF",
		55341 => x"FF",
		55342 => x"FF",
		55343 => x"FF",
		55344 => x"FF",
		55345 => x"FF",
		55346 => x"FF",
		55347 => x"FF",
		55348 => x"FF",
		55349 => x"FF",
		55350 => x"FF",
		55351 => x"FF",
		55352 => x"FF",
		55353 => x"FF",
		55354 => x"FF",
		56329 => x"FF",
		56330 => x"FF",
		56331 => x"FF",
		56332 => x"FF",
		56333 => x"FF",
		56334 => x"FF",
		56335 => x"FF",
		56336 => x"FF",
		56337 => x"FF",
		56338 => x"FF",
		56339 => x"FF",
		56340 => x"FF",
		56341 => x"FF",
		56342 => x"FF",
		56343 => x"FF",
		56344 => x"FF",
		56345 => x"FF",
		56346 => x"FF",
		56347 => x"FF",
		56348 => x"FF",
		56349 => x"FF",
		56350 => x"FF",
		56351 => x"FF",
		56352 => x"FF",
		56353 => x"FF",
		56354 => x"FF",
		56355 => x"FF",
		56356 => x"FF",
		56357 => x"FF",
		56358 => x"FF",
		56359 => x"FF",
		56360 => x"FF",
		56361 => x"FF",
		56362 => x"FF",
		56363 => x"FF",
		56364 => x"FF",
		56365 => x"FF",
		56366 => x"FF",
		56367 => x"FF",
		56368 => x"FF",
		56369 => x"FF",
		56370 => x"FF",
		56371 => x"FF",
		56372 => x"FF",
		56373 => x"FF",
		56374 => x"FF",
		56375 => x"FF",
		56376 => x"FF",
		56377 => x"FF",
		56378 => x"FF",
		57353 => x"FF",
		57354 => x"FF",
		57355 => x"FF",
		57356 => x"FF",
		57357 => x"FF",
		57358 => x"FF",
		57359 => x"FF",
		57360 => x"FF",
		57361 => x"FF",
		57362 => x"FF",
		57363 => x"FF",
		57364 => x"FF",
		57365 => x"FF",
		57366 => x"FF",
		57367 => x"FF",
		57368 => x"FF",
		57369 => x"FF",
		57370 => x"FF",
		57371 => x"FF",
		57372 => x"FF",
		57373 => x"FF",
		57374 => x"FF",
		57375 => x"FF",
		57376 => x"FF",
		57377 => x"FF",
		57378 => x"FF",
		57379 => x"FF",
		57380 => x"FF",
		57381 => x"FF",
		57382 => x"FF",
		57383 => x"FF",
		57384 => x"FF",
		57385 => x"FF",
		57386 => x"FF",
		57387 => x"FF",
		57388 => x"FF",
		57389 => x"FF",
		57390 => x"FF",
		57391 => x"FF",
		57392 => x"FF",
		57393 => x"FF",
		57394 => x"FF",
		57395 => x"FF",
		57396 => x"FF",
		57397 => x"FF",
		57398 => x"FF",
		57399 => x"FF",
		57400 => x"FF",
		57401 => x"FF",
		57402 => x"FF",
		58377 => x"FF",
		58378 => x"FF",
		58379 => x"FF",
		58380 => x"FF",
		58381 => x"FF",
		58382 => x"FF",
		58383 => x"FF",
		58384 => x"FF",
		58385 => x"FF",
		58386 => x"FF",
		58387 => x"FF",
		58388 => x"FF",
		58389 => x"FF",
		58390 => x"FF",
		58391 => x"FF",
		58392 => x"FF",
		58393 => x"FF",
		58394 => x"FF",
		58395 => x"FF",
		58396 => x"FF",
		58397 => x"FF",
		58398 => x"FF",
		58399 => x"FF",
		58400 => x"FF",
		58401 => x"FF",
		58402 => x"FF",
		58403 => x"FF",
		58404 => x"FF",
		58405 => x"FF",
		58406 => x"FF",
		58407 => x"FF",
		58408 => x"FF",
		58409 => x"FF",
		58410 => x"FF",
		58411 => x"FF",
		58412 => x"FF",
		58413 => x"FF",
		58414 => x"FF",
		58415 => x"FF",
		58416 => x"FF",
		58417 => x"FF",
		58418 => x"FF",
		58419 => x"FF",
		58420 => x"FF",
		58421 => x"FF",
		58422 => x"FF",
		58423 => x"FF",
		58424 => x"FF",
		58425 => x"FF",
		58426 => x"FF",
		59401 => x"FF",
		59402 => x"FF",
		59403 => x"FF",
		59404 => x"FF",
		59405 => x"FF",
		59406 => x"FF",
		59407 => x"FF",
		59408 => x"FF",
		59409 => x"FF",
		59410 => x"FF",
		59411 => x"FF",
		59412 => x"FF",
		59413 => x"FF",
		59414 => x"FF",
		59415 => x"FF",
		59416 => x"FF",
		59417 => x"FF",
		59418 => x"FF",
		59419 => x"FF",
		59420 => x"FF",
		59421 => x"FF",
		59422 => x"FF",
		59423 => x"FF",
		59424 => x"FF",
		59425 => x"FF",
		59426 => x"FF",
		59427 => x"FF",
		59428 => x"FF",
		59429 => x"FF",
		59430 => x"FF",
		59431 => x"FF",
		59432 => x"FF",
		59433 => x"FF",
		59434 => x"FF",
		59435 => x"FF",
		59436 => x"FF",
		59437 => x"FF",
		59438 => x"FF",
		59439 => x"FF",
		59440 => x"FF",
		59441 => x"FF",
		59442 => x"FF",
		59443 => x"FF",
		59444 => x"FF",
		59445 => x"FF",
		59446 => x"FF",
		59447 => x"FF",
		59448 => x"FF",
		59449 => x"FF",
		59450 => x"FF",
