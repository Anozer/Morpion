		6939 to 7130 => "11111111",
		7195 to 7386 => "11111111",
		7451 to 7642 => "11111111",
		7707 to 7709 => "11111111",
		7770 to 7772 => "11111111",
		7833 to 7835 => "11111111",
		7896 to 7898 => "11111111",
		7963 to 7965 => "11111111",
		8026 to 8028 => "11111111",
		8089 to 8091 => "11111111",
		8152 to 8154 => "11111111",
		8219 to 8221 => "11111111",
		8282 to 8284 => "11111111",
		8345 to 8347 => "11111111",
		8408 to 8410 => "11111111",
		8475 to 8477 => "11111111",
		8538 to 8540 => "11111111",
		8601 to 8603 => "11111111",
		8664 to 8666 => "11111111",
		8731 to 8733 => "11111111",
		8794 to 8796 => "11111111",
		8857 to 8859 => "11111111",
		8920 to 8922 => "11111111",
		8987 to 8989 => "11111111",
		9050 to 9052 => "11111111",
		9113 to 9115 => "11111111",
		9176 to 9178 => "11111111",
		9243 to 9245 => "11111111",
		9306 to 9308 => "11111111",
		9369 to 9371 => "11111111",
		9432 to 9434 => "11111111",
		9499 to 9501 => "11111111",
		9562 to 9564 => "11111111",
		9625 to 9627 => "11111111",
		9688 to 9690 => "11111111",
		9755 to 9757 => "11111111",
		9818 to 9820 => "11111111",
		9881 to 9883 => "11111111",
		9944 to 9946 => "11111111",
		10011 to 10013 => "11111111",
		10074 to 10076 => "11111111",
		10137 to 10139 => "11111111",
		10200 to 10202 => "11111111",
		10267 to 10269 => "11111111",
		10330 to 10332 => "11111111",
		10393 to 10395 => "11111111",
		10456 to 10458 => "11111111",
		10523 to 10525 => "11111111",
		10586 to 10588 => "11111111",
		10649 to 10651 => "11111111",
		10712 to 10714 => "11111111",
		10779 to 10781 => "11111111",
		10842 to 10844 => "11111111",
		10905 to 10907 => "11111111",
		10968 to 10970 => "11111111",
		11035 to 11037 => "11111111",
		11098 to 11100 => "11111111",
		11161 to 11163 => "11111111",
		11224 to 11226 => "11111111",
		11291 to 11293 => "11111111",
		11354 to 11356 => "11111111",
		11417 to 11419 => "11111111",
		11480 to 11482 => "11111111",
		11547 to 11549 => "11111111",
		11610 to 11612 => "11111111",
		11673 to 11675 => "11111111",
		11736 to 11738 => "11111111",
		11803 to 11805 => "11111111",
		11866 to 11868 => "11111111",
		11929 to 11931 => "11111111",
		11992 to 11994 => "11111111",
		12059 to 12061 => "11111111",
		12122 to 12124 => "11111111",
		12185 to 12187 => "11111111",
		12248 to 12250 => "11111111",
		12315 to 12317 => "11111111",
		12378 to 12380 => "11111111",
		12441 to 12443 => "11111111",
		12504 to 12506 => "11111111",
		12571 to 12573 => "11111111",
		12634 to 12636 => "11111111",
		12697 to 12699 => "11111111",
		12760 to 12762 => "11111111",
		12827 to 12829 => "11111111",
		12890 to 12892 => "11111111",
		12953 to 12955 => "11111111",
		13016 to 13018 => "11111111",
		13083 to 13085 => "11111111",
		13146 to 13148 => "11111111",
		13209 to 13211 => "11111111",
		13272 to 13274 => "11111111",
		13339 to 13341 => "11111111",
		13402 to 13404 => "11111111",
		13465 to 13467 => "11111111",
		13528 to 13530 => "11111111",
		13595 to 13597 => "11111111",
		13658 to 13660 => "11111111",
		13721 to 13723 => "11111111",
		13784 to 13786 => "11111111",
		13851 to 13853 => "11111111",
		13914 to 13916 => "11111111",
		13977 to 13979 => "11111111",
		14040 to 14042 => "11111111",
		14107 to 14109 => "11111111",
		14170 to 14172 => "11111111",
		14233 to 14235 => "11111111",
		14296 to 14298 => "11111111",
		14363 to 14365 => "11111111",
		14426 to 14428 => "11111111",
		14489 to 14491 => "11111111",
		14552 to 14554 => "11111111",
		14619 to 14621 => "11111111",
		14682 to 14684 => "11111111",
		14745 to 14747 => "11111111",
		14808 to 14810 => "11111111",
		14875 to 14877 => "11111111",
		14938 to 14940 => "11111111",
		15001 to 15003 => "11111111",
		15064 to 15066 => "11111111",
		15131 to 15133 => "11111111",
		15194 to 15196 => "11111111",
		15257 to 15259 => "11111111",
		15320 to 15322 => "11111111",
		15387 to 15389 => "11111111",
		15450 to 15452 => "11111111",
		15513 to 15515 => "11111111",
		15576 to 15578 => "11111111",
		15643 to 15645 => "11111111",
		15706 to 15708 => "11111111",
		15769 to 15771 => "11111111",
		15832 to 15834 => "11111111",
		15899 to 15901 => "11111111",
		15962 to 15964 => "11111111",
		16025 to 16027 => "11111111",
		16088 to 16090 => "11111111",
		16155 to 16157 => "11111111",
		16218 to 16220 => "11111111",
		16281 to 16283 => "11111111",
		16344 to 16346 => "11111111",
		16411 to 16413 => "11111111",
		16474 to 16476 => "11111111",
		16537 to 16539 => "11111111",
		16600 to 16602 => "11111111",
		16667 to 16669 => "11111111",
		16730 to 16732 => "11111111",
		16793 to 16795 => "11111111",
		16856 to 16858 => "11111111",
		16923 to 16925 => "11111111",
		16986 to 16988 => "11111111",
		17049 to 17051 => "11111111",
		17112 to 17114 => "11111111",
		17179 to 17181 => "11111111",
		17242 to 17244 => "11111111",
		17305 to 17307 => "11111111",
		17368 to 17370 => "11111111",
		17435 to 17437 => "11111111",
		17498 to 17500 => "11111111",
		17561 to 17563 => "11111111",
		17624 to 17626 => "11111111",
		17691 to 17693 => "11111111",
		17754 to 17756 => "11111111",
		17817 to 17819 => "11111111",
		17880 to 17882 => "11111111",
		17947 to 17949 => "11111111",
		18010 to 18012 => "11111111",
		18073 to 18075 => "11111111",
		18136 to 18138 => "11111111",
		18203 to 18205 => "11111111",
		18266 to 18268 => "11111111",
		18329 to 18331 => "11111111",
		18392 to 18394 => "11111111",
		18459 to 18461 => "11111111",
		18522 to 18524 => "11111111",
		18585 to 18587 => "11111111",
		18648 to 18650 => "11111111",
		18715 to 18717 => "11111111",
		18778 to 18780 => "11111111",
		18841 to 18843 => "11111111",
		18904 to 18906 => "11111111",
		18971 to 18973 => "11111111",
		19034 to 19036 => "11111111",
		19097 to 19099 => "11111111",
		19160 to 19162 => "11111111",
		19227 to 19229 => "11111111",
		19290 to 19292 => "11111111",
		19353 to 19355 => "11111111",
		19416 to 19418 => "11111111",
		19483 to 19485 => "11111111",
		19546 to 19548 => "11111111",
		19609 to 19611 => "11111111",
		19672 to 19674 => "11111111",
		19739 to 19741 => "11111111",
		19802 to 19804 => "11111111",
		19865 to 19867 => "11111111",
		19928 to 19930 => "11111111",
		19995 to 19997 => "11111111",
		20058 to 20060 => "11111111",
		20121 to 20123 => "11111111",
		20184 to 20186 => "11111111",
		20251 to 20253 => "11111111",
		20314 to 20316 => "11111111",
		20377 to 20379 => "11111111",
		20440 to 20442 => "11111111",
		20507 to 20509 => "11111111",
		20570 to 20572 => "11111111",
		20633 to 20635 => "11111111",
		20696 to 20698 => "11111111",
		20763 to 20765 => "11111111",
		20826 to 20828 => "11111111",
		20889 to 20891 => "11111111",
		20952 to 20954 => "11111111",
		21019 to 21021 => "11111111",
		21082 to 21084 => "11111111",
		21145 to 21147 => "11111111",
		21208 to 21210 => "11111111",
		21275 to 21277 => "11111111",
		21338 to 21340 => "11111111",
		21401 to 21403 => "11111111",
		21464 to 21466 => "11111111",
		21531 to 21533 => "11111111",
		21594 to 21596 => "11111111",
		21657 to 21659 => "11111111",
		21720 to 21722 => "11111111",
		21787 to 21789 => "11111111",
		21850 to 21852 => "11111111",
		21913 to 21915 => "11111111",
		21976 to 21978 => "11111111",
		22043 to 22045 => "11111111",
		22106 to 22108 => "11111111",
		22169 to 22171 => "11111111",
		22232 to 22234 => "11111111",
		22299 to 22301 => "11111111",
		22362 to 22364 => "11111111",
		22425 to 22427 => "11111111",
		22488 to 22490 => "11111111",
		22555 to 22557 => "11111111",
		22618 to 22620 => "11111111",
		22681 to 22683 => "11111111",
		22744 to 22746 => "11111111",
		22811 to 22813 => "11111111",
		22874 to 22876 => "11111111",
		22937 to 22939 => "11111111",
		23000 to 23002 => "11111111",
		23067 to 23258 => "11111111",
		23323 to 23514 => "11111111",
		23579 to 23770 => "11111111",
		23835 to 23837 => "11111111",
		23898 to 23900 => "11111111",
		23961 to 23963 => "11111111",
		24024 to 24026 => "11111111",
		24091 to 24093 => "11111111",
		24154 to 24156 => "11111111",
		24217 to 24219 => "11111111",
		24280 to 24282 => "11111111",
		24347 to 24349 => "11111111",
		24410 to 24412 => "11111111",
		24473 to 24475 => "11111111",
		24536 to 24538 => "11111111",
		24603 to 24605 => "11111111",
		24666 to 24668 => "11111111",
		24729 to 24731 => "11111111",
		24792 to 24794 => "11111111",
		24859 to 24861 => "11111111",
		24922 to 24924 => "11111111",
		24985 to 24987 => "11111111",
		25048 to 25050 => "11111111",
		25115 to 25117 => "11111111",
		25178 to 25180 => "11111111",
		25241 to 25243 => "11111111",
		25304 to 25306 => "11111111",
		25371 to 25373 => "11111111",
		25434 to 25436 => "11111111",
		25497 to 25499 => "11111111",
		25560 to 25562 => "11111111",
		25627 to 25629 => "11111111",
		25690 to 25692 => "11111111",
		25753 to 25755 => "11111111",
		25816 to 25818 => "11111111",
		25883 to 25885 => "11111111",
		25946 to 25948 => "11111111",
		26009 to 26011 => "11111111",
		26072 to 26074 => "11111111",
		26139 to 26141 => "11111111",
		26202 to 26204 => "11111111",
		26265 to 26267 => "11111111",
		26328 to 26330 => "11111111",
		26395 to 26397 => "11111111",
		26458 to 26460 => "11111111",
		26521 to 26523 => "11111111",
		26584 to 26586 => "11111111",
		26651 to 26653 => "11111111",
		26714 to 26716 => "11111111",
		26777 to 26779 => "11111111",
		26840 to 26842 => "11111111",
		26907 to 26909 => "11111111",
		26970 to 26972 => "11111111",
		27033 to 27035 => "11111111",
		27096 to 27098 => "11111111",
		27163 to 27165 => "11111111",
		27226 to 27228 => "11111111",
		27289 to 27291 => "11111111",
		27352 to 27354 => "11111111",
		27419 to 27421 => "11111111",
		27482 to 27484 => "11111111",
		27545 to 27547 => "11111111",
		27608 to 27610 => "11111111",
		27675 to 27677 => "11111111",
		27738 to 27740 => "11111111",
		27801 to 27803 => "11111111",
		27864 to 27866 => "11111111",
		27931 to 27933 => "11111111",
		27994 to 27996 => "11111111",
		28057 to 28059 => "11111111",
		28120 to 28122 => "11111111",
		28187 to 28189 => "11111111",
		28250 to 28252 => "11111111",
		28313 to 28315 => "11111111",
		28376 to 28378 => "11111111",
		28443 to 28445 => "11111111",
		28506 to 28508 => "11111111",
		28569 to 28571 => "11111111",
		28632 to 28634 => "11111111",
		28699 to 28701 => "11111111",
		28762 to 28764 => "11111111",
		28825 to 28827 => "11111111",
		28888 to 28890 => "11111111",
		28955 to 28957 => "11111111",
		29018 to 29020 => "11111111",
		29081 to 29083 => "11111111",
		29144 to 29146 => "11111111",
		29211 to 29213 => "11111111",
		29274 to 29276 => "11111111",
		29337 to 29339 => "11111111",
		29400 to 29402 => "11111111",
		29467 to 29469 => "11111111",
		29530 to 29532 => "11111111",
		29593 to 29595 => "11111111",
		29656 to 29658 => "11111111",
		29723 to 29725 => "11111111",
		29786 to 29788 => "11111111",
		29849 to 29851 => "11111111",
		29912 to 29914 => "11111111",
		29979 to 29981 => "11111111",
		30042 to 30044 => "11111111",
		30105 to 30107 => "11111111",
		30168 to 30170 => "11111111",
		30235 to 30237 => "11111111",
		30298 to 30300 => "11111111",
		30361 to 30363 => "11111111",
		30424 to 30426 => "11111111",
		30491 to 30493 => "11111111",
		30554 to 30556 => "11111111",
		30617 to 30619 => "11111111",
		30680 to 30682 => "11111111",
		30747 to 30749 => "11111111",
		30810 to 30812 => "11111111",
		30873 to 30875 => "11111111",
		30936 to 30938 => "11111111",
		31003 to 31005 => "11111111",
		31066 to 31068 => "11111111",
		31129 to 31131 => "11111111",
		31192 to 31194 => "11111111",
		31259 to 31261 => "11111111",
		31322 to 31324 => "11111111",
		31385 to 31387 => "11111111",
		31448 to 31450 => "11111111",
		31515 to 31517 => "11111111",
		31578 to 31580 => "11111111",
		31641 to 31643 => "11111111",
		31704 to 31706 => "11111111",
		31771 to 31773 => "11111111",
		31834 to 31836 => "11111111",
		31897 to 31899 => "11111111",
		31960 to 31962 => "11111111",
		32027 to 32029 => "11111111",
		32090 to 32092 => "11111111",
		32153 to 32155 => "11111111",
		32216 to 32218 => "11111111",
		32283 to 32285 => "11111111",
		32346 to 32348 => "11111111",
		32409 to 32411 => "11111111",
		32472 to 32474 => "11111111",
		32539 to 32541 => "11111111",
		32602 to 32604 => "11111111",
		32665 to 32667 => "11111111",
		32728 to 32730 => "11111111",
		32795 to 32797 => "11111111",
		32858 to 32860 => "11111111",
		32921 to 32923 => "11111111",
		32984 to 32986 => "11111111",
		33051 to 33053 => "11111111",
		33114 to 33116 => "11111111",
		33177 to 33179 => "11111111",
		33240 to 33242 => "11111111",
		33307 to 33309 => "11111111",
		33370 to 33372 => "11111111",
		33433 to 33435 => "11111111",
		33496 to 33498 => "11111111",
		33563 to 33565 => "11111111",
		33626 to 33628 => "11111111",
		33689 to 33691 => "11111111",
		33752 to 33754 => "11111111",
		33819 to 33821 => "11111111",
		33882 to 33884 => "11111111",
		33945 to 33947 => "11111111",
		34008 to 34010 => "11111111",
		34075 to 34077 => "11111111",
		34138 to 34140 => "11111111",
		34201 to 34203 => "11111111",
		34264 to 34266 => "11111111",
		34331 to 34333 => "11111111",
		34394 to 34396 => "11111111",
		34457 to 34459 => "11111111",
		34520 to 34522 => "11111111",
		34587 to 34589 => "11111111",
		34650 to 34652 => "11111111",
		34713 to 34715 => "11111111",
		34776 to 34778 => "11111111",
		34843 to 34845 => "11111111",
		34906 to 34908 => "11111111",
		34969 to 34971 => "11111111",
		35032 to 35034 => "11111111",
		35099 to 35101 => "11111111",
		35162 to 35164 => "11111111",
		35225 to 35227 => "11111111",
		35288 to 35290 => "11111111",
		35355 to 35357 => "11111111",
		35418 to 35420 => "11111111",
		35481 to 35483 => "11111111",
		35544 to 35546 => "11111111",
		35611 to 35613 => "11111111",
		35674 to 35676 => "11111111",
		35737 to 35739 => "11111111",
		35800 to 35802 => "11111111",
		35867 to 35869 => "11111111",
		35930 to 35932 => "11111111",
		35993 to 35995 => "11111111",
		36056 to 36058 => "11111111",
		36123 to 36125 => "11111111",
		36186 to 36188 => "11111111",
		36249 to 36251 => "11111111",
		36312 to 36314 => "11111111",
		36379 to 36381 => "11111111",
		36442 to 36444 => "11111111",
		36505 to 36507 => "11111111",
		36568 to 36570 => "11111111",
		36635 to 36637 => "11111111",
		36698 to 36700 => "11111111",
		36761 to 36763 => "11111111",
		36824 to 36826 => "11111111",
		36891 to 36893 => "11111111",
		36954 to 36956 => "11111111",
		37017 to 37019 => "11111111",
		37080 to 37082 => "11111111",
		37147 to 37149 => "11111111",
		37210 to 37212 => "11111111",
		37273 to 37275 => "11111111",
		37336 to 37338 => "11111111",
		37403 to 37405 => "11111111",
		37466 to 37468 => "11111111",
		37529 to 37531 => "11111111",
		37592 to 37594 => "11111111",
		37659 to 37661 => "11111111",
		37722 to 37724 => "11111111",
		37785 to 37787 => "11111111",
		37848 to 37850 => "11111111",
		37915 to 37917 => "11111111",
		37978 to 37980 => "11111111",
		38041 to 38043 => "11111111",
		38104 to 38106 => "11111111",
		38171 to 38173 => "11111111",
		38234 to 38236 => "11111111",
		38297 to 38299 => "11111111",
		38360 to 38362 => "11111111",
		38427 to 38429 => "11111111",
		38490 to 38492 => "11111111",
		38553 to 38555 => "11111111",
		38616 to 38618 => "11111111",
		38683 to 38685 => "11111111",
		38746 to 38748 => "11111111",
		38809 to 38811 => "11111111",
		38872 to 38874 => "11111111",
		38939 to 38941 => "11111111",
		39002 to 39004 => "11111111",
		39065 to 39067 => "11111111",
		39128 to 39130 => "11111111",
		39195 to 39386 => "11111111",
		39451 to 39642 => "11111111",
		39707 to 39898 => "11111111",
		39963 to 39965 => "11111111",
		40026 to 40028 => "11111111",
		40089 to 40091 => "11111111",
		40152 to 40154 => "11111111",
		40219 to 40221 => "11111111",
		40282 to 40284 => "11111111",
		40345 to 40347 => "11111111",
		40408 to 40410 => "11111111",
		40475 to 40477 => "11111111",
		40538 to 40540 => "11111111",
		40601 to 40603 => "11111111",
		40664 to 40666 => "11111111",
		40731 to 40733 => "11111111",
		40794 to 40796 => "11111111",
		40857 to 40859 => "11111111",
		40920 to 40922 => "11111111",
		40987 to 40989 => "11111111",
		41050 to 41052 => "11111111",
		41113 to 41115 => "11111111",
		41176 to 41178 => "11111111",
		41243 to 41245 => "11111111",
		41306 to 41308 => "11111111",
		41369 to 41371 => "11111111",
		41432 to 41434 => "11111111",
		41499 to 41501 => "11111111",
		41562 to 41564 => "11111111",
		41625 to 41627 => "11111111",
		41688 to 41690 => "11111111",
		41755 to 41757 => "11111111",
		41818 to 41820 => "11111111",
		41881 to 41883 => "11111111",
		41944 to 41946 => "11111111",
		42011 to 42013 => "11111111",
		42074 to 42076 => "11111111",
		42137 to 42139 => "11111111",
		42200 to 42202 => "11111111",
		42267 to 42269 => "11111111",
		42330 to 42332 => "11111111",
		42393 to 42395 => "11111111",
		42456 to 42458 => "11111111",
		42523 to 42525 => "11111111",
		42586 to 42588 => "11111111",
		42649 to 42651 => "11111111",
		42712 to 42714 => "11111111",
		42779 to 42781 => "11111111",
		42842 to 42844 => "11111111",
		42905 to 42907 => "11111111",
		42968 to 42970 => "11111111",
		43035 to 43037 => "11111111",
		43098 to 43100 => "11111111",
		43161 to 43163 => "11111111",
		43224 to 43226 => "11111111",
		43291 to 43293 => "11111111",
		43354 to 43356 => "11111111",
		43417 to 43419 => "11111111",
		43480 to 43482 => "11111111",
		43547 to 43549 => "11111111",
		43610 to 43612 => "11111111",
		43673 to 43675 => "11111111",
		43736 to 43738 => "11111111",
		43803 to 43805 => "11111111",
		43866 to 43868 => "11111111",
		43929 to 43931 => "11111111",
		43992 to 43994 => "11111111",
		44059 to 44061 => "11111111",
		44122 to 44124 => "11111111",
		44185 to 44187 => "11111111",
		44248 to 44250 => "11111111",
		44315 to 44317 => "11111111",
		44378 to 44380 => "11111111",
		44441 to 44443 => "11111111",
		44504 to 44506 => "11111111",
		44571 to 44573 => "11111111",
		44634 to 44636 => "11111111",
		44697 to 44699 => "11111111",
		44760 to 44762 => "11111111",
		44827 to 44829 => "11111111",
		44890 to 44892 => "11111111",
		44953 to 44955 => "11111111",
		45016 to 45018 => "11111111",
		45083 to 45085 => "11111111",
		45146 to 45148 => "11111111",
		45209 to 45211 => "11111111",
		45272 to 45274 => "11111111",
		45339 to 45341 => "11111111",
		45402 to 45404 => "11111111",
		45465 to 45467 => "11111111",
		45528 to 45530 => "11111111",
		45595 to 45597 => "11111111",
		45658 to 45660 => "11111111",
		45721 to 45723 => "11111111",
		45784 to 45786 => "11111111",
		45851 to 45853 => "11111111",
		45914 to 45916 => "11111111",
		45977 to 45979 => "11111111",
		46040 to 46042 => "11111111",
		46107 to 46109 => "11111111",
		46170 to 46172 => "11111111",
		46233 to 46235 => "11111111",
		46296 to 46298 => "11111111",
		46363 to 46365 => "11111111",
		46426 to 46428 => "11111111",
		46489 to 46491 => "11111111",
		46552 to 46554 => "11111111",
		46619 to 46621 => "11111111",
		46682 to 46684 => "11111111",
		46745 to 46747 => "11111111",
		46808 to 46810 => "11111111",
		46875 to 46877 => "11111111",
		46938 to 46940 => "11111111",
		47001 to 47003 => "11111111",
		47064 to 47066 => "11111111",
		47131 to 47133 => "11111111",
		47194 to 47196 => "11111111",
		47257 to 47259 => "11111111",
		47320 to 47322 => "11111111",
		47387 to 47389 => "11111111",
		47450 to 47452 => "11111111",
		47513 to 47515 => "11111111",
		47576 to 47578 => "11111111",
		47643 to 47645 => "11111111",
		47706 to 47708 => "11111111",
		47769 to 47771 => "11111111",
		47832 to 47834 => "11111111",
		47899 to 47901 => "11111111",
		47962 to 47964 => "11111111",
		48025 to 48027 => "11111111",
		48088 to 48090 => "11111111",
		48155 to 48157 => "11111111",
		48218 to 48220 => "11111111",
		48281 to 48283 => "11111111",
		48344 to 48346 => "11111111",
		48411 to 48413 => "11111111",
		48474 to 48476 => "11111111",
		48537 to 48539 => "11111111",
		48600 to 48602 => "11111111",
		48667 to 48669 => "11111111",
		48730 to 48732 => "11111111",
		48793 to 48795 => "11111111",
		48856 to 48858 => "11111111",
		48923 to 48925 => "11111111",
		48986 to 48988 => "11111111",
		49049 to 49051 => "11111111",
		49112 to 49114 => "11111111",
		49179 to 49181 => "11111111",
		49242 to 49244 => "11111111",
		49305 to 49307 => "11111111",
		49368 to 49370 => "11111111",
		49435 to 49437 => "11111111",
		49498 to 49500 => "11111111",
		49561 to 49563 => "11111111",
		49624 to 49626 => "11111111",
		49691 to 49693 => "11111111",
		49754 to 49756 => "11111111",
		49817 to 49819 => "11111111",
		49880 to 49882 => "11111111",
		49947 to 49949 => "11111111",
		50010 to 50012 => "11111111",
		50073 to 50075 => "11111111",
		50136 to 50138 => "11111111",
		50203 to 50205 => "11111111",
		50266 to 50268 => "11111111",
		50329 to 50331 => "11111111",
		50392 to 50394 => "11111111",
		50459 to 50461 => "11111111",
		50522 to 50524 => "11111111",
		50585 to 50587 => "11111111",
		50648 to 50650 => "11111111",
		50715 to 50717 => "11111111",
		50778 to 50780 => "11111111",
		50841 to 50843 => "11111111",
		50904 to 50906 => "11111111",
		50971 to 50973 => "11111111",
		51034 to 51036 => "11111111",
		51097 to 51099 => "11111111",
		51160 to 51162 => "11111111",
		51227 to 51229 => "11111111",
		51290 to 51292 => "11111111",
		51353 to 51355 => "11111111",
		51416 to 51418 => "11111111",
		51483 to 51485 => "11111111",
		51546 to 51548 => "11111111",
		51609 to 51611 => "11111111",
		51672 to 51674 => "11111111",
		51739 to 51741 => "11111111",
		51802 to 51804 => "11111111",
		51865 to 51867 => "11111111",
		51928 to 51930 => "11111111",
		51995 to 51997 => "11111111",
		52058 to 52060 => "11111111",
		52121 to 52123 => "11111111",
		52184 to 52186 => "11111111",
		52251 to 52253 => "11111111",
		52314 to 52316 => "11111111",
		52377 to 52379 => "11111111",
		52440 to 52442 => "11111111",
		52507 to 52509 => "11111111",
		52570 to 52572 => "11111111",
		52633 to 52635 => "11111111",
		52696 to 52698 => "11111111",
		52763 to 52765 => "11111111",
		52826 to 52828 => "11111111",
		52889 to 52891 => "11111111",
		52952 to 52954 => "11111111",
		53019 to 53021 => "11111111",
		53082 to 53084 => "11111111",
		53145 to 53147 => "11111111",
		53208 to 53210 => "11111111",
		53275 to 53277 => "11111111",
		53338 to 53340 => "11111111",
		53401 to 53403 => "11111111",
		53464 to 53466 => "11111111",
		53531 to 53533 => "11111111",
		53594 to 53596 => "11111111",
		53657 to 53659 => "11111111",
		53720 to 53722 => "11111111",
		53787 to 53789 => "11111111",
		53850 to 53852 => "11111111",
		53913 to 53915 => "11111111",
		53976 to 53978 => "11111111",
		54043 to 54045 => "11111111",
		54106 to 54108 => "11111111",
		54169 to 54171 => "11111111",
		54232 to 54234 => "11111111",
		54299 to 54301 => "11111111",
		54362 to 54364 => "11111111",
		54425 to 54427 => "11111111",
		54488 to 54490 => "11111111",
		54555 to 54557 => "11111111",
		54618 to 54620 => "11111111",
		54681 to 54683 => "11111111",
		54744 to 54746 => "11111111",
		54811 to 54813 => "11111111",
		54874 to 54876 => "11111111",
		54937 to 54939 => "11111111",
		55000 to 55002 => "11111111",
		55067 to 55069 => "11111111",
		55130 to 55132 => "11111111",
		55193 to 55195 => "11111111",
		55256 to 55258 => "11111111",
		55323 to 55514 => "11111111",
		55579 to 55770 => "11111111",
		55835 to 56026 => "11111111",
