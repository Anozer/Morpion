		49280 => '1',
		49281 => '1',
		49282 => '1',
		49283 => '1',
		49284 => '1',
		49285 => '1',
		49286 => '1',
		49287 => '1',
		49288 => '1',
		49289 => '1',
		49290 => '1',
		49291 => '1',
		49292 => '1',
		49293 => '1',
		49294 => '1',
		49295 => '1',
		49296 => '1',
		49297 => '1',
		49298 => '1',
		49299 => '1',
		49300 => '1',
		49301 => '1',
		49302 => '1',
		49303 => '1',
		49304 => '1',
		49305 => '1',
		49306 => '1',
		49307 => '1',
		49308 => '1',
		49309 => '1',
		49310 => '1',
		49311 => '1',
		49312 => '1',
		49313 => '1',
		49314 => '1',
		49315 => '1',
		49316 => '1',
		49317 => '1',
		49318 => '1',
		49319 => '1',
		49320 => '1',
		49321 => '1',
		49322 => '1',
		49323 => '1',
		49324 => '1',
		49325 => '1',
		49326 => '1',
		49327 => '1',
		49328 => '1',
		49329 => '1',
		49330 => '1',
		49331 => '1',
		49332 => '1',
		49333 => '1',
		49334 => '1',
		49335 => '1',
		49336 => '1',
		49337 => '1',
		49338 => '1',
		49339 => '1',
		49340 => '1',
		49341 => '1',
		49342 => '1',
		49343 => '1',
		49344 => '1',
		49345 => '1',
		49346 => '1',
		49347 => '1',
		49348 => '1',
		49349 => '1',
		49350 => '1',
		49351 => '1',
		49352 => '1',
		49353 => '1',
		49354 => '1',
		49355 => '1',
		49356 => '1',
		49357 => '1',
		49358 => '1',
		49359 => '1',
		49360 => '1',
		49361 => '1',
		49362 => '1',
		49363 => '1',
		49364 => '1',
		49365 => '1',
		49366 => '1',
		49367 => '1',
		49368 => '1',
		49369 => '1',
		49370 => '1',
		49371 => '1',
		49372 => '1',
		49373 => '1',
		49374 => '1',
		49375 => '1',
		49376 => '1',
		49377 => '1',
		49378 => '1',
		49379 => '1',
		49380 => '1',
		49381 => '1',
		49382 => '1',
		49383 => '1',
		49384 => '1',
		49385 => '1',
		49386 => '1',
		49387 => '1',
		49388 => '1',
		49389 => '1',
		49390 => '1',
		49391 => '1',
		49392 => '1',
		49393 => '1',
		49394 => '1',
		49395 => '1',
		49396 => '1',
		49397 => '1',
		49398 => '1',
		49399 => '1',
		49400 => '1',
		49401 => '1',
		49402 => '1',
		49403 => '1',
		49404 => '1',
		49405 => '1',
		49406 => '1',
		49407 => '1',
		49408 => '1',
		49409 => '1',
		49410 => '1',
		49411 => '1',
		49412 => '1',
		49413 => '1',
		49414 => '1',
		49415 => '1',
		49416 => '1',
		49417 => '1',
		49418 => '1',
		49419 => '1',
		49420 => '1',
		49421 => '1',
		49422 => '1',
		49423 => '1',
		49424 => '1',
		49425 => '1',
		49426 => '1',
		49427 => '1',
		49428 => '1',
		49429 => '1',
		49430 => '1',
		49431 => '1',
		49432 => '1',
		49433 => '1',
		49434 => '1',
		49435 => '1',
		49436 => '1',
		49437 => '1',
		49438 => '1',
		49439 => '1',
		49440 => '1',
		49441 => '1',
		49442 => '1',
		49443 => '1',
		49444 => '1',
		49445 => '1',
		49446 => '1',
		49447 => '1',
		49448 => '1',
		49449 => '1',
		49450 => '1',
		49451 => '1',
		49452 => '1',
		49453 => '1',
		49454 => '1',
		49455 => '1',
		49456 => '1',
		49457 => '1',
		49458 => '1',
		49459 => '1',
		49460 => '1',
		49461 => '1',
		49462 => '1',
		49463 => '1',
		49464 => '1',
		49465 => '1',
		49466 => '1',
		49467 => '1',
		49468 => '1',
		49469 => '1',
		49470 => '1',
		49471 => '1',
		49472 => '1',
		49473 => '1',
		49474 => '1',
		49475 => '1',
		49476 => '1',
		49477 => '1',
		49478 => '1',
		49479 => '1',
		49480 => '1',
		49481 => '1',
		49482 => '1',
		49483 => '1',
		49484 => '1',
		49485 => '1',
		49486 => '1',
		49487 => '1',
		49488 => '1',
		49489 => '1',
		49490 => '1',
		49491 => '1',
		49492 => '1',
		49493 => '1',
		49494 => '1',
		49495 => '1',
		49496 => '1',
		49497 => '1',
		49498 => '1',
		49499 => '1',
		49500 => '1',
		49501 => '1',
		49502 => '1',
		49503 => '1',
		49504 => '1',
		49505 => '1',
		49506 => '1',
		49507 => '1',
		49508 => '1',
		49509 => '1',
		49510 => '1',
		49511 => '1',
		49512 => '1',
		49513 => '1',
		49514 => '1',
		49515 => '1',
		49516 => '1',
		49517 => '1',
		49518 => '1',
		49519 => '1',
		49520 => '1',
		49521 => '1',
		49522 => '1',
		49523 => '1',
		49524 => '1',
		49525 => '1',
		49526 => '1',
		49527 => '1',
		49528 => '1',
		49529 => '1',
		49530 => '1',
		49531 => '1',
		49532 => '1',
		49533 => '1',
		49534 => '1',
		49535 => '1',
		49536 => '1',
		49537 => '1',
		49538 => '1',
		49539 => '1',
		49540 => '1',
		49541 => '1',
		49542 => '1',
		49543 => '1',
		49544 => '1',
		49545 => '1',
		49546 => '1',
		49547 => '1',
		49548 => '1',
		49549 => '1',
		49550 => '1',
		49551 => '1',
		49552 => '1',
		49553 => '1',
		49554 => '1',
		49555 => '1',
		49556 => '1',
		49557 => '1',
		49558 => '1',
		49559 => '1',
		49560 => '1',
		49561 => '1',
		49562 => '1',
		49563 => '1',
		49564 => '1',
		49565 => '1',
		49566 => '1',
		49567 => '1',
		49568 => '1',
		49569 => '1',
		49570 => '1',
		49571 => '1',
		49572 => '1',
		49573 => '1',
		49574 => '1',
		49575 => '1',
		49576 => '1',
		49577 => '1',
		49578 => '1',
		49579 => '1',
		49580 => '1',
		49581 => '1',
		49582 => '1',
		49583 => '1',
		49584 => '1',
		49585 => '1',
		49586 => '1',
		49587 => '1',
		49588 => '1',
		49589 => '1',
		49590 => '1',
		49591 => '1',
		49592 => '1',
		49593 => '1',
		49594 => '1',
		49595 => '1',
		49596 => '1',
		49597 => '1',
		49598 => '1',
		49599 => '1',
		49600 => '1',
		49601 => '1',
		49602 => '1',
		49603 => '1',
		49604 => '1',
		49605 => '1',
		49606 => '1',
		49607 => '1',
		49608 => '1',
		49609 => '1',
		49610 => '1',
		49611 => '1',
		49612 => '1',
		49613 => '1',
		49614 => '1',
		49615 => '1',
		49616 => '1',
		49617 => '1',
		49618 => '1',
		49619 => '1',
		49620 => '1',
		49621 => '1',
		49622 => '1',
		49623 => '1',
		49624 => '1',
		49625 => '1',
		49626 => '1',
		49627 => '1',
		49628 => '1',
		49629 => '1',
		49630 => '1',
		49631 => '1',
		49632 => '1',
		49633 => '1',
		49634 => '1',
		49635 => '1',
		49636 => '1',
		49637 => '1',
		49638 => '1',
		49639 => '1',
		49640 => '1',
		49641 => '1',
		49642 => '1',
		49643 => '1',
		49644 => '1',
		49645 => '1',
		49646 => '1',
		49647 => '1',
		49648 => '1',
		49649 => '1',
		49650 => '1',
		49651 => '1',
		49652 => '1',
		49653 => '1',
		49654 => '1',
		49655 => '1',
		49656 => '1',
		49657 => '1',
		49658 => '1',
		49659 => '1',
		50304 => '1',
		50305 => '1',
		50306 => '1',
		50307 => '1',
		50308 => '1',
		50309 => '1',
		50310 => '1',
		50311 => '1',
		50312 => '1',
		50313 => '1',
		50314 => '1',
		50315 => '1',
		50316 => '1',
		50317 => '1',
		50318 => '1',
		50319 => '1',
		50320 => '1',
		50321 => '1',
		50322 => '1',
		50323 => '1',
		50324 => '1',
		50325 => '1',
		50326 => '1',
		50327 => '1',
		50328 => '1',
		50329 => '1',
		50330 => '1',
		50331 => '1',
		50332 => '1',
		50333 => '1',
		50334 => '1',
		50335 => '1',
		50336 => '1',
		50337 => '1',
		50338 => '1',
		50339 => '1',
		50340 => '1',
		50341 => '1',
		50342 => '1',
		50343 => '1',
		50344 => '1',
		50345 => '1',
		50346 => '1',
		50347 => '1',
		50348 => '1',
		50349 => '1',
		50350 => '1',
		50351 => '1',
		50352 => '1',
		50353 => '1',
		50354 => '1',
		50355 => '1',
		50356 => '1',
		50357 => '1',
		50358 => '1',
		50359 => '1',
		50360 => '1',
		50361 => '1',
		50362 => '1',
		50363 => '1',
		50364 => '1',
		50365 => '1',
		50366 => '1',
		50367 => '1',
		50368 => '1',
		50369 => '1',
		50370 => '1',
		50371 => '1',
		50372 => '1',
		50373 => '1',
		50374 => '1',
		50375 => '1',
		50376 => '1',
		50377 => '1',
		50378 => '1',
		50379 => '1',
		50380 => '1',
		50381 => '1',
		50382 => '1',
		50383 => '1',
		50384 => '1',
		50385 => '1',
		50386 => '1',
		50387 => '1',
		50388 => '1',
		50389 => '1',
		50390 => '1',
		50391 => '1',
		50392 => '1',
		50393 => '1',
		50394 => '1',
		50395 => '1',
		50396 => '1',
		50397 => '1',
		50398 => '1',
		50399 => '1',
		50400 => '1',
		50401 => '1',
		50402 => '1',
		50403 => '1',
		50404 => '1',
		50405 => '1',
		50406 => '1',
		50407 => '1',
		50408 => '1',
		50409 => '1',
		50410 => '1',
		50411 => '1',
		50412 => '1',
		50413 => '1',
		50414 => '1',
		50415 => '1',
		50416 => '1',
		50417 => '1',
		50418 => '1',
		50419 => '1',
		50420 => '1',
		50421 => '1',
		50422 => '1',
		50423 => '1',
		50424 => '1',
		50425 => '1',
		50426 => '1',
		50427 => '1',
		50428 => '1',
		50429 => '1',
		50430 => '1',
		50431 => '1',
		50432 => '1',
		50433 => '1',
		50434 => '1',
		50435 => '1',
		50436 => '1',
		50437 => '1',
		50438 => '1',
		50439 => '1',
		50440 => '1',
		50441 => '1',
		50442 => '1',
		50443 => '1',
		50444 => '1',
		50445 => '1',
		50446 => '1',
		50447 => '1',
		50448 => '1',
		50449 => '1',
		50450 => '1',
		50451 => '1',
		50452 => '1',
		50453 => '1',
		50454 => '1',
		50455 => '1',
		50456 => '1',
		50457 => '1',
		50458 => '1',
		50459 => '1',
		50460 => '1',
		50461 => '1',
		50462 => '1',
		50463 => '1',
		50464 => '1',
		50465 => '1',
		50466 => '1',
		50467 => '1',
		50468 => '1',
		50469 => '1',
		50470 => '1',
		50471 => '1',
		50472 => '1',
		50473 => '1',
		50474 => '1',
		50475 => '1',
		50476 => '1',
		50477 => '1',
		50478 => '1',
		50479 => '1',
		50480 => '1',
		50481 => '1',
		50482 => '1',
		50483 => '1',
		50484 => '1',
		50485 => '1',
		50486 => '1',
		50487 => '1',
		50488 => '1',
		50489 => '1',
		50490 => '1',
		50491 => '1',
		50492 => '1',
		50493 => '1',
		50494 => '1',
		50495 => '1',
		50496 => '1',
		50497 => '1',
		50498 => '1',
		50499 => '1',
		50500 => '1',
		50501 => '1',
		50502 => '1',
		50503 => '1',
		50504 => '1',
		50505 => '1',
		50506 => '1',
		50507 => '1',
		50508 => '1',
		50509 => '1',
		50510 => '1',
		50511 => '1',
		50512 => '1',
		50513 => '1',
		50514 => '1',
		50515 => '1',
		50516 => '1',
		50517 => '1',
		50518 => '1',
		50519 => '1',
		50520 => '1',
		50521 => '1',
		50522 => '1',
		50523 => '1',
		50524 => '1',
		50525 => '1',
		50526 => '1',
		50527 => '1',
		50528 => '1',
		50529 => '1',
		50530 => '1',
		50531 => '1',
		50532 => '1',
		50533 => '1',
		50534 => '1',
		50535 => '1',
		50536 => '1',
		50537 => '1',
		50538 => '1',
		50539 => '1',
		50540 => '1',
		50541 => '1',
		50542 => '1',
		50543 => '1',
		50544 => '1',
		50545 => '1',
		50546 => '1',
		50547 => '1',
		50548 => '1',
		50549 => '1',
		50550 => '1',
		50551 => '1',
		50552 => '1',
		50553 => '1',
		50554 => '1',
		50555 => '1',
		50556 => '1',
		50557 => '1',
		50558 => '1',
		50559 => '1',
		50560 => '1',
		50561 => '1',
		50562 => '1',
		50563 => '1',
		50564 => '1',
		50565 => '1',
		50566 => '1',
		50567 => '1',
		50568 => '1',
		50569 => '1',
		50570 => '1',
		50571 => '1',
		50572 => '1',
		50573 => '1',
		50574 => '1',
		50575 => '1',
		50576 => '1',
		50577 => '1',
		50578 => '1',
		50579 => '1',
		50580 => '1',
		50581 => '1',
		50582 => '1',
		50583 => '1',
		50584 => '1',
		50585 => '1',
		50586 => '1',
		50587 => '1',
		50588 => '1',
		50589 => '1',
		50590 => '1',
		50591 => '1',
		50592 => '1',
		50593 => '1',
		50594 => '1',
		50595 => '1',
		50596 => '1',
		50597 => '1',
		50598 => '1',
		50599 => '1',
		50600 => '1',
		50601 => '1',
		50602 => '1',
		50603 => '1',
		50604 => '1',
		50605 => '1',
		50606 => '1',
		50607 => '1',
		50608 => '1',
		50609 => '1',
		50610 => '1',
		50611 => '1',
		50612 => '1',
		50613 => '1',
		50614 => '1',
		50615 => '1',
		50616 => '1',
		50617 => '1',
		50618 => '1',
		50619 => '1',
		50620 => '1',
		50621 => '1',
		50622 => '1',
		50623 => '1',
		50624 => '1',
		50625 => '1',
		50626 => '1',
		50627 => '1',
		50628 => '1',
		50629 => '1',
		50630 => '1',
		50631 => '1',
		50632 => '1',
		50633 => '1',
		50634 => '1',
		50635 => '1',
		50636 => '1',
		50637 => '1',
		50638 => '1',
		50639 => '1',
		50640 => '1',
		50641 => '1',
		50642 => '1',
		50643 => '1',
		50644 => '1',
		50645 => '1',
		50646 => '1',
		50647 => '1',
		50648 => '1',
		50649 => '1',
		50650 => '1',
		50651 => '1',
		50652 => '1',
		50653 => '1',
		50654 => '1',
		50655 => '1',
		50656 => '1',
		50657 => '1',
		50658 => '1',
		50659 => '1',
		50660 => '1',
		50661 => '1',
		50662 => '1',
		50663 => '1',
		50664 => '1',
		50665 => '1',
		50666 => '1',
		50667 => '1',
		50668 => '1',
		50669 => '1',
		50670 => '1',
		50671 => '1',
		50672 => '1',
		50673 => '1',
		50674 => '1',
		50675 => '1',
		50676 => '1',
		50677 => '1',
		50678 => '1',
		50679 => '1',
		50680 => '1',
		50681 => '1',
		50682 => '1',
		50683 => '1',
		51328 => '1',
		51329 => '1',
		51330 => '1',
		51331 => '1',
		51332 => '1',
		51333 => '1',
		51334 => '1',
		51335 => '1',
		51336 => '1',
		51337 => '1',
		51338 => '1',
		51339 => '1',
		51340 => '1',
		51341 => '1',
		51342 => '1',
		51343 => '1',
		51344 => '1',
		51345 => '1',
		51346 => '1',
		51347 => '1',
		51348 => '1',
		51349 => '1',
		51350 => '1',
		51351 => '1',
		51352 => '1',
		51353 => '1',
		51354 => '1',
		51355 => '1',
		51356 => '1',
		51357 => '1',
		51358 => '1',
		51359 => '1',
		51360 => '1',
		51361 => '1',
		51362 => '1',
		51363 => '1',
		51364 => '1',
		51365 => '1',
		51366 => '1',
		51367 => '1',
		51368 => '1',
		51369 => '1',
		51370 => '1',
		51371 => '1',
		51372 => '1',
		51373 => '1',
		51374 => '1',
		51375 => '1',
		51376 => '1',
		51377 => '1',
		51378 => '1',
		51379 => '1',
		51380 => '1',
		51381 => '1',
		51382 => '1',
		51383 => '1',
		51384 => '1',
		51385 => '1',
		51386 => '1',
		51387 => '1',
		51388 => '1',
		51389 => '1',
		51390 => '1',
		51391 => '1',
		51392 => '1',
		51393 => '1',
		51394 => '1',
		51395 => '1',
		51396 => '1',
		51397 => '1',
		51398 => '1',
		51399 => '1',
		51400 => '1',
		51401 => '1',
		51402 => '1',
		51403 => '1',
		51404 => '1',
		51405 => '1',
		51406 => '1',
		51407 => '1',
		51408 => '1',
		51409 => '1',
		51410 => '1',
		51411 => '1',
		51412 => '1',
		51413 => '1',
		51414 => '1',
		51415 => '1',
		51416 => '1',
		51417 => '1',
		51418 => '1',
		51419 => '1',
		51420 => '1',
		51421 => '1',
		51422 => '1',
		51423 => '1',
		51424 => '1',
		51425 => '1',
		51426 => '1',
		51427 => '1',
		51428 => '1',
		51429 => '1',
		51430 => '1',
		51431 => '1',
		51432 => '1',
		51433 => '1',
		51434 => '1',
		51435 => '1',
		51436 => '1',
		51437 => '1',
		51438 => '1',
		51439 => '1',
		51440 => '1',
		51441 => '1',
		51442 => '1',
		51443 => '1',
		51444 => '1',
		51445 => '1',
		51446 => '1',
		51447 => '1',
		51448 => '1',
		51449 => '1',
		51450 => '1',
		51451 => '1',
		51452 => '1',
		51453 => '1',
		51454 => '1',
		51455 => '1',
		51456 => '1',
		51457 => '1',
		51458 => '1',
		51459 => '1',
		51460 => '1',
		51461 => '1',
		51462 => '1',
		51463 => '1',
		51464 => '1',
		51465 => '1',
		51466 => '1',
		51467 => '1',
		51468 => '1',
		51469 => '1',
		51470 => '1',
		51471 => '1',
		51472 => '1',
		51473 => '1',
		51474 => '1',
		51475 => '1',
		51476 => '1',
		51477 => '1',
		51478 => '1',
		51479 => '1',
		51480 => '1',
		51481 => '1',
		51482 => '1',
		51483 => '1',
		51484 => '1',
		51485 => '1',
		51486 => '1',
		51487 => '1',
		51488 => '1',
		51489 => '1',
		51490 => '1',
		51491 => '1',
		51492 => '1',
		51493 => '1',
		51494 => '1',
		51495 => '1',
		51496 => '1',
		51497 => '1',
		51498 => '1',
		51499 => '1',
		51500 => '1',
		51501 => '1',
		51502 => '1',
		51503 => '1',
		51504 => '1',
		51505 => '1',
		51506 => '1',
		51507 => '1',
		51508 => '1',
		51509 => '1',
		51510 => '1',
		51511 => '1',
		51512 => '1',
		51513 => '1',
		51514 => '1',
		51515 => '1',
		51516 => '1',
		51517 => '1',
		51518 => '1',
		51519 => '1',
		51520 => '1',
		51521 => '1',
		51522 => '1',
		51523 => '1',
		51524 => '1',
		51525 => '1',
		51526 => '1',
		51527 => '1',
		51528 => '1',
		51529 => '1',
		51530 => '1',
		51531 => '1',
		51532 => '1',
		51533 => '1',
		51534 => '1',
		51535 => '1',
		51536 => '1',
		51537 => '1',
		51538 => '1',
		51539 => '1',
		51540 => '1',
		51541 => '1',
		51542 => '1',
		51543 => '1',
		51544 => '1',
		51545 => '1',
		51546 => '1',
		51547 => '1',
		51548 => '1',
		51549 => '1',
		51550 => '1',
		51551 => '1',
		51552 => '1',
		51553 => '1',
		51554 => '1',
		51555 => '1',
		51556 => '1',
		51557 => '1',
		51558 => '1',
		51559 => '1',
		51560 => '1',
		51561 => '1',
		51562 => '1',
		51563 => '1',
		51564 => '1',
		51565 => '1',
		51566 => '1',
		51567 => '1',
		51568 => '1',
		51569 => '1',
		51570 => '1',
		51571 => '1',
		51572 => '1',
		51573 => '1',
		51574 => '1',
		51575 => '1',
		51576 => '1',
		51577 => '1',
		51578 => '1',
		51579 => '1',
		51580 => '1',
		51581 => '1',
		51582 => '1',
		51583 => '1',
		51584 => '1',
		51585 => '1',
		51586 => '1',
		51587 => '1',
		51588 => '1',
		51589 => '1',
		51590 => '1',
		51591 => '1',
		51592 => '1',
		51593 => '1',
		51594 => '1',
		51595 => '1',
		51596 => '1',
		51597 => '1',
		51598 => '1',
		51599 => '1',
		51600 => '1',
		51601 => '1',
		51602 => '1',
		51603 => '1',
		51604 => '1',
		51605 => '1',
		51606 => '1',
		51607 => '1',
		51608 => '1',
		51609 => '1',
		51610 => '1',
		51611 => '1',
		51612 => '1',
		51613 => '1',
		51614 => '1',
		51615 => '1',
		51616 => '1',
		51617 => '1',
		51618 => '1',
		51619 => '1',
		51620 => '1',
		51621 => '1',
		51622 => '1',
		51623 => '1',
		51624 => '1',
		51625 => '1',
		51626 => '1',
		51627 => '1',
		51628 => '1',
		51629 => '1',
		51630 => '1',
		51631 => '1',
		51632 => '1',
		51633 => '1',
		51634 => '1',
		51635 => '1',
		51636 => '1',
		51637 => '1',
		51638 => '1',
		51639 => '1',
		51640 => '1',
		51641 => '1',
		51642 => '1',
		51643 => '1',
		51644 => '1',
		51645 => '1',
		51646 => '1',
		51647 => '1',
		51648 => '1',
		51649 => '1',
		51650 => '1',
		51651 => '1',
		51652 => '1',
		51653 => '1',
		51654 => '1',
		51655 => '1',
		51656 => '1',
		51657 => '1',
		51658 => '1',
		51659 => '1',
		51660 => '1',
		51661 => '1',
		51662 => '1',
		51663 => '1',
		51664 => '1',
		51665 => '1',
		51666 => '1',
		51667 => '1',
		51668 => '1',
		51669 => '1',
		51670 => '1',
		51671 => '1',
		51672 => '1',
		51673 => '1',
		51674 => '1',
		51675 => '1',
		51676 => '1',
		51677 => '1',
		51678 => '1',
		51679 => '1',
		51680 => '1',
		51681 => '1',
		51682 => '1',
		51683 => '1',
		51684 => '1',
		51685 => '1',
		51686 => '1',
		51687 => '1',
		51688 => '1',
		51689 => '1',
		51690 => '1',
		51691 => '1',
		51692 => '1',
		51693 => '1',
		51694 => '1',
		51695 => '1',
		51696 => '1',
		51697 => '1',
		51698 => '1',
		51699 => '1',
		51700 => '1',
		51701 => '1',
		51702 => '1',
		51703 => '1',
		51704 => '1',
		51705 => '1',
		51706 => '1',
		51707 => '1',
		52352 => '1',
		52353 => '1',
		52354 => '1',
		52355 => '1',
		52356 => '1',
		52357 => '1',
		52358 => '1',
		52359 => '1',
		52360 => '1',
		52361 => '1',
		52362 => '1',
		52363 => '1',
		52364 => '1',
		52365 => '1',
		52366 => '1',
		52367 => '1',
		52368 => '1',
		52369 => '1',
		52370 => '1',
		52371 => '1',
		52372 => '1',
		52373 => '1',
		52374 => '1',
		52375 => '1',
		52376 => '1',
		52377 => '1',
		52378 => '1',
		52379 => '1',
		52380 => '1',
		52381 => '1',
		52382 => '1',
		52383 => '1',
		52384 => '1',
		52385 => '1',
		52386 => '1',
		52387 => '1',
		52388 => '1',
		52389 => '1',
		52390 => '1',
		52391 => '1',
		52392 => '1',
		52393 => '1',
		52394 => '1',
		52395 => '1',
		52396 => '1',
		52397 => '1',
		52398 => '1',
		52399 => '1',
		52400 => '1',
		52401 => '1',
		52402 => '1',
		52403 => '1',
		52404 => '1',
		52405 => '1',
		52406 => '1',
		52407 => '1',
		52408 => '1',
		52409 => '1',
		52410 => '1',
		52411 => '1',
		52412 => '1',
		52413 => '1',
		52414 => '1',
		52415 => '1',
		52416 => '1',
		52417 => '1',
		52418 => '1',
		52419 => '1',
		52420 => '1',
		52421 => '1',
		52422 => '1',
		52423 => '1',
		52424 => '1',
		52425 => '1',
		52426 => '1',
		52427 => '1',
		52428 => '1',
		52429 => '1',
		52430 => '1',
		52431 => '1',
		52432 => '1',
		52433 => '1',
		52434 => '1',
		52435 => '1',
		52436 => '1',
		52437 => '1',
		52438 => '1',
		52439 => '1',
		52440 => '1',
		52441 => '1',
		52442 => '1',
		52443 => '1',
		52444 => '1',
		52445 => '1',
		52446 => '1',
		52447 => '1',
		52448 => '1',
		52449 => '1',
		52450 => '1',
		52451 => '1',
		52452 => '1',
		52453 => '1',
		52454 => '1',
		52455 => '1',
		52456 => '1',
		52457 => '1',
		52458 => '1',
		52459 => '1',
		52460 => '1',
		52461 => '1',
		52462 => '1',
		52463 => '1',
		52464 => '1',
		52465 => '1',
		52466 => '1',
		52467 => '1',
		52468 => '1',
		52469 => '1',
		52470 => '1',
		52471 => '1',
		52472 => '1',
		52473 => '1',
		52474 => '1',
		52475 => '1',
		52476 => '1',
		52477 => '1',
		52478 => '1',
		52479 => '1',
		52480 => '1',
		52481 => '1',
		52482 => '1',
		52483 => '1',
		52484 => '1',
		52485 => '1',
		52486 => '1',
		52487 => '1',
		52488 => '1',
		52489 => '1',
		52490 => '1',
		52491 => '1',
		52492 => '1',
		52493 => '1',
		52494 => '1',
		52495 => '1',
		52496 => '1',
		52497 => '1',
		52498 => '1',
		52499 => '1',
		52500 => '1',
		52501 => '1',
		52502 => '1',
		52503 => '1',
		52504 => '1',
		52505 => '1',
		52506 => '1',
		52507 => '1',
		52508 => '1',
		52509 => '1',
		52510 => '1',
		52511 => '1',
		52512 => '1',
		52513 => '1',
		52514 => '1',
		52515 => '1',
		52516 => '1',
		52517 => '1',
		52518 => '1',
		52519 => '1',
		52520 => '1',
		52521 => '1',
		52522 => '1',
		52523 => '1',
		52524 => '1',
		52525 => '1',
		52526 => '1',
		52527 => '1',
		52528 => '1',
		52529 => '1',
		52530 => '1',
		52531 => '1',
		52532 => '1',
		52533 => '1',
		52534 => '1',
		52535 => '1',
		52536 => '1',
		52537 => '1',
		52538 => '1',
		52539 => '1',
		52540 => '1',
		52541 => '1',
		52542 => '1',
		52543 => '1',
		52544 => '1',
		52545 => '1',
		52546 => '1',
		52547 => '1',
		52548 => '1',
		52549 => '1',
		52550 => '1',
		52551 => '1',
		52552 => '1',
		52553 => '1',
		52554 => '1',
		52555 => '1',
		52556 => '1',
		52557 => '1',
		52558 => '1',
		52559 => '1',
		52560 => '1',
		52561 => '1',
		52562 => '1',
		52563 => '1',
		52564 => '1',
		52565 => '1',
		52566 => '1',
		52567 => '1',
		52568 => '1',
		52569 => '1',
		52570 => '1',
		52571 => '1',
		52572 => '1',
		52573 => '1',
		52574 => '1',
		52575 => '1',
		52576 => '1',
		52577 => '1',
		52578 => '1',
		52579 => '1',
		52580 => '1',
		52581 => '1',
		52582 => '1',
		52583 => '1',
		52584 => '1',
		52585 => '1',
		52586 => '1',
		52587 => '1',
		52588 => '1',
		52589 => '1',
		52590 => '1',
		52591 => '1',
		52592 => '1',
		52593 => '1',
		52594 => '1',
		52595 => '1',
		52596 => '1',
		52597 => '1',
		52598 => '1',
		52599 => '1',
		52600 => '1',
		52601 => '1',
		52602 => '1',
		52603 => '1',
		52604 => '1',
		52605 => '1',
		52606 => '1',
		52607 => '1',
		52608 => '1',
		52609 => '1',
		52610 => '1',
		52611 => '1',
		52612 => '1',
		52613 => '1',
		52614 => '1',
		52615 => '1',
		52616 => '1',
		52617 => '1',
		52618 => '1',
		52619 => '1',
		52620 => '1',
		52621 => '1',
		52622 => '1',
		52623 => '1',
		52624 => '1',
		52625 => '1',
		52626 => '1',
		52627 => '1',
		52628 => '1',
		52629 => '1',
		52630 => '1',
		52631 => '1',
		52632 => '1',
		52633 => '1',
		52634 => '1',
		52635 => '1',
		52636 => '1',
		52637 => '1',
		52638 => '1',
		52639 => '1',
		52640 => '1',
		52641 => '1',
		52642 => '1',
		52643 => '1',
		52644 => '1',
		52645 => '1',
		52646 => '1',
		52647 => '1',
		52648 => '1',
		52649 => '1',
		52650 => '1',
		52651 => '1',
		52652 => '1',
		52653 => '1',
		52654 => '1',
		52655 => '1',
		52656 => '1',
		52657 => '1',
		52658 => '1',
		52659 => '1',
		52660 => '1',
		52661 => '1',
		52662 => '1',
		52663 => '1',
		52664 => '1',
		52665 => '1',
		52666 => '1',
		52667 => '1',
		52668 => '1',
		52669 => '1',
		52670 => '1',
		52671 => '1',
		52672 => '1',
		52673 => '1',
		52674 => '1',
		52675 => '1',
		52676 => '1',
		52677 => '1',
		52678 => '1',
		52679 => '1',
		52680 => '1',
		52681 => '1',
		52682 => '1',
		52683 => '1',
		52684 => '1',
		52685 => '1',
		52686 => '1',
		52687 => '1',
		52688 => '1',
		52689 => '1',
		52690 => '1',
		52691 => '1',
		52692 => '1',
		52693 => '1',
		52694 => '1',
		52695 => '1',
		52696 => '1',
		52697 => '1',
		52698 => '1',
		52699 => '1',
		52700 => '1',
		52701 => '1',
		52702 => '1',
		52703 => '1',
		52704 => '1',
		52705 => '1',
		52706 => '1',
		52707 => '1',
		52708 => '1',
		52709 => '1',
		52710 => '1',
		52711 => '1',
		52712 => '1',
		52713 => '1',
		52714 => '1',
		52715 => '1',
		52716 => '1',
		52717 => '1',
		52718 => '1',
		52719 => '1',
		52720 => '1',
		52721 => '1',
		52722 => '1',
		52723 => '1',
		52724 => '1',
		52725 => '1',
		52726 => '1',
		52727 => '1',
		52728 => '1',
		52729 => '1',
		52730 => '1',
		52731 => '1',
		53376 => '1',
		53377 => '1',
		53378 => '1',
		53379 => '1',
		53380 => '1',
		53381 => '1',
		53382 => '1',
		53383 => '1',
		53384 => '1',
		53385 => '1',
		53386 => '1',
		53387 => '1',
		53388 => '1',
		53389 => '1',
		53390 => '1',
		53391 => '1',
		53392 => '1',
		53393 => '1',
		53394 => '1',
		53395 => '1',
		53396 => '1',
		53397 => '1',
		53398 => '1',
		53399 => '1',
		53400 => '1',
		53401 => '1',
		53402 => '1',
		53403 => '1',
		53404 => '1',
		53405 => '1',
		53406 => '1',
		53407 => '1',
		53408 => '1',
		53409 => '1',
		53410 => '1',
		53411 => '1',
		53412 => '1',
		53413 => '1',
		53414 => '1',
		53415 => '1',
		53416 => '1',
		53417 => '1',
		53418 => '1',
		53419 => '1',
		53420 => '1',
		53421 => '1',
		53422 => '1',
		53423 => '1',
		53424 => '1',
		53425 => '1',
		53426 => '1',
		53427 => '1',
		53428 => '1',
		53429 => '1',
		53430 => '1',
		53431 => '1',
		53432 => '1',
		53433 => '1',
		53434 => '1',
		53435 => '1',
		53436 => '1',
		53437 => '1',
		53438 => '1',
		53439 => '1',
		53440 => '1',
		53441 => '1',
		53442 => '1',
		53443 => '1',
		53444 => '1',
		53445 => '1',
		53446 => '1',
		53447 => '1',
		53448 => '1',
		53449 => '1',
		53450 => '1',
		53451 => '1',
		53452 => '1',
		53453 => '1',
		53454 => '1',
		53455 => '1',
		53456 => '1',
		53457 => '1',
		53458 => '1',
		53459 => '1',
		53460 => '1',
		53461 => '1',
		53462 => '1',
		53463 => '1',
		53464 => '1',
		53465 => '1',
		53466 => '1',
		53467 => '1',
		53468 => '1',
		53469 => '1',
		53470 => '1',
		53471 => '1',
		53472 => '1',
		53473 => '1',
		53474 => '1',
		53475 => '1',
		53476 => '1',
		53477 => '1',
		53478 => '1',
		53479 => '1',
		53480 => '1',
		53481 => '1',
		53482 => '1',
		53483 => '1',
		53484 => '1',
		53485 => '1',
		53486 => '1',
		53487 => '1',
		53488 => '1',
		53489 => '1',
		53490 => '1',
		53491 => '1',
		53492 => '1',
		53493 => '1',
		53494 => '1',
		53495 => '1',
		53496 => '1',
		53497 => '1',
		53498 => '1',
		53499 => '1',
		53500 => '1',
		53501 => '1',
		53502 => '1',
		53503 => '1',
		53504 => '1',
		53505 => '1',
		53506 => '1',
		53507 => '1',
		53508 => '1',
		53509 => '1',
		53510 => '1',
		53511 => '1',
		53512 => '1',
		53513 => '1',
		53514 => '1',
		53515 => '1',
		53516 => '1',
		53517 => '1',
		53518 => '1',
		53519 => '1',
		53520 => '1',
		53521 => '1',
		53522 => '1',
		53523 => '1',
		53524 => '1',
		53525 => '1',
		53526 => '1',
		53527 => '1',
		53528 => '1',
		53529 => '1',
		53530 => '1',
		53531 => '1',
		53532 => '1',
		53533 => '1',
		53534 => '1',
		53535 => '1',
		53536 => '1',
		53537 => '1',
		53538 => '1',
		53539 => '1',
		53540 => '1',
		53541 => '1',
		53542 => '1',
		53543 => '1',
		53544 => '1',
		53545 => '1',
		53546 => '1',
		53547 => '1',
		53548 => '1',
		53549 => '1',
		53550 => '1',
		53551 => '1',
		53552 => '1',
		53553 => '1',
		53554 => '1',
		53555 => '1',
		53556 => '1',
		53557 => '1',
		53558 => '1',
		53559 => '1',
		53560 => '1',
		53561 => '1',
		53562 => '1',
		53563 => '1',
		53564 => '1',
		53565 => '1',
		53566 => '1',
		53567 => '1',
		53568 => '1',
		53569 => '1',
		53570 => '1',
		53571 => '1',
		53572 => '1',
		53573 => '1',
		53574 => '1',
		53575 => '1',
		53576 => '1',
		53577 => '1',
		53578 => '1',
		53579 => '1',
		53580 => '1',
		53581 => '1',
		53582 => '1',
		53583 => '1',
		53584 => '1',
		53585 => '1',
		53586 => '1',
		53587 => '1',
		53588 => '1',
		53589 => '1',
		53590 => '1',
		53591 => '1',
		53592 => '1',
		53593 => '1',
		53594 => '1',
		53595 => '1',
		53596 => '1',
		53597 => '1',
		53598 => '1',
		53599 => '1',
		53600 => '1',
		53601 => '1',
		53602 => '1',
		53603 => '1',
		53604 => '1',
		53605 => '1',
		53606 => '1',
		53607 => '1',
		53608 => '1',
		53609 => '1',
		53610 => '1',
		53611 => '1',
		53612 => '1',
		53613 => '1',
		53614 => '1',
		53615 => '1',
		53616 => '1',
		53617 => '1',
		53618 => '1',
		53619 => '1',
		53620 => '1',
		53621 => '1',
		53622 => '1',
		53623 => '1',
		53624 => '1',
		53625 => '1',
		53626 => '1',
		53627 => '1',
		53628 => '1',
		53629 => '1',
		53630 => '1',
		53631 => '1',
		53632 => '1',
		53633 => '1',
		53634 => '1',
		53635 => '1',
		53636 => '1',
		53637 => '1',
		53638 => '1',
		53639 => '1',
		53640 => '1',
		53641 => '1',
		53642 => '1',
		53643 => '1',
		53644 => '1',
		53645 => '1',
		53646 => '1',
		53647 => '1',
		53648 => '1',
		53649 => '1',
		53650 => '1',
		53651 => '1',
		53652 => '1',
		53653 => '1',
		53654 => '1',
		53655 => '1',
		53656 => '1',
		53657 => '1',
		53658 => '1',
		53659 => '1',
		53660 => '1',
		53661 => '1',
		53662 => '1',
		53663 => '1',
		53664 => '1',
		53665 => '1',
		53666 => '1',
		53667 => '1',
		53668 => '1',
		53669 => '1',
		53670 => '1',
		53671 => '1',
		53672 => '1',
		53673 => '1',
		53674 => '1',
		53675 => '1',
		53676 => '1',
		53677 => '1',
		53678 => '1',
		53679 => '1',
		53680 => '1',
		53681 => '1',
		53682 => '1',
		53683 => '1',
		53684 => '1',
		53685 => '1',
		53686 => '1',
		53687 => '1',
		53688 => '1',
		53689 => '1',
		53690 => '1',
		53691 => '1',
		53692 => '1',
		53693 => '1',
		53694 => '1',
		53695 => '1',
		53696 => '1',
		53697 => '1',
		53698 => '1',
		53699 => '1',
		53700 => '1',
		53701 => '1',
		53702 => '1',
		53703 => '1',
		53704 => '1',
		53705 => '1',
		53706 => '1',
		53707 => '1',
		53708 => '1',
		53709 => '1',
		53710 => '1',
		53711 => '1',
		53712 => '1',
		53713 => '1',
		53714 => '1',
		53715 => '1',
		53716 => '1',
		53717 => '1',
		53718 => '1',
		53719 => '1',
		53720 => '1',
		53721 => '1',
		53722 => '1',
		53723 => '1',
		53724 => '1',
		53725 => '1',
		53726 => '1',
		53727 => '1',
		53728 => '1',
		53729 => '1',
		53730 => '1',
		53731 => '1',
		53732 => '1',
		53733 => '1',
		53734 => '1',
		53735 => '1',
		53736 => '1',
		53737 => '1',
		53738 => '1',
		53739 => '1',
		53740 => '1',
		53741 => '1',
		53742 => '1',
		53743 => '1',
		53744 => '1',
		53745 => '1',
		53746 => '1',
		53747 => '1',
		53748 => '1',
		53749 => '1',
		53750 => '1',
		53751 => '1',
		53752 => '1',
		53753 => '1',
		53754 => '1',
		53755 => '1',
		54400 => '1',
		54401 => '1',
		54402 => '1',
		54403 => '1',
		54404 => '1',
		54525 => '1',
		54526 => '1',
		54527 => '1',
		54528 => '1',
		54529 => '1',
		54650 => '1',
		54651 => '1',
		54652 => '1',
		54653 => '1',
		54654 => '1',
		54775 => '1',
		54776 => '1',
		54777 => '1',
		54778 => '1',
		54779 => '1',
		55424 => '1',
		55425 => '1',
		55426 => '1',
		55427 => '1',
		55428 => '1',
		55549 => '1',
		55550 => '1',
		55551 => '1',
		55552 => '1',
		55553 => '1',
		55674 => '1',
		55675 => '1',
		55676 => '1',
		55677 => '1',
		55678 => '1',
		55799 => '1',
		55800 => '1',
		55801 => '1',
		55802 => '1',
		55803 => '1',
		56448 => '1',
		56449 => '1',
		56450 => '1',
		56451 => '1',
		56452 => '1',
		56573 => '1',
		56574 => '1',
		56575 => '1',
		56576 => '1',
		56577 => '1',
		56698 => '1',
		56699 => '1',
		56700 => '1',
		56701 => '1',
		56702 => '1',
		56823 => '1',
		56824 => '1',
		56825 => '1',
		56826 => '1',
		56827 => '1',
		57472 => '1',
		57473 => '1',
		57474 => '1',
		57475 => '1',
		57476 => '1',
		57597 => '1',
		57598 => '1',
		57599 => '1',
		57600 => '1',
		57601 => '1',
		57722 => '1',
		57723 => '1',
		57724 => '1',
		57725 => '1',
		57726 => '1',
		57847 => '1',
		57848 => '1',
		57849 => '1',
		57850 => '1',
		57851 => '1',
		58496 => '1',
		58497 => '1',
		58498 => '1',
		58499 => '1',
		58500 => '1',
		58621 => '1',
		58622 => '1',
		58623 => '1',
		58624 => '1',
		58625 => '1',
		58746 => '1',
		58747 => '1',
		58748 => '1',
		58749 => '1',
		58750 => '1',
		58871 => '1',
		58872 => '1',
		58873 => '1',
		58874 => '1',
		58875 => '1',
		59520 => '1',
		59521 => '1',
		59522 => '1',
		59523 => '1',
		59524 => '1',
		59645 => '1',
		59646 => '1',
		59647 => '1',
		59648 => '1',
		59649 => '1',
		59770 => '1',
		59771 => '1',
		59772 => '1',
		59773 => '1',
		59774 => '1',
		59895 => '1',
		59896 => '1',
		59897 => '1',
		59898 => '1',
		59899 => '1',
		60544 => '1',
		60545 => '1',
		60546 => '1',
		60547 => '1',
		60548 => '1',
		60669 => '1',
		60670 => '1',
		60671 => '1',
		60672 => '1',
		60673 => '1',
		60794 => '1',
		60795 => '1',
		60796 => '1',
		60797 => '1',
		60798 => '1',
		60919 => '1',
		60920 => '1',
		60921 => '1',
		60922 => '1',
		60923 => '1',
		61568 => '1',
		61569 => '1',
		61570 => '1',
		61571 => '1',
		61572 => '1',
		61693 => '1',
		61694 => '1',
		61695 => '1',
		61696 => '1',
		61697 => '1',
		61818 => '1',
		61819 => '1',
		61820 => '1',
		61821 => '1',
		61822 => '1',
		61943 => '1',
		61944 => '1',
		61945 => '1',
		61946 => '1',
		61947 => '1',
		62592 => '1',
		62593 => '1',
		62594 => '1',
		62595 => '1',
		62596 => '1',
		62717 => '1',
		62718 => '1',
		62719 => '1',
		62720 => '1',
		62721 => '1',
		62842 => '1',
		62843 => '1',
		62844 => '1',
		62845 => '1',
		62846 => '1',
		62967 => '1',
		62968 => '1',
		62969 => '1',
		62970 => '1',
		62971 => '1',
		63616 => '1',
		63617 => '1',
		63618 => '1',
		63619 => '1',
		63620 => '1',
		63741 => '1',
		63742 => '1',
		63743 => '1',
		63744 => '1',
		63745 => '1',
		63866 => '1',
		63867 => '1',
		63868 => '1',
		63869 => '1',
		63870 => '1',
		63991 => '1',
		63992 => '1',
		63993 => '1',
		63994 => '1',
		63995 => '1',
		64640 => '1',
		64641 => '1',
		64642 => '1',
		64643 => '1',
		64644 => '1',
		64765 => '1',
		64766 => '1',
		64767 => '1',
		64768 => '1',
		64769 => '1',
		64890 => '1',
		64891 => '1',
		64892 => '1',
		64893 => '1',
		64894 => '1',
		65015 => '1',
		65016 => '1',
		65017 => '1',
		65018 => '1',
		65019 => '1',
		65664 => '1',
		65665 => '1',
		65666 => '1',
		65667 => '1',
		65668 => '1',
		65789 => '1',
		65790 => '1',
		65791 => '1',
		65792 => '1',
		65793 => '1',
		65914 => '1',
		65915 => '1',
		65916 => '1',
		65917 => '1',
		65918 => '1',
		66039 => '1',
		66040 => '1',
		66041 => '1',
		66042 => '1',
		66043 => '1',
		66688 => '1',
		66689 => '1',
		66690 => '1',
		66691 => '1',
		66692 => '1',
		66813 => '1',
		66814 => '1',
		66815 => '1',
		66816 => '1',
		66817 => '1',
		66938 => '1',
		66939 => '1',
		66940 => '1',
		66941 => '1',
		66942 => '1',
		67063 => '1',
		67064 => '1',
		67065 => '1',
		67066 => '1',
		67067 => '1',
		67712 => '1',
		67713 => '1',
		67714 => '1',
		67715 => '1',
		67716 => '1',
		67837 => '1',
		67838 => '1',
		67839 => '1',
		67840 => '1',
		67841 => '1',
		67962 => '1',
		67963 => '1',
		67964 => '1',
		67965 => '1',
		67966 => '1',
		68087 => '1',
		68088 => '1',
		68089 => '1',
		68090 => '1',
		68091 => '1',
		68736 => '1',
		68737 => '1',
		68738 => '1',
		68739 => '1',
		68740 => '1',
		68861 => '1',
		68862 => '1',
		68863 => '1',
		68864 => '1',
		68865 => '1',
		68986 => '1',
		68987 => '1',
		68988 => '1',
		68989 => '1',
		68990 => '1',
		69111 => '1',
		69112 => '1',
		69113 => '1',
		69114 => '1',
		69115 => '1',
		69760 => '1',
		69761 => '1',
		69762 => '1',
		69763 => '1',
		69764 => '1',
		69885 => '1',
		69886 => '1',
		69887 => '1',
		69888 => '1',
		69889 => '1',
		70010 => '1',
		70011 => '1',
		70012 => '1',
		70013 => '1',
		70014 => '1',
		70135 => '1',
		70136 => '1',
		70137 => '1',
		70138 => '1',
		70139 => '1',
		70784 => '1',
		70785 => '1',
		70786 => '1',
		70787 => '1',
		70788 => '1',
		70909 => '1',
		70910 => '1',
		70911 => '1',
		70912 => '1',
		70913 => '1',
		71034 => '1',
		71035 => '1',
		71036 => '1',
		71037 => '1',
		71038 => '1',
		71159 => '1',
		71160 => '1',
		71161 => '1',
		71162 => '1',
		71163 => '1',
		71808 => '1',
		71809 => '1',
		71810 => '1',
		71811 => '1',
		71812 => '1',
		71933 => '1',
		71934 => '1',
		71935 => '1',
		71936 => '1',
		71937 => '1',
		72058 => '1',
		72059 => '1',
		72060 => '1',
		72061 => '1',
		72062 => '1',
		72183 => '1',
		72184 => '1',
		72185 => '1',
		72186 => '1',
		72187 => '1',
		72832 => '1',
		72833 => '1',
		72834 => '1',
		72835 => '1',
		72836 => '1',
		72957 => '1',
		72958 => '1',
		72959 => '1',
		72960 => '1',
		72961 => '1',
		73082 => '1',
		73083 => '1',
		73084 => '1',
		73085 => '1',
		73086 => '1',
		73207 => '1',
		73208 => '1',
		73209 => '1',
		73210 => '1',
		73211 => '1',
		73856 => '1',
		73857 => '1',
		73858 => '1',
		73859 => '1',
		73860 => '1',
		73981 => '1',
		73982 => '1',
		73983 => '1',
		73984 => '1',
		73985 => '1',
		74106 => '1',
		74107 => '1',
		74108 => '1',
		74109 => '1',
		74110 => '1',
		74231 => '1',
		74232 => '1',
		74233 => '1',
		74234 => '1',
		74235 => '1',
		74880 => '1',
		74881 => '1',
		74882 => '1',
		74883 => '1',
		74884 => '1',
		75005 => '1',
		75006 => '1',
		75007 => '1',
		75008 => '1',
		75009 => '1',
		75130 => '1',
		75131 => '1',
		75132 => '1',
		75133 => '1',
		75134 => '1',
		75255 => '1',
		75256 => '1',
		75257 => '1',
		75258 => '1',
		75259 => '1',
		75904 => '1',
		75905 => '1',
		75906 => '1',
		75907 => '1',
		75908 => '1',
		76029 => '1',
		76030 => '1',
		76031 => '1',
		76032 => '1',
		76033 => '1',
		76154 => '1',
		76155 => '1',
		76156 => '1',
		76157 => '1',
		76158 => '1',
		76279 => '1',
		76280 => '1',
		76281 => '1',
		76282 => '1',
		76283 => '1',
		76928 => '1',
		76929 => '1',
		76930 => '1',
		76931 => '1',
		76932 => '1',
		77053 => '1',
		77054 => '1',
		77055 => '1',
		77056 => '1',
		77057 => '1',
		77178 => '1',
		77179 => '1',
		77180 => '1',
		77181 => '1',
		77182 => '1',
		77303 => '1',
		77304 => '1',
		77305 => '1',
		77306 => '1',
		77307 => '1',
		77952 => '1',
		77953 => '1',
		77954 => '1',
		77955 => '1',
		77956 => '1',
		78077 => '1',
		78078 => '1',
		78079 => '1',
		78080 => '1',
		78081 => '1',
		78202 => '1',
		78203 => '1',
		78204 => '1',
		78205 => '1',
		78206 => '1',
		78327 => '1',
		78328 => '1',
		78329 => '1',
		78330 => '1',
		78331 => '1',
		78976 => '1',
		78977 => '1',
		78978 => '1',
		78979 => '1',
		78980 => '1',
		79101 => '1',
		79102 => '1',
		79103 => '1',
		79104 => '1',
		79105 => '1',
		79226 => '1',
		79227 => '1',
		79228 => '1',
		79229 => '1',
		79230 => '1',
		79351 => '1',
		79352 => '1',
		79353 => '1',
		79354 => '1',
		79355 => '1',
		80000 => '1',
		80001 => '1',
		80002 => '1',
		80003 => '1',
		80004 => '1',
		80125 => '1',
		80126 => '1',
		80127 => '1',
		80128 => '1',
		80129 => '1',
		80250 => '1',
		80251 => '1',
		80252 => '1',
		80253 => '1',
		80254 => '1',
		80375 => '1',
		80376 => '1',
		80377 => '1',
		80378 => '1',
		80379 => '1',
		81024 => '1',
		81025 => '1',
		81026 => '1',
		81027 => '1',
		81028 => '1',
		81149 => '1',
		81150 => '1',
		81151 => '1',
		81152 => '1',
		81153 => '1',
		81274 => '1',
		81275 => '1',
		81276 => '1',
		81277 => '1',
		81278 => '1',
		81399 => '1',
		81400 => '1',
		81401 => '1',
		81402 => '1',
		81403 => '1',
		82048 => '1',
		82049 => '1',
		82050 => '1',
		82051 => '1',
		82052 => '1',
		82173 => '1',
		82174 => '1',
		82175 => '1',
		82176 => '1',
		82177 => '1',
		82298 => '1',
		82299 => '1',
		82300 => '1',
		82301 => '1',
		82302 => '1',
		82423 => '1',
		82424 => '1',
		82425 => '1',
		82426 => '1',
		82427 => '1',
		83072 => '1',
		83073 => '1',
		83074 => '1',
		83075 => '1',
		83076 => '1',
		83197 => '1',
		83198 => '1',
		83199 => '1',
		83200 => '1',
		83201 => '1',
		83322 => '1',
		83323 => '1',
		83324 => '1',
		83325 => '1',
		83326 => '1',
		83447 => '1',
		83448 => '1',
		83449 => '1',
		83450 => '1',
		83451 => '1',
		84096 => '1',
		84097 => '1',
		84098 => '1',
		84099 => '1',
		84100 => '1',
		84221 => '1',
		84222 => '1',
		84223 => '1',
		84224 => '1',
		84225 => '1',
		84346 => '1',
		84347 => '1',
		84348 => '1',
		84349 => '1',
		84350 => '1',
		84471 => '1',
		84472 => '1',
		84473 => '1',
		84474 => '1',
		84475 => '1',
		85120 => '1',
		85121 => '1',
		85122 => '1',
		85123 => '1',
		85124 => '1',
		85245 => '1',
		85246 => '1',
		85247 => '1',
		85248 => '1',
		85249 => '1',
		85370 => '1',
		85371 => '1',
		85372 => '1',
		85373 => '1',
		85374 => '1',
		85495 => '1',
		85496 => '1',
		85497 => '1',
		85498 => '1',
		85499 => '1',
		86144 => '1',
		86145 => '1',
		86146 => '1',
		86147 => '1',
		86148 => '1',
		86269 => '1',
		86270 => '1',
		86271 => '1',
		86272 => '1',
		86273 => '1',
		86394 => '1',
		86395 => '1',
		86396 => '1',
		86397 => '1',
		86398 => '1',
		86519 => '1',
		86520 => '1',
		86521 => '1',
		86522 => '1',
		86523 => '1',
		87168 => '1',
		87169 => '1',
		87170 => '1',
		87171 => '1',
		87172 => '1',
		87293 => '1',
		87294 => '1',
		87295 => '1',
		87296 => '1',
		87297 => '1',
		87418 => '1',
		87419 => '1',
		87420 => '1',
		87421 => '1',
		87422 => '1',
		87543 => '1',
		87544 => '1',
		87545 => '1',
		87546 => '1',
		87547 => '1',
		88192 => '1',
		88193 => '1',
		88194 => '1',
		88195 => '1',
		88196 => '1',
		88317 => '1',
		88318 => '1',
		88319 => '1',
		88320 => '1',
		88321 => '1',
		88442 => '1',
		88443 => '1',
		88444 => '1',
		88445 => '1',
		88446 => '1',
		88567 => '1',
		88568 => '1',
		88569 => '1',
		88570 => '1',
		88571 => '1',
		89216 => '1',
		89217 => '1',
		89218 => '1',
		89219 => '1',
		89220 => '1',
		89341 => '1',
		89342 => '1',
		89343 => '1',
		89344 => '1',
		89345 => '1',
		89466 => '1',
		89467 => '1',
		89468 => '1',
		89469 => '1',
		89470 => '1',
		89591 => '1',
		89592 => '1',
		89593 => '1',
		89594 => '1',
		89595 => '1',
		90240 => '1',
		90241 => '1',
		90242 => '1',
		90243 => '1',
		90244 => '1',
		90365 => '1',
		90366 => '1',
		90367 => '1',
		90368 => '1',
		90369 => '1',
		90490 => '1',
		90491 => '1',
		90492 => '1',
		90493 => '1',
		90494 => '1',
		90615 => '1',
		90616 => '1',
		90617 => '1',
		90618 => '1',
		90619 => '1',
		91264 => '1',
		91265 => '1',
		91266 => '1',
		91267 => '1',
		91268 => '1',
		91389 => '1',
		91390 => '1',
		91391 => '1',
		91392 => '1',
		91393 => '1',
		91514 => '1',
		91515 => '1',
		91516 => '1',
		91517 => '1',
		91518 => '1',
		91639 => '1',
		91640 => '1',
		91641 => '1',
		91642 => '1',
		91643 => '1',
		92288 => '1',
		92289 => '1',
		92290 => '1',
		92291 => '1',
		92292 => '1',
		92413 => '1',
		92414 => '1',
		92415 => '1',
		92416 => '1',
		92417 => '1',
		92538 => '1',
		92539 => '1',
		92540 => '1',
		92541 => '1',
		92542 => '1',
		92663 => '1',
		92664 => '1',
		92665 => '1',
		92666 => '1',
		92667 => '1',
		93312 => '1',
		93313 => '1',
		93314 => '1',
		93315 => '1',
		93316 => '1',
		93437 => '1',
		93438 => '1',
		93439 => '1',
		93440 => '1',
		93441 => '1',
		93562 => '1',
		93563 => '1',
		93564 => '1',
		93565 => '1',
		93566 => '1',
		93687 => '1',
		93688 => '1',
		93689 => '1',
		93690 => '1',
		93691 => '1',
		94336 => '1',
		94337 => '1',
		94338 => '1',
		94339 => '1',
		94340 => '1',
		94461 => '1',
		94462 => '1',
		94463 => '1',
		94464 => '1',
		94465 => '1',
		94586 => '1',
		94587 => '1',
		94588 => '1',
		94589 => '1',
		94590 => '1',
		94711 => '1',
		94712 => '1',
		94713 => '1',
		94714 => '1',
		94715 => '1',
		95360 => '1',
		95361 => '1',
		95362 => '1',
		95363 => '1',
		95364 => '1',
		95485 => '1',
		95486 => '1',
		95487 => '1',
		95488 => '1',
		95489 => '1',
		95610 => '1',
		95611 => '1',
		95612 => '1',
		95613 => '1',
		95614 => '1',
		95735 => '1',
		95736 => '1',
		95737 => '1',
		95738 => '1',
		95739 => '1',
		96384 => '1',
		96385 => '1',
		96386 => '1',
		96387 => '1',
		96388 => '1',
		96509 => '1',
		96510 => '1',
		96511 => '1',
		96512 => '1',
		96513 => '1',
		96634 => '1',
		96635 => '1',
		96636 => '1',
		96637 => '1',
		96638 => '1',
		96759 => '1',
		96760 => '1',
		96761 => '1',
		96762 => '1',
		96763 => '1',
		97408 => '1',
		97409 => '1',
		97410 => '1',
		97411 => '1',
		97412 => '1',
		97533 => '1',
		97534 => '1',
		97535 => '1',
		97536 => '1',
		97537 => '1',
		97658 => '1',
		97659 => '1',
		97660 => '1',
		97661 => '1',
		97662 => '1',
		97783 => '1',
		97784 => '1',
		97785 => '1',
		97786 => '1',
		97787 => '1',
		98432 => '1',
		98433 => '1',
		98434 => '1',
		98435 => '1',
		98436 => '1',
		98557 => '1',
		98558 => '1',
		98559 => '1',
		98560 => '1',
		98561 => '1',
		98682 => '1',
		98683 => '1',
		98684 => '1',
		98685 => '1',
		98686 => '1',
		98807 => '1',
		98808 => '1',
		98809 => '1',
		98810 => '1',
		98811 => '1',
		99456 => '1',
		99457 => '1',
		99458 => '1',
		99459 => '1',
		99460 => '1',
		99581 => '1',
		99582 => '1',
		99583 => '1',
		99584 => '1',
		99585 => '1',
		99706 => '1',
		99707 => '1',
		99708 => '1',
		99709 => '1',
		99710 => '1',
		99831 => '1',
		99832 => '1',
		99833 => '1',
		99834 => '1',
		99835 => '1',
		100480 => '1',
		100481 => '1',
		100482 => '1',
		100483 => '1',
		100484 => '1',
		100605 => '1',
		100606 => '1',
		100607 => '1',
		100608 => '1',
		100609 => '1',
		100730 => '1',
		100731 => '1',
		100732 => '1',
		100733 => '1',
		100734 => '1',
		100855 => '1',
		100856 => '1',
		100857 => '1',
		100858 => '1',
		100859 => '1',
		101504 => '1',
		101505 => '1',
		101506 => '1',
		101507 => '1',
		101508 => '1',
		101629 => '1',
		101630 => '1',
		101631 => '1',
		101632 => '1',
		101633 => '1',
		101754 => '1',
		101755 => '1',
		101756 => '1',
		101757 => '1',
		101758 => '1',
		101879 => '1',
		101880 => '1',
		101881 => '1',
		101882 => '1',
		101883 => '1',
		102528 => '1',
		102529 => '1',
		102530 => '1',
		102531 => '1',
		102532 => '1',
		102653 => '1',
		102654 => '1',
		102655 => '1',
		102656 => '1',
		102657 => '1',
		102778 => '1',
		102779 => '1',
		102780 => '1',
		102781 => '1',
		102782 => '1',
		102903 => '1',
		102904 => '1',
		102905 => '1',
		102906 => '1',
		102907 => '1',
		103552 => '1',
		103553 => '1',
		103554 => '1',
		103555 => '1',
		103556 => '1',
		103677 => '1',
		103678 => '1',
		103679 => '1',
		103680 => '1',
		103681 => '1',
		103802 => '1',
		103803 => '1',
		103804 => '1',
		103805 => '1',
		103806 => '1',
		103927 => '1',
		103928 => '1',
		103929 => '1',
		103930 => '1',
		103931 => '1',
		104576 => '1',
		104577 => '1',
		104578 => '1',
		104579 => '1',
		104580 => '1',
		104701 => '1',
		104702 => '1',
		104703 => '1',
		104704 => '1',
		104705 => '1',
		104826 => '1',
		104827 => '1',
		104828 => '1',
		104829 => '1',
		104830 => '1',
		104951 => '1',
		104952 => '1',
		104953 => '1',
		104954 => '1',
		104955 => '1',
		105600 => '1',
		105601 => '1',
		105602 => '1',
		105603 => '1',
		105604 => '1',
		105725 => '1',
		105726 => '1',
		105727 => '1',
		105728 => '1',
		105729 => '1',
		105850 => '1',
		105851 => '1',
		105852 => '1',
		105853 => '1',
		105854 => '1',
		105975 => '1',
		105976 => '1',
		105977 => '1',
		105978 => '1',
		105979 => '1',
		106624 => '1',
		106625 => '1',
		106626 => '1',
		106627 => '1',
		106628 => '1',
		106749 => '1',
		106750 => '1',
		106751 => '1',
		106752 => '1',
		106753 => '1',
		106874 => '1',
		106875 => '1',
		106876 => '1',
		106877 => '1',
		106878 => '1',
		106999 => '1',
		107000 => '1',
		107001 => '1',
		107002 => '1',
		107003 => '1',
		107648 => '1',
		107649 => '1',
		107650 => '1',
		107651 => '1',
		107652 => '1',
		107773 => '1',
		107774 => '1',
		107775 => '1',
		107776 => '1',
		107777 => '1',
		107898 => '1',
		107899 => '1',
		107900 => '1',
		107901 => '1',
		107902 => '1',
		108023 => '1',
		108024 => '1',
		108025 => '1',
		108026 => '1',
		108027 => '1',
		108672 => '1',
		108673 => '1',
		108674 => '1',
		108675 => '1',
		108676 => '1',
		108797 => '1',
		108798 => '1',
		108799 => '1',
		108800 => '1',
		108801 => '1',
		108922 => '1',
		108923 => '1',
		108924 => '1',
		108925 => '1',
		108926 => '1',
		109047 => '1',
		109048 => '1',
		109049 => '1',
		109050 => '1',
		109051 => '1',
		109696 => '1',
		109697 => '1',
		109698 => '1',
		109699 => '1',
		109700 => '1',
		109821 => '1',
		109822 => '1',
		109823 => '1',
		109824 => '1',
		109825 => '1',
		109946 => '1',
		109947 => '1',
		109948 => '1',
		109949 => '1',
		109950 => '1',
		110071 => '1',
		110072 => '1',
		110073 => '1',
		110074 => '1',
		110075 => '1',
		110720 => '1',
		110721 => '1',
		110722 => '1',
		110723 => '1',
		110724 => '1',
		110845 => '1',
		110846 => '1',
		110847 => '1',
		110848 => '1',
		110849 => '1',
		110970 => '1',
		110971 => '1',
		110972 => '1',
		110973 => '1',
		110974 => '1',
		111095 => '1',
		111096 => '1',
		111097 => '1',
		111098 => '1',
		111099 => '1',
		111744 => '1',
		111745 => '1',
		111746 => '1',
		111747 => '1',
		111748 => '1',
		111869 => '1',
		111870 => '1',
		111871 => '1',
		111872 => '1',
		111873 => '1',
		111994 => '1',
		111995 => '1',
		111996 => '1',
		111997 => '1',
		111998 => '1',
		112119 => '1',
		112120 => '1',
		112121 => '1',
		112122 => '1',
		112123 => '1',
		112768 => '1',
		112769 => '1',
		112770 => '1',
		112771 => '1',
		112772 => '1',
		112893 => '1',
		112894 => '1',
		112895 => '1',
		112896 => '1',
		112897 => '1',
		113018 => '1',
		113019 => '1',
		113020 => '1',
		113021 => '1',
		113022 => '1',
		113143 => '1',
		113144 => '1',
		113145 => '1',
		113146 => '1',
		113147 => '1',
		113792 => '1',
		113793 => '1',
		113794 => '1',
		113795 => '1',
		113796 => '1',
		113917 => '1',
		113918 => '1',
		113919 => '1',
		113920 => '1',
		113921 => '1',
		114042 => '1',
		114043 => '1',
		114044 => '1',
		114045 => '1',
		114046 => '1',
		114167 => '1',
		114168 => '1',
		114169 => '1',
		114170 => '1',
		114171 => '1',
		114816 => '1',
		114817 => '1',
		114818 => '1',
		114819 => '1',
		114820 => '1',
		114941 => '1',
		114942 => '1',
		114943 => '1',
		114944 => '1',
		114945 => '1',
		115066 => '1',
		115067 => '1',
		115068 => '1',
		115069 => '1',
		115070 => '1',
		115191 => '1',
		115192 => '1',
		115193 => '1',
		115194 => '1',
		115195 => '1',
		115840 => '1',
		115841 => '1',
		115842 => '1',
		115843 => '1',
		115844 => '1',
		115965 => '1',
		115966 => '1',
		115967 => '1',
		115968 => '1',
		115969 => '1',
		116090 => '1',
		116091 => '1',
		116092 => '1',
		116093 => '1',
		116094 => '1',
		116215 => '1',
		116216 => '1',
		116217 => '1',
		116218 => '1',
		116219 => '1',
		116864 => '1',
		116865 => '1',
		116866 => '1',
		116867 => '1',
		116868 => '1',
		116989 => '1',
		116990 => '1',
		116991 => '1',
		116992 => '1',
		116993 => '1',
		117114 => '1',
		117115 => '1',
		117116 => '1',
		117117 => '1',
		117118 => '1',
		117239 => '1',
		117240 => '1',
		117241 => '1',
		117242 => '1',
		117243 => '1',
		117888 => '1',
		117889 => '1',
		117890 => '1',
		117891 => '1',
		117892 => '1',
		118013 => '1',
		118014 => '1',
		118015 => '1',
		118016 => '1',
		118017 => '1',
		118138 => '1',
		118139 => '1',
		118140 => '1',
		118141 => '1',
		118142 => '1',
		118263 => '1',
		118264 => '1',
		118265 => '1',
		118266 => '1',
		118267 => '1',
		118912 => '1',
		118913 => '1',
		118914 => '1',
		118915 => '1',
		118916 => '1',
		119037 => '1',
		119038 => '1',
		119039 => '1',
		119040 => '1',
		119041 => '1',
		119162 => '1',
		119163 => '1',
		119164 => '1',
		119165 => '1',
		119166 => '1',
		119287 => '1',
		119288 => '1',
		119289 => '1',
		119290 => '1',
		119291 => '1',
		119936 => '1',
		119937 => '1',
		119938 => '1',
		119939 => '1',
		119940 => '1',
		120061 => '1',
		120062 => '1',
		120063 => '1',
		120064 => '1',
		120065 => '1',
		120186 => '1',
		120187 => '1',
		120188 => '1',
		120189 => '1',
		120190 => '1',
		120311 => '1',
		120312 => '1',
		120313 => '1',
		120314 => '1',
		120315 => '1',
		120960 => '1',
		120961 => '1',
		120962 => '1',
		120963 => '1',
		120964 => '1',
		121085 => '1',
		121086 => '1',
		121087 => '1',
		121088 => '1',
		121089 => '1',
		121210 => '1',
		121211 => '1',
		121212 => '1',
		121213 => '1',
		121214 => '1',
		121335 => '1',
		121336 => '1',
		121337 => '1',
		121338 => '1',
		121339 => '1',
		121984 => '1',
		121985 => '1',
		121986 => '1',
		121987 => '1',
		121988 => '1',
		122109 => '1',
		122110 => '1',
		122111 => '1',
		122112 => '1',
		122113 => '1',
		122234 => '1',
		122235 => '1',
		122236 => '1',
		122237 => '1',
		122238 => '1',
		122359 => '1',
		122360 => '1',
		122361 => '1',
		122362 => '1',
		122363 => '1',
		123008 => '1',
		123009 => '1',
		123010 => '1',
		123011 => '1',
		123012 => '1',
		123133 => '1',
		123134 => '1',
		123135 => '1',
		123136 => '1',
		123137 => '1',
		123258 => '1',
		123259 => '1',
		123260 => '1',
		123261 => '1',
		123262 => '1',
		123383 => '1',
		123384 => '1',
		123385 => '1',
		123386 => '1',
		123387 => '1',
		124032 => '1',
		124033 => '1',
		124034 => '1',
		124035 => '1',
		124036 => '1',
		124157 => '1',
		124158 => '1',
		124159 => '1',
		124160 => '1',
		124161 => '1',
		124282 => '1',
		124283 => '1',
		124284 => '1',
		124285 => '1',
		124286 => '1',
		124407 => '1',
		124408 => '1',
		124409 => '1',
		124410 => '1',
		124411 => '1',
		125056 => '1',
		125057 => '1',
		125058 => '1',
		125059 => '1',
		125060 => '1',
		125181 => '1',
		125182 => '1',
		125183 => '1',
		125184 => '1',
		125185 => '1',
		125306 => '1',
		125307 => '1',
		125308 => '1',
		125309 => '1',
		125310 => '1',
		125431 => '1',
		125432 => '1',
		125433 => '1',
		125434 => '1',
		125435 => '1',
		126080 => '1',
		126081 => '1',
		126082 => '1',
		126083 => '1',
		126084 => '1',
		126205 => '1',
		126206 => '1',
		126207 => '1',
		126208 => '1',
		126209 => '1',
		126330 => '1',
		126331 => '1',
		126332 => '1',
		126333 => '1',
		126334 => '1',
		126455 => '1',
		126456 => '1',
		126457 => '1',
		126458 => '1',
		126459 => '1',
		127104 => '1',
		127105 => '1',
		127106 => '1',
		127107 => '1',
		127108 => '1',
		127229 => '1',
		127230 => '1',
		127231 => '1',
		127232 => '1',
		127233 => '1',
		127354 => '1',
		127355 => '1',
		127356 => '1',
		127357 => '1',
		127358 => '1',
		127479 => '1',
		127480 => '1',
		127481 => '1',
		127482 => '1',
		127483 => '1',
		128128 => '1',
		128129 => '1',
		128130 => '1',
		128131 => '1',
		128132 => '1',
		128253 => '1',
		128254 => '1',
		128255 => '1',
		128256 => '1',
		128257 => '1',
		128378 => '1',
		128379 => '1',
		128380 => '1',
		128381 => '1',
		128382 => '1',
		128503 => '1',
		128504 => '1',
		128505 => '1',
		128506 => '1',
		128507 => '1',
		129152 => '1',
		129153 => '1',
		129154 => '1',
		129155 => '1',
		129156 => '1',
		129277 => '1',
		129278 => '1',
		129279 => '1',
		129280 => '1',
		129281 => '1',
		129402 => '1',
		129403 => '1',
		129404 => '1',
		129405 => '1',
		129406 => '1',
		129527 => '1',
		129528 => '1',
		129529 => '1',
		129530 => '1',
		129531 => '1',
		130176 => '1',
		130177 => '1',
		130178 => '1',
		130179 => '1',
		130180 => '1',
		130301 => '1',
		130302 => '1',
		130303 => '1',
		130304 => '1',
		130305 => '1',
		130426 => '1',
		130427 => '1',
		130428 => '1',
		130429 => '1',
		130430 => '1',
		130551 => '1',
		130552 => '1',
		130553 => '1',
		130554 => '1',
		130555 => '1',
		131200 => '1',
		131201 => '1',
		131202 => '1',
		131203 => '1',
		131204 => '1',
		131325 => '1',
		131326 => '1',
		131327 => '1',
		131328 => '1',
		131329 => '1',
		131450 => '1',
		131451 => '1',
		131452 => '1',
		131453 => '1',
		131454 => '1',
		131575 => '1',
		131576 => '1',
		131577 => '1',
		131578 => '1',
		131579 => '1',
		132224 => '1',
		132225 => '1',
		132226 => '1',
		132227 => '1',
		132228 => '1',
		132349 => '1',
		132350 => '1',
		132351 => '1',
		132352 => '1',
		132353 => '1',
		132474 => '1',
		132475 => '1',
		132476 => '1',
		132477 => '1',
		132478 => '1',
		132599 => '1',
		132600 => '1',
		132601 => '1',
		132602 => '1',
		132603 => '1',
		133248 => '1',
		133249 => '1',
		133250 => '1',
		133251 => '1',
		133252 => '1',
		133373 => '1',
		133374 => '1',
		133375 => '1',
		133376 => '1',
		133377 => '1',
		133498 => '1',
		133499 => '1',
		133500 => '1',
		133501 => '1',
		133502 => '1',
		133623 => '1',
		133624 => '1',
		133625 => '1',
		133626 => '1',
		133627 => '1',
		134272 => '1',
		134273 => '1',
		134274 => '1',
		134275 => '1',
		134276 => '1',
		134397 => '1',
		134398 => '1',
		134399 => '1',
		134400 => '1',
		134401 => '1',
		134522 => '1',
		134523 => '1',
		134524 => '1',
		134525 => '1',
		134526 => '1',
		134647 => '1',
		134648 => '1',
		134649 => '1',
		134650 => '1',
		134651 => '1',
		135296 => '1',
		135297 => '1',
		135298 => '1',
		135299 => '1',
		135300 => '1',
		135421 => '1',
		135422 => '1',
		135423 => '1',
		135424 => '1',
		135425 => '1',
		135546 => '1',
		135547 => '1',
		135548 => '1',
		135549 => '1',
		135550 => '1',
		135671 => '1',
		135672 => '1',
		135673 => '1',
		135674 => '1',
		135675 => '1',
		136320 => '1',
		136321 => '1',
		136322 => '1',
		136323 => '1',
		136324 => '1',
		136445 => '1',
		136446 => '1',
		136447 => '1',
		136448 => '1',
		136449 => '1',
		136570 => '1',
		136571 => '1',
		136572 => '1',
		136573 => '1',
		136574 => '1',
		136695 => '1',
		136696 => '1',
		136697 => '1',
		136698 => '1',
		136699 => '1',
		137344 => '1',
		137345 => '1',
		137346 => '1',
		137347 => '1',
		137348 => '1',
		137469 => '1',
		137470 => '1',
		137471 => '1',
		137472 => '1',
		137473 => '1',
		137594 => '1',
		137595 => '1',
		137596 => '1',
		137597 => '1',
		137598 => '1',
		137719 => '1',
		137720 => '1',
		137721 => '1',
		137722 => '1',
		137723 => '1',
		138368 => '1',
		138369 => '1',
		138370 => '1',
		138371 => '1',
		138372 => '1',
		138493 => '1',
		138494 => '1',
		138495 => '1',
		138496 => '1',
		138497 => '1',
		138618 => '1',
		138619 => '1',
		138620 => '1',
		138621 => '1',
		138622 => '1',
		138743 => '1',
		138744 => '1',
		138745 => '1',
		138746 => '1',
		138747 => '1',
		139392 => '1',
		139393 => '1',
		139394 => '1',
		139395 => '1',
		139396 => '1',
		139517 => '1',
		139518 => '1',
		139519 => '1',
		139520 => '1',
		139521 => '1',
		139642 => '1',
		139643 => '1',
		139644 => '1',
		139645 => '1',
		139646 => '1',
		139767 => '1',
		139768 => '1',
		139769 => '1',
		139770 => '1',
		139771 => '1',
		140416 => '1',
		140417 => '1',
		140418 => '1',
		140419 => '1',
		140420 => '1',
		140541 => '1',
		140542 => '1',
		140543 => '1',
		140544 => '1',
		140545 => '1',
		140666 => '1',
		140667 => '1',
		140668 => '1',
		140669 => '1',
		140670 => '1',
		140791 => '1',
		140792 => '1',
		140793 => '1',
		140794 => '1',
		140795 => '1',
		141440 => '1',
		141441 => '1',
		141442 => '1',
		141443 => '1',
		141444 => '1',
		141565 => '1',
		141566 => '1',
		141567 => '1',
		141568 => '1',
		141569 => '1',
		141690 => '1',
		141691 => '1',
		141692 => '1',
		141693 => '1',
		141694 => '1',
		141815 => '1',
		141816 => '1',
		141817 => '1',
		141818 => '1',
		141819 => '1',
		142464 => '1',
		142465 => '1',
		142466 => '1',
		142467 => '1',
		142468 => '1',
		142589 => '1',
		142590 => '1',
		142591 => '1',
		142592 => '1',
		142593 => '1',
		142714 => '1',
		142715 => '1',
		142716 => '1',
		142717 => '1',
		142718 => '1',
		142839 => '1',
		142840 => '1',
		142841 => '1',
		142842 => '1',
		142843 => '1',
		143488 => '1',
		143489 => '1',
		143490 => '1',
		143491 => '1',
		143492 => '1',
		143613 => '1',
		143614 => '1',
		143615 => '1',
		143616 => '1',
		143617 => '1',
		143738 => '1',
		143739 => '1',
		143740 => '1',
		143741 => '1',
		143742 => '1',
		143863 => '1',
		143864 => '1',
		143865 => '1',
		143866 => '1',
		143867 => '1',
		144512 => '1',
		144513 => '1',
		144514 => '1',
		144515 => '1',
		144516 => '1',
		144637 => '1',
		144638 => '1',
		144639 => '1',
		144640 => '1',
		144641 => '1',
		144762 => '1',
		144763 => '1',
		144764 => '1',
		144765 => '1',
		144766 => '1',
		144887 => '1',
		144888 => '1',
		144889 => '1',
		144890 => '1',
		144891 => '1',
		145536 => '1',
		145537 => '1',
		145538 => '1',
		145539 => '1',
		145540 => '1',
		145661 => '1',
		145662 => '1',
		145663 => '1',
		145664 => '1',
		145665 => '1',
		145786 => '1',
		145787 => '1',
		145788 => '1',
		145789 => '1',
		145790 => '1',
		145911 => '1',
		145912 => '1',
		145913 => '1',
		145914 => '1',
		145915 => '1',
		146560 => '1',
		146561 => '1',
		146562 => '1',
		146563 => '1',
		146564 => '1',
		146685 => '1',
		146686 => '1',
		146687 => '1',
		146688 => '1',
		146689 => '1',
		146810 => '1',
		146811 => '1',
		146812 => '1',
		146813 => '1',
		146814 => '1',
		146935 => '1',
		146936 => '1',
		146937 => '1',
		146938 => '1',
		146939 => '1',
		147584 => '1',
		147585 => '1',
		147586 => '1',
		147587 => '1',
		147588 => '1',
		147709 => '1',
		147710 => '1',
		147711 => '1',
		147712 => '1',
		147713 => '1',
		147834 => '1',
		147835 => '1',
		147836 => '1',
		147837 => '1',
		147838 => '1',
		147959 => '1',
		147960 => '1',
		147961 => '1',
		147962 => '1',
		147963 => '1',
		148608 => '1',
		148609 => '1',
		148610 => '1',
		148611 => '1',
		148612 => '1',
		148733 => '1',
		148734 => '1',
		148735 => '1',
		148736 => '1',
		148737 => '1',
		148858 => '1',
		148859 => '1',
		148860 => '1',
		148861 => '1',
		148862 => '1',
		148983 => '1',
		148984 => '1',
		148985 => '1',
		148986 => '1',
		148987 => '1',
		149632 => '1',
		149633 => '1',
		149634 => '1',
		149635 => '1',
		149636 => '1',
		149757 => '1',
		149758 => '1',
		149759 => '1',
		149760 => '1',
		149761 => '1',
		149882 => '1',
		149883 => '1',
		149884 => '1',
		149885 => '1',
		149886 => '1',
		150007 => '1',
		150008 => '1',
		150009 => '1',
		150010 => '1',
		150011 => '1',
		150656 => '1',
		150657 => '1',
		150658 => '1',
		150659 => '1',
		150660 => '1',
		150781 => '1',
		150782 => '1',
		150783 => '1',
		150784 => '1',
		150785 => '1',
		150906 => '1',
		150907 => '1',
		150908 => '1',
		150909 => '1',
		150910 => '1',
		151031 => '1',
		151032 => '1',
		151033 => '1',
		151034 => '1',
		151035 => '1',
		151680 => '1',
		151681 => '1',
		151682 => '1',
		151683 => '1',
		151684 => '1',
		151805 => '1',
		151806 => '1',
		151807 => '1',
		151808 => '1',
		151809 => '1',
		151930 => '1',
		151931 => '1',
		151932 => '1',
		151933 => '1',
		151934 => '1',
		152055 => '1',
		152056 => '1',
		152057 => '1',
		152058 => '1',
		152059 => '1',
		152704 => '1',
		152705 => '1',
		152706 => '1',
		152707 => '1',
		152708 => '1',
		152829 => '1',
		152830 => '1',
		152831 => '1',
		152832 => '1',
		152833 => '1',
		152954 => '1',
		152955 => '1',
		152956 => '1',
		152957 => '1',
		152958 => '1',
		153079 => '1',
		153080 => '1',
		153081 => '1',
		153082 => '1',
		153083 => '1',
		153728 => '1',
		153729 => '1',
		153730 => '1',
		153731 => '1',
		153732 => '1',
		153853 => '1',
		153854 => '1',
		153855 => '1',
		153856 => '1',
		153857 => '1',
		153978 => '1',
		153979 => '1',
		153980 => '1',
		153981 => '1',
		153982 => '1',
		154103 => '1',
		154104 => '1',
		154105 => '1',
		154106 => '1',
		154107 => '1',
		154752 => '1',
		154753 => '1',
		154754 => '1',
		154755 => '1',
		154756 => '1',
		154877 => '1',
		154878 => '1',
		154879 => '1',
		154880 => '1',
		154881 => '1',
		155002 => '1',
		155003 => '1',
		155004 => '1',
		155005 => '1',
		155006 => '1',
		155127 => '1',
		155128 => '1',
		155129 => '1',
		155130 => '1',
		155131 => '1',
		155776 => '1',
		155777 => '1',
		155778 => '1',
		155779 => '1',
		155780 => '1',
		155901 => '1',
		155902 => '1',
		155903 => '1',
		155904 => '1',
		155905 => '1',
		156026 => '1',
		156027 => '1',
		156028 => '1',
		156029 => '1',
		156030 => '1',
		156151 => '1',
		156152 => '1',
		156153 => '1',
		156154 => '1',
		156155 => '1',
		156800 => '1',
		156801 => '1',
		156802 => '1',
		156803 => '1',
		156804 => '1',
		156925 => '1',
		156926 => '1',
		156927 => '1',
		156928 => '1',
		156929 => '1',
		157050 => '1',
		157051 => '1',
		157052 => '1',
		157053 => '1',
		157054 => '1',
		157175 => '1',
		157176 => '1',
		157177 => '1',
		157178 => '1',
		157179 => '1',
		157824 => '1',
		157825 => '1',
		157826 => '1',
		157827 => '1',
		157828 => '1',
		157949 => '1',
		157950 => '1',
		157951 => '1',
		157952 => '1',
		157953 => '1',
		158074 => '1',
		158075 => '1',
		158076 => '1',
		158077 => '1',
		158078 => '1',
		158199 => '1',
		158200 => '1',
		158201 => '1',
		158202 => '1',
		158203 => '1',
		158848 => '1',
		158849 => '1',
		158850 => '1',
		158851 => '1',
		158852 => '1',
		158973 => '1',
		158974 => '1',
		158975 => '1',
		158976 => '1',
		158977 => '1',
		159098 => '1',
		159099 => '1',
		159100 => '1',
		159101 => '1',
		159102 => '1',
		159223 => '1',
		159224 => '1',
		159225 => '1',
		159226 => '1',
		159227 => '1',
		159872 => '1',
		159873 => '1',
		159874 => '1',
		159875 => '1',
		159876 => '1',
		159997 => '1',
		159998 => '1',
		159999 => '1',
		160000 => '1',
		160001 => '1',
		160122 => '1',
		160123 => '1',
		160124 => '1',
		160125 => '1',
		160126 => '1',
		160247 => '1',
		160248 => '1',
		160249 => '1',
		160250 => '1',
		160251 => '1',
		160896 => '1',
		160897 => '1',
		160898 => '1',
		160899 => '1',
		160900 => '1',
		161021 => '1',
		161022 => '1',
		161023 => '1',
		161024 => '1',
		161025 => '1',
		161146 => '1',
		161147 => '1',
		161148 => '1',
		161149 => '1',
		161150 => '1',
		161271 => '1',
		161272 => '1',
		161273 => '1',
		161274 => '1',
		161275 => '1',
		161920 => '1',
		161921 => '1',
		161922 => '1',
		161923 => '1',
		161924 => '1',
		162045 => '1',
		162046 => '1',
		162047 => '1',
		162048 => '1',
		162049 => '1',
		162170 => '1',
		162171 => '1',
		162172 => '1',
		162173 => '1',
		162174 => '1',
		162295 => '1',
		162296 => '1',
		162297 => '1',
		162298 => '1',
		162299 => '1',
		162944 => '1',
		162945 => '1',
		162946 => '1',
		162947 => '1',
		162948 => '1',
		163069 => '1',
		163070 => '1',
		163071 => '1',
		163072 => '1',
		163073 => '1',
		163194 => '1',
		163195 => '1',
		163196 => '1',
		163197 => '1',
		163198 => '1',
		163319 => '1',
		163320 => '1',
		163321 => '1',
		163322 => '1',
		163323 => '1',
		163968 => '1',
		163969 => '1',
		163970 => '1',
		163971 => '1',
		163972 => '1',
		164093 => '1',
		164094 => '1',
		164095 => '1',
		164096 => '1',
		164097 => '1',
		164218 => '1',
		164219 => '1',
		164220 => '1',
		164221 => '1',
		164222 => '1',
		164343 => '1',
		164344 => '1',
		164345 => '1',
		164346 => '1',
		164347 => '1',
		164992 => '1',
		164993 => '1',
		164994 => '1',
		164995 => '1',
		164996 => '1',
		165117 => '1',
		165118 => '1',
		165119 => '1',
		165120 => '1',
		165121 => '1',
		165242 => '1',
		165243 => '1',
		165244 => '1',
		165245 => '1',
		165246 => '1',
		165367 => '1',
		165368 => '1',
		165369 => '1',
		165370 => '1',
		165371 => '1',
		166016 => '1',
		166017 => '1',
		166018 => '1',
		166019 => '1',
		166020 => '1',
		166141 => '1',
		166142 => '1',
		166143 => '1',
		166144 => '1',
		166145 => '1',
		166266 => '1',
		166267 => '1',
		166268 => '1',
		166269 => '1',
		166270 => '1',
		166391 => '1',
		166392 => '1',
		166393 => '1',
		166394 => '1',
		166395 => '1',
		167040 => '1',
		167041 => '1',
		167042 => '1',
		167043 => '1',
		167044 => '1',
		167165 => '1',
		167166 => '1',
		167167 => '1',
		167168 => '1',
		167169 => '1',
		167290 => '1',
		167291 => '1',
		167292 => '1',
		167293 => '1',
		167294 => '1',
		167415 => '1',
		167416 => '1',
		167417 => '1',
		167418 => '1',
		167419 => '1',
		168064 => '1',
		168065 => '1',
		168066 => '1',
		168067 => '1',
		168068 => '1',
		168189 => '1',
		168190 => '1',
		168191 => '1',
		168192 => '1',
		168193 => '1',
		168314 => '1',
		168315 => '1',
		168316 => '1',
		168317 => '1',
		168318 => '1',
		168439 => '1',
		168440 => '1',
		168441 => '1',
		168442 => '1',
		168443 => '1',
		169088 => '1',
		169089 => '1',
		169090 => '1',
		169091 => '1',
		169092 => '1',
		169213 => '1',
		169214 => '1',
		169215 => '1',
		169216 => '1',
		169217 => '1',
		169338 => '1',
		169339 => '1',
		169340 => '1',
		169341 => '1',
		169342 => '1',
		169463 => '1',
		169464 => '1',
		169465 => '1',
		169466 => '1',
		169467 => '1',
		170112 => '1',
		170113 => '1',
		170114 => '1',
		170115 => '1',
		170116 => '1',
		170237 => '1',
		170238 => '1',
		170239 => '1',
		170240 => '1',
		170241 => '1',
		170362 => '1',
		170363 => '1',
		170364 => '1',
		170365 => '1',
		170366 => '1',
		170487 => '1',
		170488 => '1',
		170489 => '1',
		170490 => '1',
		170491 => '1',
		171136 => '1',
		171137 => '1',
		171138 => '1',
		171139 => '1',
		171140 => '1',
		171261 => '1',
		171262 => '1',
		171263 => '1',
		171264 => '1',
		171265 => '1',
		171386 => '1',
		171387 => '1',
		171388 => '1',
		171389 => '1',
		171390 => '1',
		171511 => '1',
		171512 => '1',
		171513 => '1',
		171514 => '1',
		171515 => '1',
		172160 => '1',
		172161 => '1',
		172162 => '1',
		172163 => '1',
		172164 => '1',
		172285 => '1',
		172286 => '1',
		172287 => '1',
		172288 => '1',
		172289 => '1',
		172410 => '1',
		172411 => '1',
		172412 => '1',
		172413 => '1',
		172414 => '1',
		172535 => '1',
		172536 => '1',
		172537 => '1',
		172538 => '1',
		172539 => '1',
		173184 => '1',
		173185 => '1',
		173186 => '1',
		173187 => '1',
		173188 => '1',
		173309 => '1',
		173310 => '1',
		173311 => '1',
		173312 => '1',
		173313 => '1',
		173434 => '1',
		173435 => '1',
		173436 => '1',
		173437 => '1',
		173438 => '1',
		173559 => '1',
		173560 => '1',
		173561 => '1',
		173562 => '1',
		173563 => '1',
		174208 => '1',
		174209 => '1',
		174210 => '1',
		174211 => '1',
		174212 => '1',
		174333 => '1',
		174334 => '1',
		174335 => '1',
		174336 => '1',
		174337 => '1',
		174458 => '1',
		174459 => '1',
		174460 => '1',
		174461 => '1',
		174462 => '1',
		174583 => '1',
		174584 => '1',
		174585 => '1',
		174586 => '1',
		174587 => '1',
		175232 => '1',
		175233 => '1',
		175234 => '1',
		175235 => '1',
		175236 => '1',
		175357 => '1',
		175358 => '1',
		175359 => '1',
		175360 => '1',
		175361 => '1',
		175482 => '1',
		175483 => '1',
		175484 => '1',
		175485 => '1',
		175486 => '1',
		175607 => '1',
		175608 => '1',
		175609 => '1',
		175610 => '1',
		175611 => '1',
		176256 => '1',
		176257 => '1',
		176258 => '1',
		176259 => '1',
		176260 => '1',
		176381 => '1',
		176382 => '1',
		176383 => '1',
		176384 => '1',
		176385 => '1',
		176506 => '1',
		176507 => '1',
		176508 => '1',
		176509 => '1',
		176510 => '1',
		176631 => '1',
		176632 => '1',
		176633 => '1',
		176634 => '1',
		176635 => '1',
		177280 => '1',
		177281 => '1',
		177282 => '1',
		177283 => '1',
		177284 => '1',
		177285 => '1',
		177286 => '1',
		177287 => '1',
		177288 => '1',
		177289 => '1',
		177290 => '1',
		177291 => '1',
		177292 => '1',
		177293 => '1',
		177294 => '1',
		177295 => '1',
		177296 => '1',
		177297 => '1',
		177298 => '1',
		177299 => '1',
		177300 => '1',
		177301 => '1',
		177302 => '1',
		177303 => '1',
		177304 => '1',
		177305 => '1',
		177306 => '1',
		177307 => '1',
		177308 => '1',
		177309 => '1',
		177310 => '1',
		177311 => '1',
		177312 => '1',
		177313 => '1',
		177314 => '1',
		177315 => '1',
		177316 => '1',
		177317 => '1',
		177318 => '1',
		177319 => '1',
		177320 => '1',
		177321 => '1',
		177322 => '1',
		177323 => '1',
		177324 => '1',
		177325 => '1',
		177326 => '1',
		177327 => '1',
		177328 => '1',
		177329 => '1',
		177330 => '1',
		177331 => '1',
		177332 => '1',
		177333 => '1',
		177334 => '1',
		177335 => '1',
		177336 => '1',
		177337 => '1',
		177338 => '1',
		177339 => '1',
		177340 => '1',
		177341 => '1',
		177342 => '1',
		177343 => '1',
		177344 => '1',
		177345 => '1',
		177346 => '1',
		177347 => '1',
		177348 => '1',
		177349 => '1',
		177350 => '1',
		177351 => '1',
		177352 => '1',
		177353 => '1',
		177354 => '1',
		177355 => '1',
		177356 => '1',
		177357 => '1',
		177358 => '1',
		177359 => '1',
		177360 => '1',
		177361 => '1',
		177362 => '1',
		177363 => '1',
		177364 => '1',
		177365 => '1',
		177366 => '1',
		177367 => '1',
		177368 => '1',
		177369 => '1',
		177370 => '1',
		177371 => '1',
		177372 => '1',
		177373 => '1',
		177374 => '1',
		177375 => '1',
		177376 => '1',
		177377 => '1',
		177378 => '1',
		177379 => '1',
		177380 => '1',
		177381 => '1',
		177382 => '1',
		177383 => '1',
		177384 => '1',
		177385 => '1',
		177386 => '1',
		177387 => '1',
		177388 => '1',
		177389 => '1',
		177390 => '1',
		177391 => '1',
		177392 => '1',
		177393 => '1',
		177394 => '1',
		177395 => '1',
		177396 => '1',
		177397 => '1',
		177398 => '1',
		177399 => '1',
		177400 => '1',
		177401 => '1',
		177402 => '1',
		177403 => '1',
		177404 => '1',
		177405 => '1',
		177406 => '1',
		177407 => '1',
		177408 => '1',
		177409 => '1',
		177410 => '1',
		177411 => '1',
		177412 => '1',
		177413 => '1',
		177414 => '1',
		177415 => '1',
		177416 => '1',
		177417 => '1',
		177418 => '1',
		177419 => '1',
		177420 => '1',
		177421 => '1',
		177422 => '1',
		177423 => '1',
		177424 => '1',
		177425 => '1',
		177426 => '1',
		177427 => '1',
		177428 => '1',
		177429 => '1',
		177430 => '1',
		177431 => '1',
		177432 => '1',
		177433 => '1',
		177434 => '1',
		177435 => '1',
		177436 => '1',
		177437 => '1',
		177438 => '1',
		177439 => '1',
		177440 => '1',
		177441 => '1',
		177442 => '1',
		177443 => '1',
		177444 => '1',
		177445 => '1',
		177446 => '1',
		177447 => '1',
		177448 => '1',
		177449 => '1',
		177450 => '1',
		177451 => '1',
		177452 => '1',
		177453 => '1',
		177454 => '1',
		177455 => '1',
		177456 => '1',
		177457 => '1',
		177458 => '1',
		177459 => '1',
		177460 => '1',
		177461 => '1',
		177462 => '1',
		177463 => '1',
		177464 => '1',
		177465 => '1',
		177466 => '1',
		177467 => '1',
		177468 => '1',
		177469 => '1',
		177470 => '1',
		177471 => '1',
		177472 => '1',
		177473 => '1',
		177474 => '1',
		177475 => '1',
		177476 => '1',
		177477 => '1',
		177478 => '1',
		177479 => '1',
		177480 => '1',
		177481 => '1',
		177482 => '1',
		177483 => '1',
		177484 => '1',
		177485 => '1',
		177486 => '1',
		177487 => '1',
		177488 => '1',
		177489 => '1',
		177490 => '1',
		177491 => '1',
		177492 => '1',
		177493 => '1',
		177494 => '1',
		177495 => '1',
		177496 => '1',
		177497 => '1',
		177498 => '1',
		177499 => '1',
		177500 => '1',
		177501 => '1',
		177502 => '1',
		177503 => '1',
		177504 => '1',
		177505 => '1',
		177506 => '1',
		177507 => '1',
		177508 => '1',
		177509 => '1',
		177510 => '1',
		177511 => '1',
		177512 => '1',
		177513 => '1',
		177514 => '1',
		177515 => '1',
		177516 => '1',
		177517 => '1',
		177518 => '1',
		177519 => '1',
		177520 => '1',
		177521 => '1',
		177522 => '1',
		177523 => '1',
		177524 => '1',
		177525 => '1',
		177526 => '1',
		177527 => '1',
		177528 => '1',
		177529 => '1',
		177530 => '1',
		177531 => '1',
		177532 => '1',
		177533 => '1',
		177534 => '1',
		177535 => '1',
		177536 => '1',
		177537 => '1',
		177538 => '1',
		177539 => '1',
		177540 => '1',
		177541 => '1',
		177542 => '1',
		177543 => '1',
		177544 => '1',
		177545 => '1',
		177546 => '1',
		177547 => '1',
		177548 => '1',
		177549 => '1',
		177550 => '1',
		177551 => '1',
		177552 => '1',
		177553 => '1',
		177554 => '1',
		177555 => '1',
		177556 => '1',
		177557 => '1',
		177558 => '1',
		177559 => '1',
		177560 => '1',
		177561 => '1',
		177562 => '1',
		177563 => '1',
		177564 => '1',
		177565 => '1',
		177566 => '1',
		177567 => '1',
		177568 => '1',
		177569 => '1',
		177570 => '1',
		177571 => '1',
		177572 => '1',
		177573 => '1',
		177574 => '1',
		177575 => '1',
		177576 => '1',
		177577 => '1',
		177578 => '1',
		177579 => '1',
		177580 => '1',
		177581 => '1',
		177582 => '1',
		177583 => '1',
		177584 => '1',
		177585 => '1',
		177586 => '1',
		177587 => '1',
		177588 => '1',
		177589 => '1',
		177590 => '1',
		177591 => '1',
		177592 => '1',
		177593 => '1',
		177594 => '1',
		177595 => '1',
		177596 => '1',
		177597 => '1',
		177598 => '1',
		177599 => '1',
		177600 => '1',
		177601 => '1',
		177602 => '1',
		177603 => '1',
		177604 => '1',
		177605 => '1',
		177606 => '1',
		177607 => '1',
		177608 => '1',
		177609 => '1',
		177610 => '1',
		177611 => '1',
		177612 => '1',
		177613 => '1',
		177614 => '1',
		177615 => '1',
		177616 => '1',
		177617 => '1',
		177618 => '1',
		177619 => '1',
		177620 => '1',
		177621 => '1',
		177622 => '1',
		177623 => '1',
		177624 => '1',
		177625 => '1',
		177626 => '1',
		177627 => '1',
		177628 => '1',
		177629 => '1',
		177630 => '1',
		177631 => '1',
		177632 => '1',
		177633 => '1',
		177634 => '1',
		177635 => '1',
		177636 => '1',
		177637 => '1',
		177638 => '1',
		177639 => '1',
		177640 => '1',
		177641 => '1',
		177642 => '1',
		177643 => '1',
		177644 => '1',
		177645 => '1',
		177646 => '1',
		177647 => '1',
		177648 => '1',
		177649 => '1',
		177650 => '1',
		177651 => '1',
		177652 => '1',
		177653 => '1',
		177654 => '1',
		177655 => '1',
		177656 => '1',
		177657 => '1',
		177658 => '1',
		177659 => '1',
		178304 => '1',
		178305 => '1',
		178306 => '1',
		178307 => '1',
		178308 => '1',
		178309 => '1',
		178310 => '1',
		178311 => '1',
		178312 => '1',
		178313 => '1',
		178314 => '1',
		178315 => '1',
		178316 => '1',
		178317 => '1',
		178318 => '1',
		178319 => '1',
		178320 => '1',
		178321 => '1',
		178322 => '1',
		178323 => '1',
		178324 => '1',
		178325 => '1',
		178326 => '1',
		178327 => '1',
		178328 => '1',
		178329 => '1',
		178330 => '1',
		178331 => '1',
		178332 => '1',
		178333 => '1',
		178334 => '1',
		178335 => '1',
		178336 => '1',
		178337 => '1',
		178338 => '1',
		178339 => '1',
		178340 => '1',
		178341 => '1',
		178342 => '1',
		178343 => '1',
		178344 => '1',
		178345 => '1',
		178346 => '1',
		178347 => '1',
		178348 => '1',
		178349 => '1',
		178350 => '1',
		178351 => '1',
		178352 => '1',
		178353 => '1',
		178354 => '1',
		178355 => '1',
		178356 => '1',
		178357 => '1',
		178358 => '1',
		178359 => '1',
		178360 => '1',
		178361 => '1',
		178362 => '1',
		178363 => '1',
		178364 => '1',
		178365 => '1',
		178366 => '1',
		178367 => '1',
		178368 => '1',
		178369 => '1',
		178370 => '1',
		178371 => '1',
		178372 => '1',
		178373 => '1',
		178374 => '1',
		178375 => '1',
		178376 => '1',
		178377 => '1',
		178378 => '1',
		178379 => '1',
		178380 => '1',
		178381 => '1',
		178382 => '1',
		178383 => '1',
		178384 => '1',
		178385 => '1',
		178386 => '1',
		178387 => '1',
		178388 => '1',
		178389 => '1',
		178390 => '1',
		178391 => '1',
		178392 => '1',
		178393 => '1',
		178394 => '1',
		178395 => '1',
		178396 => '1',
		178397 => '1',
		178398 => '1',
		178399 => '1',
		178400 => '1',
		178401 => '1',
		178402 => '1',
		178403 => '1',
		178404 => '1',
		178405 => '1',
		178406 => '1',
		178407 => '1',
		178408 => '1',
		178409 => '1',
		178410 => '1',
		178411 => '1',
		178412 => '1',
		178413 => '1',
		178414 => '1',
		178415 => '1',
		178416 => '1',
		178417 => '1',
		178418 => '1',
		178419 => '1',
		178420 => '1',
		178421 => '1',
		178422 => '1',
		178423 => '1',
		178424 => '1',
		178425 => '1',
		178426 => '1',
		178427 => '1',
		178428 => '1',
		178429 => '1',
		178430 => '1',
		178431 => '1',
		178432 => '1',
		178433 => '1',
		178434 => '1',
		178435 => '1',
		178436 => '1',
		178437 => '1',
		178438 => '1',
		178439 => '1',
		178440 => '1',
		178441 => '1',
		178442 => '1',
		178443 => '1',
		178444 => '1',
		178445 => '1',
		178446 => '1',
		178447 => '1',
		178448 => '1',
		178449 => '1',
		178450 => '1',
		178451 => '1',
		178452 => '1',
		178453 => '1',
		178454 => '1',
		178455 => '1',
		178456 => '1',
		178457 => '1',
		178458 => '1',
		178459 => '1',
		178460 => '1',
		178461 => '1',
		178462 => '1',
		178463 => '1',
		178464 => '1',
		178465 => '1',
		178466 => '1',
		178467 => '1',
		178468 => '1',
		178469 => '1',
		178470 => '1',
		178471 => '1',
		178472 => '1',
		178473 => '1',
		178474 => '1',
		178475 => '1',
		178476 => '1',
		178477 => '1',
		178478 => '1',
		178479 => '1',
		178480 => '1',
		178481 => '1',
		178482 => '1',
		178483 => '1',
		178484 => '1',
		178485 => '1',
		178486 => '1',
		178487 => '1',
		178488 => '1',
		178489 => '1',
		178490 => '1',
		178491 => '1',
		178492 => '1',
		178493 => '1',
		178494 => '1',
		178495 => '1',
		178496 => '1',
		178497 => '1',
		178498 => '1',
		178499 => '1',
		178500 => '1',
		178501 => '1',
		178502 => '1',
		178503 => '1',
		178504 => '1',
		178505 => '1',
		178506 => '1',
		178507 => '1',
		178508 => '1',
		178509 => '1',
		178510 => '1',
		178511 => '1',
		178512 => '1',
		178513 => '1',
		178514 => '1',
		178515 => '1',
		178516 => '1',
		178517 => '1',
		178518 => '1',
		178519 => '1',
		178520 => '1',
		178521 => '1',
		178522 => '1',
		178523 => '1',
		178524 => '1',
		178525 => '1',
		178526 => '1',
		178527 => '1',
		178528 => '1',
		178529 => '1',
		178530 => '1',
		178531 => '1',
		178532 => '1',
		178533 => '1',
		178534 => '1',
		178535 => '1',
		178536 => '1',
		178537 => '1',
		178538 => '1',
		178539 => '1',
		178540 => '1',
		178541 => '1',
		178542 => '1',
		178543 => '1',
		178544 => '1',
		178545 => '1',
		178546 => '1',
		178547 => '1',
		178548 => '1',
		178549 => '1',
		178550 => '1',
		178551 => '1',
		178552 => '1',
		178553 => '1',
		178554 => '1',
		178555 => '1',
		178556 => '1',
		178557 => '1',
		178558 => '1',
		178559 => '1',
		178560 => '1',
		178561 => '1',
		178562 => '1',
		178563 => '1',
		178564 => '1',
		178565 => '1',
		178566 => '1',
		178567 => '1',
		178568 => '1',
		178569 => '1',
		178570 => '1',
		178571 => '1',
		178572 => '1',
		178573 => '1',
		178574 => '1',
		178575 => '1',
		178576 => '1',
		178577 => '1',
		178578 => '1',
		178579 => '1',
		178580 => '1',
		178581 => '1',
		178582 => '1',
		178583 => '1',
		178584 => '1',
		178585 => '1',
		178586 => '1',
		178587 => '1',
		178588 => '1',
		178589 => '1',
		178590 => '1',
		178591 => '1',
		178592 => '1',
		178593 => '1',
		178594 => '1',
		178595 => '1',
		178596 => '1',
		178597 => '1',
		178598 => '1',
		178599 => '1',
		178600 => '1',
		178601 => '1',
		178602 => '1',
		178603 => '1',
		178604 => '1',
		178605 => '1',
		178606 => '1',
		178607 => '1',
		178608 => '1',
		178609 => '1',
		178610 => '1',
		178611 => '1',
		178612 => '1',
		178613 => '1',
		178614 => '1',
		178615 => '1',
		178616 => '1',
		178617 => '1',
		178618 => '1',
		178619 => '1',
		178620 => '1',
		178621 => '1',
		178622 => '1',
		178623 => '1',
		178624 => '1',
		178625 => '1',
		178626 => '1',
		178627 => '1',
		178628 => '1',
		178629 => '1',
		178630 => '1',
		178631 => '1',
		178632 => '1',
		178633 => '1',
		178634 => '1',
		178635 => '1',
		178636 => '1',
		178637 => '1',
		178638 => '1',
		178639 => '1',
		178640 => '1',
		178641 => '1',
		178642 => '1',
		178643 => '1',
		178644 => '1',
		178645 => '1',
		178646 => '1',
		178647 => '1',
		178648 => '1',
		178649 => '1',
		178650 => '1',
		178651 => '1',
		178652 => '1',
		178653 => '1',
		178654 => '1',
		178655 => '1',
		178656 => '1',
		178657 => '1',
		178658 => '1',
		178659 => '1',
		178660 => '1',
		178661 => '1',
		178662 => '1',
		178663 => '1',
		178664 => '1',
		178665 => '1',
		178666 => '1',
		178667 => '1',
		178668 => '1',
		178669 => '1',
		178670 => '1',
		178671 => '1',
		178672 => '1',
		178673 => '1',
		178674 => '1',
		178675 => '1',
		178676 => '1',
		178677 => '1',
		178678 => '1',
		178679 => '1',
		178680 => '1',
		178681 => '1',
		178682 => '1',
		178683 => '1',
		179328 => '1',
		179329 => '1',
		179330 => '1',
		179331 => '1',
		179332 => '1',
		179333 => '1',
		179334 => '1',
		179335 => '1',
		179336 => '1',
		179337 => '1',
		179338 => '1',
		179339 => '1',
		179340 => '1',
		179341 => '1',
		179342 => '1',
		179343 => '1',
		179344 => '1',
		179345 => '1',
		179346 => '1',
		179347 => '1',
		179348 => '1',
		179349 => '1',
		179350 => '1',
		179351 => '1',
		179352 => '1',
		179353 => '1',
		179354 => '1',
		179355 => '1',
		179356 => '1',
		179357 => '1',
		179358 => '1',
		179359 => '1',
		179360 => '1',
		179361 => '1',
		179362 => '1',
		179363 => '1',
		179364 => '1',
		179365 => '1',
		179366 => '1',
		179367 => '1',
		179368 => '1',
		179369 => '1',
		179370 => '1',
		179371 => '1',
		179372 => '1',
		179373 => '1',
		179374 => '1',
		179375 => '1',
		179376 => '1',
		179377 => '1',
		179378 => '1',
		179379 => '1',
		179380 => '1',
		179381 => '1',
		179382 => '1',
		179383 => '1',
		179384 => '1',
		179385 => '1',
		179386 => '1',
		179387 => '1',
		179388 => '1',
		179389 => '1',
		179390 => '1',
		179391 => '1',
		179392 => '1',
		179393 => '1',
		179394 => '1',
		179395 => '1',
		179396 => '1',
		179397 => '1',
		179398 => '1',
		179399 => '1',
		179400 => '1',
		179401 => '1',
		179402 => '1',
		179403 => '1',
		179404 => '1',
		179405 => '1',
		179406 => '1',
		179407 => '1',
		179408 => '1',
		179409 => '1',
		179410 => '1',
		179411 => '1',
		179412 => '1',
		179413 => '1',
		179414 => '1',
		179415 => '1',
		179416 => '1',
		179417 => '1',
		179418 => '1',
		179419 => '1',
		179420 => '1',
		179421 => '1',
		179422 => '1',
		179423 => '1',
		179424 => '1',
		179425 => '1',
		179426 => '1',
		179427 => '1',
		179428 => '1',
		179429 => '1',
		179430 => '1',
		179431 => '1',
		179432 => '1',
		179433 => '1',
		179434 => '1',
		179435 => '1',
		179436 => '1',
		179437 => '1',
		179438 => '1',
		179439 => '1',
		179440 => '1',
		179441 => '1',
		179442 => '1',
		179443 => '1',
		179444 => '1',
		179445 => '1',
		179446 => '1',
		179447 => '1',
		179448 => '1',
		179449 => '1',
		179450 => '1',
		179451 => '1',
		179452 => '1',
		179453 => '1',
		179454 => '1',
		179455 => '1',
		179456 => '1',
		179457 => '1',
		179458 => '1',
		179459 => '1',
		179460 => '1',
		179461 => '1',
		179462 => '1',
		179463 => '1',
		179464 => '1',
		179465 => '1',
		179466 => '1',
		179467 => '1',
		179468 => '1',
		179469 => '1',
		179470 => '1',
		179471 => '1',
		179472 => '1',
		179473 => '1',
		179474 => '1',
		179475 => '1',
		179476 => '1',
		179477 => '1',
		179478 => '1',
		179479 => '1',
		179480 => '1',
		179481 => '1',
		179482 => '1',
		179483 => '1',
		179484 => '1',
		179485 => '1',
		179486 => '1',
		179487 => '1',
		179488 => '1',
		179489 => '1',
		179490 => '1',
		179491 => '1',
		179492 => '1',
		179493 => '1',
		179494 => '1',
		179495 => '1',
		179496 => '1',
		179497 => '1',
		179498 => '1',
		179499 => '1',
		179500 => '1',
		179501 => '1',
		179502 => '1',
		179503 => '1',
		179504 => '1',
		179505 => '1',
		179506 => '1',
		179507 => '1',
		179508 => '1',
		179509 => '1',
		179510 => '1',
		179511 => '1',
		179512 => '1',
		179513 => '1',
		179514 => '1',
		179515 => '1',
		179516 => '1',
		179517 => '1',
		179518 => '1',
		179519 => '1',
		179520 => '1',
		179521 => '1',
		179522 => '1',
		179523 => '1',
		179524 => '1',
		179525 => '1',
		179526 => '1',
		179527 => '1',
		179528 => '1',
		179529 => '1',
		179530 => '1',
		179531 => '1',
		179532 => '1',
		179533 => '1',
		179534 => '1',
		179535 => '1',
		179536 => '1',
		179537 => '1',
		179538 => '1',
		179539 => '1',
		179540 => '1',
		179541 => '1',
		179542 => '1',
		179543 => '1',
		179544 => '1',
		179545 => '1',
		179546 => '1',
		179547 => '1',
		179548 => '1',
		179549 => '1',
		179550 => '1',
		179551 => '1',
		179552 => '1',
		179553 => '1',
		179554 => '1',
		179555 => '1',
		179556 => '1',
		179557 => '1',
		179558 => '1',
		179559 => '1',
		179560 => '1',
		179561 => '1',
		179562 => '1',
		179563 => '1',
		179564 => '1',
		179565 => '1',
		179566 => '1',
		179567 => '1',
		179568 => '1',
		179569 => '1',
		179570 => '1',
		179571 => '1',
		179572 => '1',
		179573 => '1',
		179574 => '1',
		179575 => '1',
		179576 => '1',
		179577 => '1',
		179578 => '1',
		179579 => '1',
		179580 => '1',
		179581 => '1',
		179582 => '1',
		179583 => '1',
		179584 => '1',
		179585 => '1',
		179586 => '1',
		179587 => '1',
		179588 => '1',
		179589 => '1',
		179590 => '1',
		179591 => '1',
		179592 => '1',
		179593 => '1',
		179594 => '1',
		179595 => '1',
		179596 => '1',
		179597 => '1',
		179598 => '1',
		179599 => '1',
		179600 => '1',
		179601 => '1',
		179602 => '1',
		179603 => '1',
		179604 => '1',
		179605 => '1',
		179606 => '1',
		179607 => '1',
		179608 => '1',
		179609 => '1',
		179610 => '1',
		179611 => '1',
		179612 => '1',
		179613 => '1',
		179614 => '1',
		179615 => '1',
		179616 => '1',
		179617 => '1',
		179618 => '1',
		179619 => '1',
		179620 => '1',
		179621 => '1',
		179622 => '1',
		179623 => '1',
		179624 => '1',
		179625 => '1',
		179626 => '1',
		179627 => '1',
		179628 => '1',
		179629 => '1',
		179630 => '1',
		179631 => '1',
		179632 => '1',
		179633 => '1',
		179634 => '1',
		179635 => '1',
		179636 => '1',
		179637 => '1',
		179638 => '1',
		179639 => '1',
		179640 => '1',
		179641 => '1',
		179642 => '1',
		179643 => '1',
		179644 => '1',
		179645 => '1',
		179646 => '1',
		179647 => '1',
		179648 => '1',
		179649 => '1',
		179650 => '1',
		179651 => '1',
		179652 => '1',
		179653 => '1',
		179654 => '1',
		179655 => '1',
		179656 => '1',
		179657 => '1',
		179658 => '1',
		179659 => '1',
		179660 => '1',
		179661 => '1',
		179662 => '1',
		179663 => '1',
		179664 => '1',
		179665 => '1',
		179666 => '1',
		179667 => '1',
		179668 => '1',
		179669 => '1',
		179670 => '1',
		179671 => '1',
		179672 => '1',
		179673 => '1',
		179674 => '1',
		179675 => '1',
		179676 => '1',
		179677 => '1',
		179678 => '1',
		179679 => '1',
		179680 => '1',
		179681 => '1',
		179682 => '1',
		179683 => '1',
		179684 => '1',
		179685 => '1',
		179686 => '1',
		179687 => '1',
		179688 => '1',
		179689 => '1',
		179690 => '1',
		179691 => '1',
		179692 => '1',
		179693 => '1',
		179694 => '1',
		179695 => '1',
		179696 => '1',
		179697 => '1',
		179698 => '1',
		179699 => '1',
		179700 => '1',
		179701 => '1',
		179702 => '1',
		179703 => '1',
		179704 => '1',
		179705 => '1',
		179706 => '1',
		179707 => '1',
		180352 => '1',
		180353 => '1',
		180354 => '1',
		180355 => '1',
		180356 => '1',
		180357 => '1',
		180358 => '1',
		180359 => '1',
		180360 => '1',
		180361 => '1',
		180362 => '1',
		180363 => '1',
		180364 => '1',
		180365 => '1',
		180366 => '1',
		180367 => '1',
		180368 => '1',
		180369 => '1',
		180370 => '1',
		180371 => '1',
		180372 => '1',
		180373 => '1',
		180374 => '1',
		180375 => '1',
		180376 => '1',
		180377 => '1',
		180378 => '1',
		180379 => '1',
		180380 => '1',
		180381 => '1',
		180382 => '1',
		180383 => '1',
		180384 => '1',
		180385 => '1',
		180386 => '1',
		180387 => '1',
		180388 => '1',
		180389 => '1',
		180390 => '1',
		180391 => '1',
		180392 => '1',
		180393 => '1',
		180394 => '1',
		180395 => '1',
		180396 => '1',
		180397 => '1',
		180398 => '1',
		180399 => '1',
		180400 => '1',
		180401 => '1',
		180402 => '1',
		180403 => '1',
		180404 => '1',
		180405 => '1',
		180406 => '1',
		180407 => '1',
		180408 => '1',
		180409 => '1',
		180410 => '1',
		180411 => '1',
		180412 => '1',
		180413 => '1',
		180414 => '1',
		180415 => '1',
		180416 => '1',
		180417 => '1',
		180418 => '1',
		180419 => '1',
		180420 => '1',
		180421 => '1',
		180422 => '1',
		180423 => '1',
		180424 => '1',
		180425 => '1',
		180426 => '1',
		180427 => '1',
		180428 => '1',
		180429 => '1',
		180430 => '1',
		180431 => '1',
		180432 => '1',
		180433 => '1',
		180434 => '1',
		180435 => '1',
		180436 => '1',
		180437 => '1',
		180438 => '1',
		180439 => '1',
		180440 => '1',
		180441 => '1',
		180442 => '1',
		180443 => '1',
		180444 => '1',
		180445 => '1',
		180446 => '1',
		180447 => '1',
		180448 => '1',
		180449 => '1',
		180450 => '1',
		180451 => '1',
		180452 => '1',
		180453 => '1',
		180454 => '1',
		180455 => '1',
		180456 => '1',
		180457 => '1',
		180458 => '1',
		180459 => '1',
		180460 => '1',
		180461 => '1',
		180462 => '1',
		180463 => '1',
		180464 => '1',
		180465 => '1',
		180466 => '1',
		180467 => '1',
		180468 => '1',
		180469 => '1',
		180470 => '1',
		180471 => '1',
		180472 => '1',
		180473 => '1',
		180474 => '1',
		180475 => '1',
		180476 => '1',
		180477 => '1',
		180478 => '1',
		180479 => '1',
		180480 => '1',
		180481 => '1',
		180482 => '1',
		180483 => '1',
		180484 => '1',
		180485 => '1',
		180486 => '1',
		180487 => '1',
		180488 => '1',
		180489 => '1',
		180490 => '1',
		180491 => '1',
		180492 => '1',
		180493 => '1',
		180494 => '1',
		180495 => '1',
		180496 => '1',
		180497 => '1',
		180498 => '1',
		180499 => '1',
		180500 => '1',
		180501 => '1',
		180502 => '1',
		180503 => '1',
		180504 => '1',
		180505 => '1',
		180506 => '1',
		180507 => '1',
		180508 => '1',
		180509 => '1',
		180510 => '1',
		180511 => '1',
		180512 => '1',
		180513 => '1',
		180514 => '1',
		180515 => '1',
		180516 => '1',
		180517 => '1',
		180518 => '1',
		180519 => '1',
		180520 => '1',
		180521 => '1',
		180522 => '1',
		180523 => '1',
		180524 => '1',
		180525 => '1',
		180526 => '1',
		180527 => '1',
		180528 => '1',
		180529 => '1',
		180530 => '1',
		180531 => '1',
		180532 => '1',
		180533 => '1',
		180534 => '1',
		180535 => '1',
		180536 => '1',
		180537 => '1',
		180538 => '1',
		180539 => '1',
		180540 => '1',
		180541 => '1',
		180542 => '1',
		180543 => '1',
		180544 => '1',
		180545 => '1',
		180546 => '1',
		180547 => '1',
		180548 => '1',
		180549 => '1',
		180550 => '1',
		180551 => '1',
		180552 => '1',
		180553 => '1',
		180554 => '1',
		180555 => '1',
		180556 => '1',
		180557 => '1',
		180558 => '1',
		180559 => '1',
		180560 => '1',
		180561 => '1',
		180562 => '1',
		180563 => '1',
		180564 => '1',
		180565 => '1',
		180566 => '1',
		180567 => '1',
		180568 => '1',
		180569 => '1',
		180570 => '1',
		180571 => '1',
		180572 => '1',
		180573 => '1',
		180574 => '1',
		180575 => '1',
		180576 => '1',
		180577 => '1',
		180578 => '1',
		180579 => '1',
		180580 => '1',
		180581 => '1',
		180582 => '1',
		180583 => '1',
		180584 => '1',
		180585 => '1',
		180586 => '1',
		180587 => '1',
		180588 => '1',
		180589 => '1',
		180590 => '1',
		180591 => '1',
		180592 => '1',
		180593 => '1',
		180594 => '1',
		180595 => '1',
		180596 => '1',
		180597 => '1',
		180598 => '1',
		180599 => '1',
		180600 => '1',
		180601 => '1',
		180602 => '1',
		180603 => '1',
		180604 => '1',
		180605 => '1',
		180606 => '1',
		180607 => '1',
		180608 => '1',
		180609 => '1',
		180610 => '1',
		180611 => '1',
		180612 => '1',
		180613 => '1',
		180614 => '1',
		180615 => '1',
		180616 => '1',
		180617 => '1',
		180618 => '1',
		180619 => '1',
		180620 => '1',
		180621 => '1',
		180622 => '1',
		180623 => '1',
		180624 => '1',
		180625 => '1',
		180626 => '1',
		180627 => '1',
		180628 => '1',
		180629 => '1',
		180630 => '1',
		180631 => '1',
		180632 => '1',
		180633 => '1',
		180634 => '1',
		180635 => '1',
		180636 => '1',
		180637 => '1',
		180638 => '1',
		180639 => '1',
		180640 => '1',
		180641 => '1',
		180642 => '1',
		180643 => '1',
		180644 => '1',
		180645 => '1',
		180646 => '1',
		180647 => '1',
		180648 => '1',
		180649 => '1',
		180650 => '1',
		180651 => '1',
		180652 => '1',
		180653 => '1',
		180654 => '1',
		180655 => '1',
		180656 => '1',
		180657 => '1',
		180658 => '1',
		180659 => '1',
		180660 => '1',
		180661 => '1',
		180662 => '1',
		180663 => '1',
		180664 => '1',
		180665 => '1',
		180666 => '1',
		180667 => '1',
		180668 => '1',
		180669 => '1',
		180670 => '1',
		180671 => '1',
		180672 => '1',
		180673 => '1',
		180674 => '1',
		180675 => '1',
		180676 => '1',
		180677 => '1',
		180678 => '1',
		180679 => '1',
		180680 => '1',
		180681 => '1',
		180682 => '1',
		180683 => '1',
		180684 => '1',
		180685 => '1',
		180686 => '1',
		180687 => '1',
		180688 => '1',
		180689 => '1',
		180690 => '1',
		180691 => '1',
		180692 => '1',
		180693 => '1',
		180694 => '1',
		180695 => '1',
		180696 => '1',
		180697 => '1',
		180698 => '1',
		180699 => '1',
		180700 => '1',
		180701 => '1',
		180702 => '1',
		180703 => '1',
		180704 => '1',
		180705 => '1',
		180706 => '1',
		180707 => '1',
		180708 => '1',
		180709 => '1',
		180710 => '1',
		180711 => '1',
		180712 => '1',
		180713 => '1',
		180714 => '1',
		180715 => '1',
		180716 => '1',
		180717 => '1',
		180718 => '1',
		180719 => '1',
		180720 => '1',
		180721 => '1',
		180722 => '1',
		180723 => '1',
		180724 => '1',
		180725 => '1',
		180726 => '1',
		180727 => '1',
		180728 => '1',
		180729 => '1',
		180730 => '1',
		180731 => '1',
		181376 => '1',
		181377 => '1',
		181378 => '1',
		181379 => '1',
		181380 => '1',
		181381 => '1',
		181382 => '1',
		181383 => '1',
		181384 => '1',
		181385 => '1',
		181386 => '1',
		181387 => '1',
		181388 => '1',
		181389 => '1',
		181390 => '1',
		181391 => '1',
		181392 => '1',
		181393 => '1',
		181394 => '1',
		181395 => '1',
		181396 => '1',
		181397 => '1',
		181398 => '1',
		181399 => '1',
		181400 => '1',
		181401 => '1',
		181402 => '1',
		181403 => '1',
		181404 => '1',
		181405 => '1',
		181406 => '1',
		181407 => '1',
		181408 => '1',
		181409 => '1',
		181410 => '1',
		181411 => '1',
		181412 => '1',
		181413 => '1',
		181414 => '1',
		181415 => '1',
		181416 => '1',
		181417 => '1',
		181418 => '1',
		181419 => '1',
		181420 => '1',
		181421 => '1',
		181422 => '1',
		181423 => '1',
		181424 => '1',
		181425 => '1',
		181426 => '1',
		181427 => '1',
		181428 => '1',
		181429 => '1',
		181430 => '1',
		181431 => '1',
		181432 => '1',
		181433 => '1',
		181434 => '1',
		181435 => '1',
		181436 => '1',
		181437 => '1',
		181438 => '1',
		181439 => '1',
		181440 => '1',
		181441 => '1',
		181442 => '1',
		181443 => '1',
		181444 => '1',
		181445 => '1',
		181446 => '1',
		181447 => '1',
		181448 => '1',
		181449 => '1',
		181450 => '1',
		181451 => '1',
		181452 => '1',
		181453 => '1',
		181454 => '1',
		181455 => '1',
		181456 => '1',
		181457 => '1',
		181458 => '1',
		181459 => '1',
		181460 => '1',
		181461 => '1',
		181462 => '1',
		181463 => '1',
		181464 => '1',
		181465 => '1',
		181466 => '1',
		181467 => '1',
		181468 => '1',
		181469 => '1',
		181470 => '1',
		181471 => '1',
		181472 => '1',
		181473 => '1',
		181474 => '1',
		181475 => '1',
		181476 => '1',
		181477 => '1',
		181478 => '1',
		181479 => '1',
		181480 => '1',
		181481 => '1',
		181482 => '1',
		181483 => '1',
		181484 => '1',
		181485 => '1',
		181486 => '1',
		181487 => '1',
		181488 => '1',
		181489 => '1',
		181490 => '1',
		181491 => '1',
		181492 => '1',
		181493 => '1',
		181494 => '1',
		181495 => '1',
		181496 => '1',
		181497 => '1',
		181498 => '1',
		181499 => '1',
		181500 => '1',
		181501 => '1',
		181502 => '1',
		181503 => '1',
		181504 => '1',
		181505 => '1',
		181506 => '1',
		181507 => '1',
		181508 => '1',
		181509 => '1',
		181510 => '1',
		181511 => '1',
		181512 => '1',
		181513 => '1',
		181514 => '1',
		181515 => '1',
		181516 => '1',
		181517 => '1',
		181518 => '1',
		181519 => '1',
		181520 => '1',
		181521 => '1',
		181522 => '1',
		181523 => '1',
		181524 => '1',
		181525 => '1',
		181526 => '1',
		181527 => '1',
		181528 => '1',
		181529 => '1',
		181530 => '1',
		181531 => '1',
		181532 => '1',
		181533 => '1',
		181534 => '1',
		181535 => '1',
		181536 => '1',
		181537 => '1',
		181538 => '1',
		181539 => '1',
		181540 => '1',
		181541 => '1',
		181542 => '1',
		181543 => '1',
		181544 => '1',
		181545 => '1',
		181546 => '1',
		181547 => '1',
		181548 => '1',
		181549 => '1',
		181550 => '1',
		181551 => '1',
		181552 => '1',
		181553 => '1',
		181554 => '1',
		181555 => '1',
		181556 => '1',
		181557 => '1',
		181558 => '1',
		181559 => '1',
		181560 => '1',
		181561 => '1',
		181562 => '1',
		181563 => '1',
		181564 => '1',
		181565 => '1',
		181566 => '1',
		181567 => '1',
		181568 => '1',
		181569 => '1',
		181570 => '1',
		181571 => '1',
		181572 => '1',
		181573 => '1',
		181574 => '1',
		181575 => '1',
		181576 => '1',
		181577 => '1',
		181578 => '1',
		181579 => '1',
		181580 => '1',
		181581 => '1',
		181582 => '1',
		181583 => '1',
		181584 => '1',
		181585 => '1',
		181586 => '1',
		181587 => '1',
		181588 => '1',
		181589 => '1',
		181590 => '1',
		181591 => '1',
		181592 => '1',
		181593 => '1',
		181594 => '1',
		181595 => '1',
		181596 => '1',
		181597 => '1',
		181598 => '1',
		181599 => '1',
		181600 => '1',
		181601 => '1',
		181602 => '1',
		181603 => '1',
		181604 => '1',
		181605 => '1',
		181606 => '1',
		181607 => '1',
		181608 => '1',
		181609 => '1',
		181610 => '1',
		181611 => '1',
		181612 => '1',
		181613 => '1',
		181614 => '1',
		181615 => '1',
		181616 => '1',
		181617 => '1',
		181618 => '1',
		181619 => '1',
		181620 => '1',
		181621 => '1',
		181622 => '1',
		181623 => '1',
		181624 => '1',
		181625 => '1',
		181626 => '1',
		181627 => '1',
		181628 => '1',
		181629 => '1',
		181630 => '1',
		181631 => '1',
		181632 => '1',
		181633 => '1',
		181634 => '1',
		181635 => '1',
		181636 => '1',
		181637 => '1',
		181638 => '1',
		181639 => '1',
		181640 => '1',
		181641 => '1',
		181642 => '1',
		181643 => '1',
		181644 => '1',
		181645 => '1',
		181646 => '1',
		181647 => '1',
		181648 => '1',
		181649 => '1',
		181650 => '1',
		181651 => '1',
		181652 => '1',
		181653 => '1',
		181654 => '1',
		181655 => '1',
		181656 => '1',
		181657 => '1',
		181658 => '1',
		181659 => '1',
		181660 => '1',
		181661 => '1',
		181662 => '1',
		181663 => '1',
		181664 => '1',
		181665 => '1',
		181666 => '1',
		181667 => '1',
		181668 => '1',
		181669 => '1',
		181670 => '1',
		181671 => '1',
		181672 => '1',
		181673 => '1',
		181674 => '1',
		181675 => '1',
		181676 => '1',
		181677 => '1',
		181678 => '1',
		181679 => '1',
		181680 => '1',
		181681 => '1',
		181682 => '1',
		181683 => '1',
		181684 => '1',
		181685 => '1',
		181686 => '1',
		181687 => '1',
		181688 => '1',
		181689 => '1',
		181690 => '1',
		181691 => '1',
		181692 => '1',
		181693 => '1',
		181694 => '1',
		181695 => '1',
		181696 => '1',
		181697 => '1',
		181698 => '1',
		181699 => '1',
		181700 => '1',
		181701 => '1',
		181702 => '1',
		181703 => '1',
		181704 => '1',
		181705 => '1',
		181706 => '1',
		181707 => '1',
		181708 => '1',
		181709 => '1',
		181710 => '1',
		181711 => '1',
		181712 => '1',
		181713 => '1',
		181714 => '1',
		181715 => '1',
		181716 => '1',
		181717 => '1',
		181718 => '1',
		181719 => '1',
		181720 => '1',
		181721 => '1',
		181722 => '1',
		181723 => '1',
		181724 => '1',
		181725 => '1',
		181726 => '1',
		181727 => '1',
		181728 => '1',
		181729 => '1',
		181730 => '1',
		181731 => '1',
		181732 => '1',
		181733 => '1',
		181734 => '1',
		181735 => '1',
		181736 => '1',
		181737 => '1',
		181738 => '1',
		181739 => '1',
		181740 => '1',
		181741 => '1',
		181742 => '1',
		181743 => '1',
		181744 => '1',
		181745 => '1',
		181746 => '1',
		181747 => '1',
		181748 => '1',
		181749 => '1',
		181750 => '1',
		181751 => '1',
		181752 => '1',
		181753 => '1',
		181754 => '1',
		181755 => '1',
		182400 => '1',
		182401 => '1',
		182402 => '1',
		182403 => '1',
		182404 => '1',
		182525 => '1',
		182526 => '1',
		182527 => '1',
		182528 => '1',
		182529 => '1',
		182650 => '1',
		182651 => '1',
		182652 => '1',
		182653 => '1',
		182654 => '1',
		182775 => '1',
		182776 => '1',
		182777 => '1',
		182778 => '1',
		182779 => '1',
		183424 => '1',
		183425 => '1',
		183426 => '1',
		183427 => '1',
		183428 => '1',
		183549 => '1',
		183550 => '1',
		183551 => '1',
		183552 => '1',
		183553 => '1',
		183674 => '1',
		183675 => '1',
		183676 => '1',
		183677 => '1',
		183678 => '1',
		183799 => '1',
		183800 => '1',
		183801 => '1',
		183802 => '1',
		183803 => '1',
		184448 => '1',
		184449 => '1',
		184450 => '1',
		184451 => '1',
		184452 => '1',
		184573 => '1',
		184574 => '1',
		184575 => '1',
		184576 => '1',
		184577 => '1',
		184698 => '1',
		184699 => '1',
		184700 => '1',
		184701 => '1',
		184702 => '1',
		184823 => '1',
		184824 => '1',
		184825 => '1',
		184826 => '1',
		184827 => '1',
		185472 => '1',
		185473 => '1',
		185474 => '1',
		185475 => '1',
		185476 => '1',
		185597 => '1',
		185598 => '1',
		185599 => '1',
		185600 => '1',
		185601 => '1',
		185722 => '1',
		185723 => '1',
		185724 => '1',
		185725 => '1',
		185726 => '1',
		185847 => '1',
		185848 => '1',
		185849 => '1',
		185850 => '1',
		185851 => '1',
		186496 => '1',
		186497 => '1',
		186498 => '1',
		186499 => '1',
		186500 => '1',
		186621 => '1',
		186622 => '1',
		186623 => '1',
		186624 => '1',
		186625 => '1',
		186746 => '1',
		186747 => '1',
		186748 => '1',
		186749 => '1',
		186750 => '1',
		186871 => '1',
		186872 => '1',
		186873 => '1',
		186874 => '1',
		186875 => '1',
		187520 => '1',
		187521 => '1',
		187522 => '1',
		187523 => '1',
		187524 => '1',
		187645 => '1',
		187646 => '1',
		187647 => '1',
		187648 => '1',
		187649 => '1',
		187770 => '1',
		187771 => '1',
		187772 => '1',
		187773 => '1',
		187774 => '1',
		187895 => '1',
		187896 => '1',
		187897 => '1',
		187898 => '1',
		187899 => '1',
		188544 => '1',
		188545 => '1',
		188546 => '1',
		188547 => '1',
		188548 => '1',
		188669 => '1',
		188670 => '1',
		188671 => '1',
		188672 => '1',
		188673 => '1',
		188794 => '1',
		188795 => '1',
		188796 => '1',
		188797 => '1',
		188798 => '1',
		188919 => '1',
		188920 => '1',
		188921 => '1',
		188922 => '1',
		188923 => '1',
		189568 => '1',
		189569 => '1',
		189570 => '1',
		189571 => '1',
		189572 => '1',
		189693 => '1',
		189694 => '1',
		189695 => '1',
		189696 => '1',
		189697 => '1',
		189818 => '1',
		189819 => '1',
		189820 => '1',
		189821 => '1',
		189822 => '1',
		189943 => '1',
		189944 => '1',
		189945 => '1',
		189946 => '1',
		189947 => '1',
		190592 => '1',
		190593 => '1',
		190594 => '1',
		190595 => '1',
		190596 => '1',
		190717 => '1',
		190718 => '1',
		190719 => '1',
		190720 => '1',
		190721 => '1',
		190842 => '1',
		190843 => '1',
		190844 => '1',
		190845 => '1',
		190846 => '1',
		190967 => '1',
		190968 => '1',
		190969 => '1',
		190970 => '1',
		190971 => '1',
		191616 => '1',
		191617 => '1',
		191618 => '1',
		191619 => '1',
		191620 => '1',
		191741 => '1',
		191742 => '1',
		191743 => '1',
		191744 => '1',
		191745 => '1',
		191866 => '1',
		191867 => '1',
		191868 => '1',
		191869 => '1',
		191870 => '1',
		191991 => '1',
		191992 => '1',
		191993 => '1',
		191994 => '1',
		191995 => '1',
		192640 => '1',
		192641 => '1',
		192642 => '1',
		192643 => '1',
		192644 => '1',
		192765 => '1',
		192766 => '1',
		192767 => '1',
		192768 => '1',
		192769 => '1',
		192890 => '1',
		192891 => '1',
		192892 => '1',
		192893 => '1',
		192894 => '1',
		193015 => '1',
		193016 => '1',
		193017 => '1',
		193018 => '1',
		193019 => '1',
		193664 => '1',
		193665 => '1',
		193666 => '1',
		193667 => '1',
		193668 => '1',
		193789 => '1',
		193790 => '1',
		193791 => '1',
		193792 => '1',
		193793 => '1',
		193914 => '1',
		193915 => '1',
		193916 => '1',
		193917 => '1',
		193918 => '1',
		194039 => '1',
		194040 => '1',
		194041 => '1',
		194042 => '1',
		194043 => '1',
		194688 => '1',
		194689 => '1',
		194690 => '1',
		194691 => '1',
		194692 => '1',
		194813 => '1',
		194814 => '1',
		194815 => '1',
		194816 => '1',
		194817 => '1',
		194938 => '1',
		194939 => '1',
		194940 => '1',
		194941 => '1',
		194942 => '1',
		195063 => '1',
		195064 => '1',
		195065 => '1',
		195066 => '1',
		195067 => '1',
		195712 => '1',
		195713 => '1',
		195714 => '1',
		195715 => '1',
		195716 => '1',
		195837 => '1',
		195838 => '1',
		195839 => '1',
		195840 => '1',
		195841 => '1',
		195962 => '1',
		195963 => '1',
		195964 => '1',
		195965 => '1',
		195966 => '1',
		196087 => '1',
		196088 => '1',
		196089 => '1',
		196090 => '1',
		196091 => '1',
		196736 => '1',
		196737 => '1',
		196738 => '1',
		196739 => '1',
		196740 => '1',
		196861 => '1',
		196862 => '1',
		196863 => '1',
		196864 => '1',
		196865 => '1',
		196986 => '1',
		196987 => '1',
		196988 => '1',
		196989 => '1',
		196990 => '1',
		197111 => '1',
		197112 => '1',
		197113 => '1',
		197114 => '1',
		197115 => '1',
		197760 => '1',
		197761 => '1',
		197762 => '1',
		197763 => '1',
		197764 => '1',
		197885 => '1',
		197886 => '1',
		197887 => '1',
		197888 => '1',
		197889 => '1',
		198010 => '1',
		198011 => '1',
		198012 => '1',
		198013 => '1',
		198014 => '1',
		198135 => '1',
		198136 => '1',
		198137 => '1',
		198138 => '1',
		198139 => '1',
		198784 => '1',
		198785 => '1',
		198786 => '1',
		198787 => '1',
		198788 => '1',
		198909 => '1',
		198910 => '1',
		198911 => '1',
		198912 => '1',
		198913 => '1',
		199034 => '1',
		199035 => '1',
		199036 => '1',
		199037 => '1',
		199038 => '1',
		199159 => '1',
		199160 => '1',
		199161 => '1',
		199162 => '1',
		199163 => '1',
		199808 => '1',
		199809 => '1',
		199810 => '1',
		199811 => '1',
		199812 => '1',
		199933 => '1',
		199934 => '1',
		199935 => '1',
		199936 => '1',
		199937 => '1',
		200058 => '1',
		200059 => '1',
		200060 => '1',
		200061 => '1',
		200062 => '1',
		200183 => '1',
		200184 => '1',
		200185 => '1',
		200186 => '1',
		200187 => '1',
		200832 => '1',
		200833 => '1',
		200834 => '1',
		200835 => '1',
		200836 => '1',
		200957 => '1',
		200958 => '1',
		200959 => '1',
		200960 => '1',
		200961 => '1',
		201082 => '1',
		201083 => '1',
		201084 => '1',
		201085 => '1',
		201086 => '1',
		201207 => '1',
		201208 => '1',
		201209 => '1',
		201210 => '1',
		201211 => '1',
		201856 => '1',
		201857 => '1',
		201858 => '1',
		201859 => '1',
		201860 => '1',
		201981 => '1',
		201982 => '1',
		201983 => '1',
		201984 => '1',
		201985 => '1',
		202106 => '1',
		202107 => '1',
		202108 => '1',
		202109 => '1',
		202110 => '1',
		202231 => '1',
		202232 => '1',
		202233 => '1',
		202234 => '1',
		202235 => '1',
		202880 => '1',
		202881 => '1',
		202882 => '1',
		202883 => '1',
		202884 => '1',
		203005 => '1',
		203006 => '1',
		203007 => '1',
		203008 => '1',
		203009 => '1',
		203130 => '1',
		203131 => '1',
		203132 => '1',
		203133 => '1',
		203134 => '1',
		203255 => '1',
		203256 => '1',
		203257 => '1',
		203258 => '1',
		203259 => '1',
		203904 => '1',
		203905 => '1',
		203906 => '1',
		203907 => '1',
		203908 => '1',
		204029 => '1',
		204030 => '1',
		204031 => '1',
		204032 => '1',
		204033 => '1',
		204154 => '1',
		204155 => '1',
		204156 => '1',
		204157 => '1',
		204158 => '1',
		204279 => '1',
		204280 => '1',
		204281 => '1',
		204282 => '1',
		204283 => '1',
		204928 => '1',
		204929 => '1',
		204930 => '1',
		204931 => '1',
		204932 => '1',
		205053 => '1',
		205054 => '1',
		205055 => '1',
		205056 => '1',
		205057 => '1',
		205178 => '1',
		205179 => '1',
		205180 => '1',
		205181 => '1',
		205182 => '1',
		205303 => '1',
		205304 => '1',
		205305 => '1',
		205306 => '1',
		205307 => '1',
		205952 => '1',
		205953 => '1',
		205954 => '1',
		205955 => '1',
		205956 => '1',
		206077 => '1',
		206078 => '1',
		206079 => '1',
		206080 => '1',
		206081 => '1',
		206202 => '1',
		206203 => '1',
		206204 => '1',
		206205 => '1',
		206206 => '1',
		206327 => '1',
		206328 => '1',
		206329 => '1',
		206330 => '1',
		206331 => '1',
		206976 => '1',
		206977 => '1',
		206978 => '1',
		206979 => '1',
		206980 => '1',
		207101 => '1',
		207102 => '1',
		207103 => '1',
		207104 => '1',
		207105 => '1',
		207226 => '1',
		207227 => '1',
		207228 => '1',
		207229 => '1',
		207230 => '1',
		207351 => '1',
		207352 => '1',
		207353 => '1',
		207354 => '1',
		207355 => '1',
		208000 => '1',
		208001 => '1',
		208002 => '1',
		208003 => '1',
		208004 => '1',
		208125 => '1',
		208126 => '1',
		208127 => '1',
		208128 => '1',
		208129 => '1',
		208250 => '1',
		208251 => '1',
		208252 => '1',
		208253 => '1',
		208254 => '1',
		208375 => '1',
		208376 => '1',
		208377 => '1',
		208378 => '1',
		208379 => '1',
		209024 => '1',
		209025 => '1',
		209026 => '1',
		209027 => '1',
		209028 => '1',
		209149 => '1',
		209150 => '1',
		209151 => '1',
		209152 => '1',
		209153 => '1',
		209274 => '1',
		209275 => '1',
		209276 => '1',
		209277 => '1',
		209278 => '1',
		209399 => '1',
		209400 => '1',
		209401 => '1',
		209402 => '1',
		209403 => '1',
		210048 => '1',
		210049 => '1',
		210050 => '1',
		210051 => '1',
		210052 => '1',
		210173 => '1',
		210174 => '1',
		210175 => '1',
		210176 => '1',
		210177 => '1',
		210298 => '1',
		210299 => '1',
		210300 => '1',
		210301 => '1',
		210302 => '1',
		210423 => '1',
		210424 => '1',
		210425 => '1',
		210426 => '1',
		210427 => '1',
		211072 => '1',
		211073 => '1',
		211074 => '1',
		211075 => '1',
		211076 => '1',
		211197 => '1',
		211198 => '1',
		211199 => '1',
		211200 => '1',
		211201 => '1',
		211322 => '1',
		211323 => '1',
		211324 => '1',
		211325 => '1',
		211326 => '1',
		211447 => '1',
		211448 => '1',
		211449 => '1',
		211450 => '1',
		211451 => '1',
		212096 => '1',
		212097 => '1',
		212098 => '1',
		212099 => '1',
		212100 => '1',
		212221 => '1',
		212222 => '1',
		212223 => '1',
		212224 => '1',
		212225 => '1',
		212346 => '1',
		212347 => '1',
		212348 => '1',
		212349 => '1',
		212350 => '1',
		212471 => '1',
		212472 => '1',
		212473 => '1',
		212474 => '1',
		212475 => '1',
		213120 => '1',
		213121 => '1',
		213122 => '1',
		213123 => '1',
		213124 => '1',
		213245 => '1',
		213246 => '1',
		213247 => '1',
		213248 => '1',
		213249 => '1',
		213370 => '1',
		213371 => '1',
		213372 => '1',
		213373 => '1',
		213374 => '1',
		213495 => '1',
		213496 => '1',
		213497 => '1',
		213498 => '1',
		213499 => '1',
		214144 => '1',
		214145 => '1',
		214146 => '1',
		214147 => '1',
		214148 => '1',
		214269 => '1',
		214270 => '1',
		214271 => '1',
		214272 => '1',
		214273 => '1',
		214394 => '1',
		214395 => '1',
		214396 => '1',
		214397 => '1',
		214398 => '1',
		214519 => '1',
		214520 => '1',
		214521 => '1',
		214522 => '1',
		214523 => '1',
		215168 => '1',
		215169 => '1',
		215170 => '1',
		215171 => '1',
		215172 => '1',
		215293 => '1',
		215294 => '1',
		215295 => '1',
		215296 => '1',
		215297 => '1',
		215418 => '1',
		215419 => '1',
		215420 => '1',
		215421 => '1',
		215422 => '1',
		215543 => '1',
		215544 => '1',
		215545 => '1',
		215546 => '1',
		215547 => '1',
		216192 => '1',
		216193 => '1',
		216194 => '1',
		216195 => '1',
		216196 => '1',
		216317 => '1',
		216318 => '1',
		216319 => '1',
		216320 => '1',
		216321 => '1',
		216442 => '1',
		216443 => '1',
		216444 => '1',
		216445 => '1',
		216446 => '1',
		216567 => '1',
		216568 => '1',
		216569 => '1',
		216570 => '1',
		216571 => '1',
		217216 => '1',
		217217 => '1',
		217218 => '1',
		217219 => '1',
		217220 => '1',
		217341 => '1',
		217342 => '1',
		217343 => '1',
		217344 => '1',
		217345 => '1',
		217466 => '1',
		217467 => '1',
		217468 => '1',
		217469 => '1',
		217470 => '1',
		217591 => '1',
		217592 => '1',
		217593 => '1',
		217594 => '1',
		217595 => '1',
		218240 => '1',
		218241 => '1',
		218242 => '1',
		218243 => '1',
		218244 => '1',
		218365 => '1',
		218366 => '1',
		218367 => '1',
		218368 => '1',
		218369 => '1',
		218490 => '1',
		218491 => '1',
		218492 => '1',
		218493 => '1',
		218494 => '1',
		218615 => '1',
		218616 => '1',
		218617 => '1',
		218618 => '1',
		218619 => '1',
		219264 => '1',
		219265 => '1',
		219266 => '1',
		219267 => '1',
		219268 => '1',
		219389 => '1',
		219390 => '1',
		219391 => '1',
		219392 => '1',
		219393 => '1',
		219514 => '1',
		219515 => '1',
		219516 => '1',
		219517 => '1',
		219518 => '1',
		219639 => '1',
		219640 => '1',
		219641 => '1',
		219642 => '1',
		219643 => '1',
		220288 => '1',
		220289 => '1',
		220290 => '1',
		220291 => '1',
		220292 => '1',
		220413 => '1',
		220414 => '1',
		220415 => '1',
		220416 => '1',
		220417 => '1',
		220538 => '1',
		220539 => '1',
		220540 => '1',
		220541 => '1',
		220542 => '1',
		220663 => '1',
		220664 => '1',
		220665 => '1',
		220666 => '1',
		220667 => '1',
		221312 => '1',
		221313 => '1',
		221314 => '1',
		221315 => '1',
		221316 => '1',
		221437 => '1',
		221438 => '1',
		221439 => '1',
		221440 => '1',
		221441 => '1',
		221562 => '1',
		221563 => '1',
		221564 => '1',
		221565 => '1',
		221566 => '1',
		221687 => '1',
		221688 => '1',
		221689 => '1',
		221690 => '1',
		221691 => '1',
		222336 => '1',
		222337 => '1',
		222338 => '1',
		222339 => '1',
		222340 => '1',
		222461 => '1',
		222462 => '1',
		222463 => '1',
		222464 => '1',
		222465 => '1',
		222586 => '1',
		222587 => '1',
		222588 => '1',
		222589 => '1',
		222590 => '1',
		222711 => '1',
		222712 => '1',
		222713 => '1',
		222714 => '1',
		222715 => '1',
		223360 => '1',
		223361 => '1',
		223362 => '1',
		223363 => '1',
		223364 => '1',
		223485 => '1',
		223486 => '1',
		223487 => '1',
		223488 => '1',
		223489 => '1',
		223610 => '1',
		223611 => '1',
		223612 => '1',
		223613 => '1',
		223614 => '1',
		223735 => '1',
		223736 => '1',
		223737 => '1',
		223738 => '1',
		223739 => '1',
		224384 => '1',
		224385 => '1',
		224386 => '1',
		224387 => '1',
		224388 => '1',
		224509 => '1',
		224510 => '1',
		224511 => '1',
		224512 => '1',
		224513 => '1',
		224634 => '1',
		224635 => '1',
		224636 => '1',
		224637 => '1',
		224638 => '1',
		224759 => '1',
		224760 => '1',
		224761 => '1',
		224762 => '1',
		224763 => '1',
		225408 => '1',
		225409 => '1',
		225410 => '1',
		225411 => '1',
		225412 => '1',
		225533 => '1',
		225534 => '1',
		225535 => '1',
		225536 => '1',
		225537 => '1',
		225658 => '1',
		225659 => '1',
		225660 => '1',
		225661 => '1',
		225662 => '1',
		225783 => '1',
		225784 => '1',
		225785 => '1',
		225786 => '1',
		225787 => '1',
		226432 => '1',
		226433 => '1',
		226434 => '1',
		226435 => '1',
		226436 => '1',
		226557 => '1',
		226558 => '1',
		226559 => '1',
		226560 => '1',
		226561 => '1',
		226682 => '1',
		226683 => '1',
		226684 => '1',
		226685 => '1',
		226686 => '1',
		226807 => '1',
		226808 => '1',
		226809 => '1',
		226810 => '1',
		226811 => '1',
		227456 => '1',
		227457 => '1',
		227458 => '1',
		227459 => '1',
		227460 => '1',
		227581 => '1',
		227582 => '1',
		227583 => '1',
		227584 => '1',
		227585 => '1',
		227706 => '1',
		227707 => '1',
		227708 => '1',
		227709 => '1',
		227710 => '1',
		227831 => '1',
		227832 => '1',
		227833 => '1',
		227834 => '1',
		227835 => '1',
		228480 => '1',
		228481 => '1',
		228482 => '1',
		228483 => '1',
		228484 => '1',
		228605 => '1',
		228606 => '1',
		228607 => '1',
		228608 => '1',
		228609 => '1',
		228730 => '1',
		228731 => '1',
		228732 => '1',
		228733 => '1',
		228734 => '1',
		228855 => '1',
		228856 => '1',
		228857 => '1',
		228858 => '1',
		228859 => '1',
		229504 => '1',
		229505 => '1',
		229506 => '1',
		229507 => '1',
		229508 => '1',
		229629 => '1',
		229630 => '1',
		229631 => '1',
		229632 => '1',
		229633 => '1',
		229754 => '1',
		229755 => '1',
		229756 => '1',
		229757 => '1',
		229758 => '1',
		229879 => '1',
		229880 => '1',
		229881 => '1',
		229882 => '1',
		229883 => '1',
		230528 => '1',
		230529 => '1',
		230530 => '1',
		230531 => '1',
		230532 => '1',
		230653 => '1',
		230654 => '1',
		230655 => '1',
		230656 => '1',
		230657 => '1',
		230778 => '1',
		230779 => '1',
		230780 => '1',
		230781 => '1',
		230782 => '1',
		230903 => '1',
		230904 => '1',
		230905 => '1',
		230906 => '1',
		230907 => '1',
		231552 => '1',
		231553 => '1',
		231554 => '1',
		231555 => '1',
		231556 => '1',
		231677 => '1',
		231678 => '1',
		231679 => '1',
		231680 => '1',
		231681 => '1',
		231802 => '1',
		231803 => '1',
		231804 => '1',
		231805 => '1',
		231806 => '1',
		231927 => '1',
		231928 => '1',
		231929 => '1',
		231930 => '1',
		231931 => '1',
		232576 => '1',
		232577 => '1',
		232578 => '1',
		232579 => '1',
		232580 => '1',
		232701 => '1',
		232702 => '1',
		232703 => '1',
		232704 => '1',
		232705 => '1',
		232826 => '1',
		232827 => '1',
		232828 => '1',
		232829 => '1',
		232830 => '1',
		232951 => '1',
		232952 => '1',
		232953 => '1',
		232954 => '1',
		232955 => '1',
		233600 => '1',
		233601 => '1',
		233602 => '1',
		233603 => '1',
		233604 => '1',
		233725 => '1',
		233726 => '1',
		233727 => '1',
		233728 => '1',
		233729 => '1',
		233850 => '1',
		233851 => '1',
		233852 => '1',
		233853 => '1',
		233854 => '1',
		233975 => '1',
		233976 => '1',
		233977 => '1',
		233978 => '1',
		233979 => '1',
		234624 => '1',
		234625 => '1',
		234626 => '1',
		234627 => '1',
		234628 => '1',
		234749 => '1',
		234750 => '1',
		234751 => '1',
		234752 => '1',
		234753 => '1',
		234874 => '1',
		234875 => '1',
		234876 => '1',
		234877 => '1',
		234878 => '1',
		234999 => '1',
		235000 => '1',
		235001 => '1',
		235002 => '1',
		235003 => '1',
		235648 => '1',
		235649 => '1',
		235650 => '1',
		235651 => '1',
		235652 => '1',
		235773 => '1',
		235774 => '1',
		235775 => '1',
		235776 => '1',
		235777 => '1',
		235898 => '1',
		235899 => '1',
		235900 => '1',
		235901 => '1',
		235902 => '1',
		236023 => '1',
		236024 => '1',
		236025 => '1',
		236026 => '1',
		236027 => '1',
		236672 => '1',
		236673 => '1',
		236674 => '1',
		236675 => '1',
		236676 => '1',
		236797 => '1',
		236798 => '1',
		236799 => '1',
		236800 => '1',
		236801 => '1',
		236922 => '1',
		236923 => '1',
		236924 => '1',
		236925 => '1',
		236926 => '1',
		237047 => '1',
		237048 => '1',
		237049 => '1',
		237050 => '1',
		237051 => '1',
		237696 => '1',
		237697 => '1',
		237698 => '1',
		237699 => '1',
		237700 => '1',
		237821 => '1',
		237822 => '1',
		237823 => '1',
		237824 => '1',
		237825 => '1',
		237946 => '1',
		237947 => '1',
		237948 => '1',
		237949 => '1',
		237950 => '1',
		238071 => '1',
		238072 => '1',
		238073 => '1',
		238074 => '1',
		238075 => '1',
		238720 => '1',
		238721 => '1',
		238722 => '1',
		238723 => '1',
		238724 => '1',
		238845 => '1',
		238846 => '1',
		238847 => '1',
		238848 => '1',
		238849 => '1',
		238970 => '1',
		238971 => '1',
		238972 => '1',
		238973 => '1',
		238974 => '1',
		239095 => '1',
		239096 => '1',
		239097 => '1',
		239098 => '1',
		239099 => '1',
		239744 => '1',
		239745 => '1',
		239746 => '1',
		239747 => '1',
		239748 => '1',
		239869 => '1',
		239870 => '1',
		239871 => '1',
		239872 => '1',
		239873 => '1',
		239994 => '1',
		239995 => '1',
		239996 => '1',
		239997 => '1',
		239998 => '1',
		240119 => '1',
		240120 => '1',
		240121 => '1',
		240122 => '1',
		240123 => '1',
		240768 => '1',
		240769 => '1',
		240770 => '1',
		240771 => '1',
		240772 => '1',
		240893 => '1',
		240894 => '1',
		240895 => '1',
		240896 => '1',
		240897 => '1',
		241018 => '1',
		241019 => '1',
		241020 => '1',
		241021 => '1',
		241022 => '1',
		241143 => '1',
		241144 => '1',
		241145 => '1',
		241146 => '1',
		241147 => '1',
		241792 => '1',
		241793 => '1',
		241794 => '1',
		241795 => '1',
		241796 => '1',
		241917 => '1',
		241918 => '1',
		241919 => '1',
		241920 => '1',
		241921 => '1',
		242042 => '1',
		242043 => '1',
		242044 => '1',
		242045 => '1',
		242046 => '1',
		242167 => '1',
		242168 => '1',
		242169 => '1',
		242170 => '1',
		242171 => '1',
		242816 => '1',
		242817 => '1',
		242818 => '1',
		242819 => '1',
		242820 => '1',
		242941 => '1',
		242942 => '1',
		242943 => '1',
		242944 => '1',
		242945 => '1',
		243066 => '1',
		243067 => '1',
		243068 => '1',
		243069 => '1',
		243070 => '1',
		243191 => '1',
		243192 => '1',
		243193 => '1',
		243194 => '1',
		243195 => '1',
		243840 => '1',
		243841 => '1',
		243842 => '1',
		243843 => '1',
		243844 => '1',
		243965 => '1',
		243966 => '1',
		243967 => '1',
		243968 => '1',
		243969 => '1',
		244090 => '1',
		244091 => '1',
		244092 => '1',
		244093 => '1',
		244094 => '1',
		244215 => '1',
		244216 => '1',
		244217 => '1',
		244218 => '1',
		244219 => '1',
		244864 => '1',
		244865 => '1',
		244866 => '1',
		244867 => '1',
		244868 => '1',
		244989 => '1',
		244990 => '1',
		244991 => '1',
		244992 => '1',
		244993 => '1',
		245114 => '1',
		245115 => '1',
		245116 => '1',
		245117 => '1',
		245118 => '1',
		245239 => '1',
		245240 => '1',
		245241 => '1',
		245242 => '1',
		245243 => '1',
		245888 => '1',
		245889 => '1',
		245890 => '1',
		245891 => '1',
		245892 => '1',
		246013 => '1',
		246014 => '1',
		246015 => '1',
		246016 => '1',
		246017 => '1',
		246138 => '1',
		246139 => '1',
		246140 => '1',
		246141 => '1',
		246142 => '1',
		246263 => '1',
		246264 => '1',
		246265 => '1',
		246266 => '1',
		246267 => '1',
		246912 => '1',
		246913 => '1',
		246914 => '1',
		246915 => '1',
		246916 => '1',
		247037 => '1',
		247038 => '1',
		247039 => '1',
		247040 => '1',
		247041 => '1',
		247162 => '1',
		247163 => '1',
		247164 => '1',
		247165 => '1',
		247166 => '1',
		247287 => '1',
		247288 => '1',
		247289 => '1',
		247290 => '1',
		247291 => '1',
		247936 => '1',
		247937 => '1',
		247938 => '1',
		247939 => '1',
		247940 => '1',
		248061 => '1',
		248062 => '1',
		248063 => '1',
		248064 => '1',
		248065 => '1',
		248186 => '1',
		248187 => '1',
		248188 => '1',
		248189 => '1',
		248190 => '1',
		248311 => '1',
		248312 => '1',
		248313 => '1',
		248314 => '1',
		248315 => '1',
		248960 => '1',
		248961 => '1',
		248962 => '1',
		248963 => '1',
		248964 => '1',
		249085 => '1',
		249086 => '1',
		249087 => '1',
		249088 => '1',
		249089 => '1',
		249210 => '1',
		249211 => '1',
		249212 => '1',
		249213 => '1',
		249214 => '1',
		249335 => '1',
		249336 => '1',
		249337 => '1',
		249338 => '1',
		249339 => '1',
		249984 => '1',
		249985 => '1',
		249986 => '1',
		249987 => '1',
		249988 => '1',
		250109 => '1',
		250110 => '1',
		250111 => '1',
		250112 => '1',
		250113 => '1',
		250234 => '1',
		250235 => '1',
		250236 => '1',
		250237 => '1',
		250238 => '1',
		250359 => '1',
		250360 => '1',
		250361 => '1',
		250362 => '1',
		250363 => '1',
		251008 => '1',
		251009 => '1',
		251010 => '1',
		251011 => '1',
		251012 => '1',
		251133 => '1',
		251134 => '1',
		251135 => '1',
		251136 => '1',
		251137 => '1',
		251258 => '1',
		251259 => '1',
		251260 => '1',
		251261 => '1',
		251262 => '1',
		251383 => '1',
		251384 => '1',
		251385 => '1',
		251386 => '1',
		251387 => '1',
		252032 => '1',
		252033 => '1',
		252034 => '1',
		252035 => '1',
		252036 => '1',
		252157 => '1',
		252158 => '1',
		252159 => '1',
		252160 => '1',
		252161 => '1',
		252282 => '1',
		252283 => '1',
		252284 => '1',
		252285 => '1',
		252286 => '1',
		252407 => '1',
		252408 => '1',
		252409 => '1',
		252410 => '1',
		252411 => '1',
		253056 => '1',
		253057 => '1',
		253058 => '1',
		253059 => '1',
		253060 => '1',
		253181 => '1',
		253182 => '1',
		253183 => '1',
		253184 => '1',
		253185 => '1',
		253306 => '1',
		253307 => '1',
		253308 => '1',
		253309 => '1',
		253310 => '1',
		253431 => '1',
		253432 => '1',
		253433 => '1',
		253434 => '1',
		253435 => '1',
		254080 => '1',
		254081 => '1',
		254082 => '1',
		254083 => '1',
		254084 => '1',
		254205 => '1',
		254206 => '1',
		254207 => '1',
		254208 => '1',
		254209 => '1',
		254330 => '1',
		254331 => '1',
		254332 => '1',
		254333 => '1',
		254334 => '1',
		254455 => '1',
		254456 => '1',
		254457 => '1',
		254458 => '1',
		254459 => '1',
		255104 => '1',
		255105 => '1',
		255106 => '1',
		255107 => '1',
		255108 => '1',
		255229 => '1',
		255230 => '1',
		255231 => '1',
		255232 => '1',
		255233 => '1',
		255354 => '1',
		255355 => '1',
		255356 => '1',
		255357 => '1',
		255358 => '1',
		255479 => '1',
		255480 => '1',
		255481 => '1',
		255482 => '1',
		255483 => '1',
		256128 => '1',
		256129 => '1',
		256130 => '1',
		256131 => '1',
		256132 => '1',
		256253 => '1',
		256254 => '1',
		256255 => '1',
		256256 => '1',
		256257 => '1',
		256378 => '1',
		256379 => '1',
		256380 => '1',
		256381 => '1',
		256382 => '1',
		256503 => '1',
		256504 => '1',
		256505 => '1',
		256506 => '1',
		256507 => '1',
		257152 => '1',
		257153 => '1',
		257154 => '1',
		257155 => '1',
		257156 => '1',
		257277 => '1',
		257278 => '1',
		257279 => '1',
		257280 => '1',
		257281 => '1',
		257402 => '1',
		257403 => '1',
		257404 => '1',
		257405 => '1',
		257406 => '1',
		257527 => '1',
		257528 => '1',
		257529 => '1',
		257530 => '1',
		257531 => '1',
		258176 => '1',
		258177 => '1',
		258178 => '1',
		258179 => '1',
		258180 => '1',
		258301 => '1',
		258302 => '1',
		258303 => '1',
		258304 => '1',
		258305 => '1',
		258426 => '1',
		258427 => '1',
		258428 => '1',
		258429 => '1',
		258430 => '1',
		258551 => '1',
		258552 => '1',
		258553 => '1',
		258554 => '1',
		258555 => '1',
		259200 => '1',
		259201 => '1',
		259202 => '1',
		259203 => '1',
		259204 => '1',
		259325 => '1',
		259326 => '1',
		259327 => '1',
		259328 => '1',
		259329 => '1',
		259450 => '1',
		259451 => '1',
		259452 => '1',
		259453 => '1',
		259454 => '1',
		259575 => '1',
		259576 => '1',
		259577 => '1',
		259578 => '1',
		259579 => '1',
		260224 => '1',
		260225 => '1',
		260226 => '1',
		260227 => '1',
		260228 => '1',
		260349 => '1',
		260350 => '1',
		260351 => '1',
		260352 => '1',
		260353 => '1',
		260474 => '1',
		260475 => '1',
		260476 => '1',
		260477 => '1',
		260478 => '1',
		260599 => '1',
		260600 => '1',
		260601 => '1',
		260602 => '1',
		260603 => '1',
		261248 => '1',
		261249 => '1',
		261250 => '1',
		261251 => '1',
		261252 => '1',
		261373 => '1',
		261374 => '1',
		261375 => '1',
		261376 => '1',
		261377 => '1',
		261498 => '1',
		261499 => '1',
		261500 => '1',
		261501 => '1',
		261502 => '1',
		261623 => '1',
		261624 => '1',
		261625 => '1',
		261626 => '1',
		261627 => '1',
		262272 => '1',
		262273 => '1',
		262274 => '1',
		262275 => '1',
		262276 => '1',
		262397 => '1',
		262398 => '1',
		262399 => '1',
		262400 => '1',
		262401 => '1',
		262522 => '1',
		262523 => '1',
		262524 => '1',
		262525 => '1',
		262526 => '1',
		262647 => '1',
		262648 => '1',
		262649 => '1',
		262650 => '1',
		262651 => '1',
		263296 => '1',
		263297 => '1',
		263298 => '1',
		263299 => '1',
		263300 => '1',
		263421 => '1',
		263422 => '1',
		263423 => '1',
		263424 => '1',
		263425 => '1',
		263546 => '1',
		263547 => '1',
		263548 => '1',
		263549 => '1',
		263550 => '1',
		263671 => '1',
		263672 => '1',
		263673 => '1',
		263674 => '1',
		263675 => '1',
		264320 => '1',
		264321 => '1',
		264322 => '1',
		264323 => '1',
		264324 => '1',
		264445 => '1',
		264446 => '1',
		264447 => '1',
		264448 => '1',
		264449 => '1',
		264570 => '1',
		264571 => '1',
		264572 => '1',
		264573 => '1',
		264574 => '1',
		264695 => '1',
		264696 => '1',
		264697 => '1',
		264698 => '1',
		264699 => '1',
		265344 => '1',
		265345 => '1',
		265346 => '1',
		265347 => '1',
		265348 => '1',
		265469 => '1',
		265470 => '1',
		265471 => '1',
		265472 => '1',
		265473 => '1',
		265594 => '1',
		265595 => '1',
		265596 => '1',
		265597 => '1',
		265598 => '1',
		265719 => '1',
		265720 => '1',
		265721 => '1',
		265722 => '1',
		265723 => '1',
		266368 => '1',
		266369 => '1',
		266370 => '1',
		266371 => '1',
		266372 => '1',
		266493 => '1',
		266494 => '1',
		266495 => '1',
		266496 => '1',
		266497 => '1',
		266618 => '1',
		266619 => '1',
		266620 => '1',
		266621 => '1',
		266622 => '1',
		266743 => '1',
		266744 => '1',
		266745 => '1',
		266746 => '1',
		266747 => '1',
		267392 => '1',
		267393 => '1',
		267394 => '1',
		267395 => '1',
		267396 => '1',
		267517 => '1',
		267518 => '1',
		267519 => '1',
		267520 => '1',
		267521 => '1',
		267642 => '1',
		267643 => '1',
		267644 => '1',
		267645 => '1',
		267646 => '1',
		267767 => '1',
		267768 => '1',
		267769 => '1',
		267770 => '1',
		267771 => '1',
		268416 => '1',
		268417 => '1',
		268418 => '1',
		268419 => '1',
		268420 => '1',
		268541 => '1',
		268542 => '1',
		268543 => '1',
		268544 => '1',
		268545 => '1',
		268666 => '1',
		268667 => '1',
		268668 => '1',
		268669 => '1',
		268670 => '1',
		268791 => '1',
		268792 => '1',
		268793 => '1',
		268794 => '1',
		268795 => '1',
		269440 => '1',
		269441 => '1',
		269442 => '1',
		269443 => '1',
		269444 => '1',
		269565 => '1',
		269566 => '1',
		269567 => '1',
		269568 => '1',
		269569 => '1',
		269690 => '1',
		269691 => '1',
		269692 => '1',
		269693 => '1',
		269694 => '1',
		269815 => '1',
		269816 => '1',
		269817 => '1',
		269818 => '1',
		269819 => '1',
		270464 => '1',
		270465 => '1',
		270466 => '1',
		270467 => '1',
		270468 => '1',
		270589 => '1',
		270590 => '1',
		270591 => '1',
		270592 => '1',
		270593 => '1',
		270714 => '1',
		270715 => '1',
		270716 => '1',
		270717 => '1',
		270718 => '1',
		270839 => '1',
		270840 => '1',
		270841 => '1',
		270842 => '1',
		270843 => '1',
		271488 => '1',
		271489 => '1',
		271490 => '1',
		271491 => '1',
		271492 => '1',
		271613 => '1',
		271614 => '1',
		271615 => '1',
		271616 => '1',
		271617 => '1',
		271738 => '1',
		271739 => '1',
		271740 => '1',
		271741 => '1',
		271742 => '1',
		271863 => '1',
		271864 => '1',
		271865 => '1',
		271866 => '1',
		271867 => '1',
		272512 => '1',
		272513 => '1',
		272514 => '1',
		272515 => '1',
		272516 => '1',
		272637 => '1',
		272638 => '1',
		272639 => '1',
		272640 => '1',
		272641 => '1',
		272762 => '1',
		272763 => '1',
		272764 => '1',
		272765 => '1',
		272766 => '1',
		272887 => '1',
		272888 => '1',
		272889 => '1',
		272890 => '1',
		272891 => '1',
		273536 => '1',
		273537 => '1',
		273538 => '1',
		273539 => '1',
		273540 => '1',
		273661 => '1',
		273662 => '1',
		273663 => '1',
		273664 => '1',
		273665 => '1',
		273786 => '1',
		273787 => '1',
		273788 => '1',
		273789 => '1',
		273790 => '1',
		273911 => '1',
		273912 => '1',
		273913 => '1',
		273914 => '1',
		273915 => '1',
		274560 => '1',
		274561 => '1',
		274562 => '1',
		274563 => '1',
		274564 => '1',
		274685 => '1',
		274686 => '1',
		274687 => '1',
		274688 => '1',
		274689 => '1',
		274810 => '1',
		274811 => '1',
		274812 => '1',
		274813 => '1',
		274814 => '1',
		274935 => '1',
		274936 => '1',
		274937 => '1',
		274938 => '1',
		274939 => '1',
		275584 => '1',
		275585 => '1',
		275586 => '1',
		275587 => '1',
		275588 => '1',
		275709 => '1',
		275710 => '1',
		275711 => '1',
		275712 => '1',
		275713 => '1',
		275834 => '1',
		275835 => '1',
		275836 => '1',
		275837 => '1',
		275838 => '1',
		275959 => '1',
		275960 => '1',
		275961 => '1',
		275962 => '1',
		275963 => '1',
		276608 => '1',
		276609 => '1',
		276610 => '1',
		276611 => '1',
		276612 => '1',
		276733 => '1',
		276734 => '1',
		276735 => '1',
		276736 => '1',
		276737 => '1',
		276858 => '1',
		276859 => '1',
		276860 => '1',
		276861 => '1',
		276862 => '1',
		276983 => '1',
		276984 => '1',
		276985 => '1',
		276986 => '1',
		276987 => '1',
		277632 => '1',
		277633 => '1',
		277634 => '1',
		277635 => '1',
		277636 => '1',
		277757 => '1',
		277758 => '1',
		277759 => '1',
		277760 => '1',
		277761 => '1',
		277882 => '1',
		277883 => '1',
		277884 => '1',
		277885 => '1',
		277886 => '1',
		278007 => '1',
		278008 => '1',
		278009 => '1',
		278010 => '1',
		278011 => '1',
		278656 => '1',
		278657 => '1',
		278658 => '1',
		278659 => '1',
		278660 => '1',
		278781 => '1',
		278782 => '1',
		278783 => '1',
		278784 => '1',
		278785 => '1',
		278906 => '1',
		278907 => '1',
		278908 => '1',
		278909 => '1',
		278910 => '1',
		279031 => '1',
		279032 => '1',
		279033 => '1',
		279034 => '1',
		279035 => '1',
		279680 => '1',
		279681 => '1',
		279682 => '1',
		279683 => '1',
		279684 => '1',
		279805 => '1',
		279806 => '1',
		279807 => '1',
		279808 => '1',
		279809 => '1',
		279930 => '1',
		279931 => '1',
		279932 => '1',
		279933 => '1',
		279934 => '1',
		280055 => '1',
		280056 => '1',
		280057 => '1',
		280058 => '1',
		280059 => '1',
		280704 => '1',
		280705 => '1',
		280706 => '1',
		280707 => '1',
		280708 => '1',
		280829 => '1',
		280830 => '1',
		280831 => '1',
		280832 => '1',
		280833 => '1',
		280954 => '1',
		280955 => '1',
		280956 => '1',
		280957 => '1',
		280958 => '1',
		281079 => '1',
		281080 => '1',
		281081 => '1',
		281082 => '1',
		281083 => '1',
		281728 => '1',
		281729 => '1',
		281730 => '1',
		281731 => '1',
		281732 => '1',
		281853 => '1',
		281854 => '1',
		281855 => '1',
		281856 => '1',
		281857 => '1',
		281978 => '1',
		281979 => '1',
		281980 => '1',
		281981 => '1',
		281982 => '1',
		282103 => '1',
		282104 => '1',
		282105 => '1',
		282106 => '1',
		282107 => '1',
		282752 => '1',
		282753 => '1',
		282754 => '1',
		282755 => '1',
		282756 => '1',
		282877 => '1',
		282878 => '1',
		282879 => '1',
		282880 => '1',
		282881 => '1',
		283002 => '1',
		283003 => '1',
		283004 => '1',
		283005 => '1',
		283006 => '1',
		283127 => '1',
		283128 => '1',
		283129 => '1',
		283130 => '1',
		283131 => '1',
		283776 => '1',
		283777 => '1',
		283778 => '1',
		283779 => '1',
		283780 => '1',
		283901 => '1',
		283902 => '1',
		283903 => '1',
		283904 => '1',
		283905 => '1',
		284026 => '1',
		284027 => '1',
		284028 => '1',
		284029 => '1',
		284030 => '1',
		284151 => '1',
		284152 => '1',
		284153 => '1',
		284154 => '1',
		284155 => '1',
		284800 => '1',
		284801 => '1',
		284802 => '1',
		284803 => '1',
		284804 => '1',
		284925 => '1',
		284926 => '1',
		284927 => '1',
		284928 => '1',
		284929 => '1',
		285050 => '1',
		285051 => '1',
		285052 => '1',
		285053 => '1',
		285054 => '1',
		285175 => '1',
		285176 => '1',
		285177 => '1',
		285178 => '1',
		285179 => '1',
		285824 => '1',
		285825 => '1',
		285826 => '1',
		285827 => '1',
		285828 => '1',
		285949 => '1',
		285950 => '1',
		285951 => '1',
		285952 => '1',
		285953 => '1',
		286074 => '1',
		286075 => '1',
		286076 => '1',
		286077 => '1',
		286078 => '1',
		286199 => '1',
		286200 => '1',
		286201 => '1',
		286202 => '1',
		286203 => '1',
		286848 => '1',
		286849 => '1',
		286850 => '1',
		286851 => '1',
		286852 => '1',
		286973 => '1',
		286974 => '1',
		286975 => '1',
		286976 => '1',
		286977 => '1',
		287098 => '1',
		287099 => '1',
		287100 => '1',
		287101 => '1',
		287102 => '1',
		287223 => '1',
		287224 => '1',
		287225 => '1',
		287226 => '1',
		287227 => '1',
		287872 => '1',
		287873 => '1',
		287874 => '1',
		287875 => '1',
		287876 => '1',
		287997 => '1',
		287998 => '1',
		287999 => '1',
		288000 => '1',
		288001 => '1',
		288122 => '1',
		288123 => '1',
		288124 => '1',
		288125 => '1',
		288126 => '1',
		288247 => '1',
		288248 => '1',
		288249 => '1',
		288250 => '1',
		288251 => '1',
		288896 => '1',
		288897 => '1',
		288898 => '1',
		288899 => '1',
		288900 => '1',
		289021 => '1',
		289022 => '1',
		289023 => '1',
		289024 => '1',
		289025 => '1',
		289146 => '1',
		289147 => '1',
		289148 => '1',
		289149 => '1',
		289150 => '1',
		289271 => '1',
		289272 => '1',
		289273 => '1',
		289274 => '1',
		289275 => '1',
		289920 => '1',
		289921 => '1',
		289922 => '1',
		289923 => '1',
		289924 => '1',
		290045 => '1',
		290046 => '1',
		290047 => '1',
		290048 => '1',
		290049 => '1',
		290170 => '1',
		290171 => '1',
		290172 => '1',
		290173 => '1',
		290174 => '1',
		290295 => '1',
		290296 => '1',
		290297 => '1',
		290298 => '1',
		290299 => '1',
		290944 => '1',
		290945 => '1',
		290946 => '1',
		290947 => '1',
		290948 => '1',
		291069 => '1',
		291070 => '1',
		291071 => '1',
		291072 => '1',
		291073 => '1',
		291194 => '1',
		291195 => '1',
		291196 => '1',
		291197 => '1',
		291198 => '1',
		291319 => '1',
		291320 => '1',
		291321 => '1',
		291322 => '1',
		291323 => '1',
		291968 => '1',
		291969 => '1',
		291970 => '1',
		291971 => '1',
		291972 => '1',
		292093 => '1',
		292094 => '1',
		292095 => '1',
		292096 => '1',
		292097 => '1',
		292218 => '1',
		292219 => '1',
		292220 => '1',
		292221 => '1',
		292222 => '1',
		292343 => '1',
		292344 => '1',
		292345 => '1',
		292346 => '1',
		292347 => '1',
		292992 => '1',
		292993 => '1',
		292994 => '1',
		292995 => '1',
		292996 => '1',
		293117 => '1',
		293118 => '1',
		293119 => '1',
		293120 => '1',
		293121 => '1',
		293242 => '1',
		293243 => '1',
		293244 => '1',
		293245 => '1',
		293246 => '1',
		293367 => '1',
		293368 => '1',
		293369 => '1',
		293370 => '1',
		293371 => '1',
		294016 => '1',
		294017 => '1',
		294018 => '1',
		294019 => '1',
		294020 => '1',
		294141 => '1',
		294142 => '1',
		294143 => '1',
		294144 => '1',
		294145 => '1',
		294266 => '1',
		294267 => '1',
		294268 => '1',
		294269 => '1',
		294270 => '1',
		294391 => '1',
		294392 => '1',
		294393 => '1',
		294394 => '1',
		294395 => '1',
		295040 => '1',
		295041 => '1',
		295042 => '1',
		295043 => '1',
		295044 => '1',
		295165 => '1',
		295166 => '1',
		295167 => '1',
		295168 => '1',
		295169 => '1',
		295290 => '1',
		295291 => '1',
		295292 => '1',
		295293 => '1',
		295294 => '1',
		295415 => '1',
		295416 => '1',
		295417 => '1',
		295418 => '1',
		295419 => '1',
		296064 => '1',
		296065 => '1',
		296066 => '1',
		296067 => '1',
		296068 => '1',
		296189 => '1',
		296190 => '1',
		296191 => '1',
		296192 => '1',
		296193 => '1',
		296314 => '1',
		296315 => '1',
		296316 => '1',
		296317 => '1',
		296318 => '1',
		296439 => '1',
		296440 => '1',
		296441 => '1',
		296442 => '1',
		296443 => '1',
		297088 => '1',
		297089 => '1',
		297090 => '1',
		297091 => '1',
		297092 => '1',
		297213 => '1',
		297214 => '1',
		297215 => '1',
		297216 => '1',
		297217 => '1',
		297338 => '1',
		297339 => '1',
		297340 => '1',
		297341 => '1',
		297342 => '1',
		297463 => '1',
		297464 => '1',
		297465 => '1',
		297466 => '1',
		297467 => '1',
		298112 => '1',
		298113 => '1',
		298114 => '1',
		298115 => '1',
		298116 => '1',
		298237 => '1',
		298238 => '1',
		298239 => '1',
		298240 => '1',
		298241 => '1',
		298362 => '1',
		298363 => '1',
		298364 => '1',
		298365 => '1',
		298366 => '1',
		298487 => '1',
		298488 => '1',
		298489 => '1',
		298490 => '1',
		298491 => '1',
		299136 => '1',
		299137 => '1',
		299138 => '1',
		299139 => '1',
		299140 => '1',
		299261 => '1',
		299262 => '1',
		299263 => '1',
		299264 => '1',
		299265 => '1',
		299386 => '1',
		299387 => '1',
		299388 => '1',
		299389 => '1',
		299390 => '1',
		299511 => '1',
		299512 => '1',
		299513 => '1',
		299514 => '1',
		299515 => '1',
		300160 => '1',
		300161 => '1',
		300162 => '1',
		300163 => '1',
		300164 => '1',
		300285 => '1',
		300286 => '1',
		300287 => '1',
		300288 => '1',
		300289 => '1',
		300410 => '1',
		300411 => '1',
		300412 => '1',
		300413 => '1',
		300414 => '1',
		300535 => '1',
		300536 => '1',
		300537 => '1',
		300538 => '1',
		300539 => '1',
		301184 => '1',
		301185 => '1',
		301186 => '1',
		301187 => '1',
		301188 => '1',
		301309 => '1',
		301310 => '1',
		301311 => '1',
		301312 => '1',
		301313 => '1',
		301434 => '1',
		301435 => '1',
		301436 => '1',
		301437 => '1',
		301438 => '1',
		301559 => '1',
		301560 => '1',
		301561 => '1',
		301562 => '1',
		301563 => '1',
		302208 => '1',
		302209 => '1',
		302210 => '1',
		302211 => '1',
		302212 => '1',
		302333 => '1',
		302334 => '1',
		302335 => '1',
		302336 => '1',
		302337 => '1',
		302458 => '1',
		302459 => '1',
		302460 => '1',
		302461 => '1',
		302462 => '1',
		302583 => '1',
		302584 => '1',
		302585 => '1',
		302586 => '1',
		302587 => '1',
		303232 => '1',
		303233 => '1',
		303234 => '1',
		303235 => '1',
		303236 => '1',
		303357 => '1',
		303358 => '1',
		303359 => '1',
		303360 => '1',
		303361 => '1',
		303482 => '1',
		303483 => '1',
		303484 => '1',
		303485 => '1',
		303486 => '1',
		303607 => '1',
		303608 => '1',
		303609 => '1',
		303610 => '1',
		303611 => '1',
		304256 => '1',
		304257 => '1',
		304258 => '1',
		304259 => '1',
		304260 => '1',
		304381 => '1',
		304382 => '1',
		304383 => '1',
		304384 => '1',
		304385 => '1',
		304506 => '1',
		304507 => '1',
		304508 => '1',
		304509 => '1',
		304510 => '1',
		304631 => '1',
		304632 => '1',
		304633 => '1',
		304634 => '1',
		304635 => '1',
		305280 => '1',
		305281 => '1',
		305282 => '1',
		305283 => '1',
		305284 => '1',
		305285 => '1',
		305286 => '1',
		305287 => '1',
		305288 => '1',
		305289 => '1',
		305290 => '1',
		305291 => '1',
		305292 => '1',
		305293 => '1',
		305294 => '1',
		305295 => '1',
		305296 => '1',
		305297 => '1',
		305298 => '1',
		305299 => '1',
		305300 => '1',
		305301 => '1',
		305302 => '1',
		305303 => '1',
		305304 => '1',
		305305 => '1',
		305306 => '1',
		305307 => '1',
		305308 => '1',
		305309 => '1',
		305310 => '1',
		305311 => '1',
		305312 => '1',
		305313 => '1',
		305314 => '1',
		305315 => '1',
		305316 => '1',
		305317 => '1',
		305318 => '1',
		305319 => '1',
		305320 => '1',
		305321 => '1',
		305322 => '1',
		305323 => '1',
		305324 => '1',
		305325 => '1',
		305326 => '1',
		305327 => '1',
		305328 => '1',
		305329 => '1',
		305330 => '1',
		305331 => '1',
		305332 => '1',
		305333 => '1',
		305334 => '1',
		305335 => '1',
		305336 => '1',
		305337 => '1',
		305338 => '1',
		305339 => '1',
		305340 => '1',
		305341 => '1',
		305342 => '1',
		305343 => '1',
		305344 => '1',
		305345 => '1',
		305346 => '1',
		305347 => '1',
		305348 => '1',
		305349 => '1',
		305350 => '1',
		305351 => '1',
		305352 => '1',
		305353 => '1',
		305354 => '1',
		305355 => '1',
		305356 => '1',
		305357 => '1',
		305358 => '1',
		305359 => '1',
		305360 => '1',
		305361 => '1',
		305362 => '1',
		305363 => '1',
		305364 => '1',
		305365 => '1',
		305366 => '1',
		305367 => '1',
		305368 => '1',
		305369 => '1',
		305370 => '1',
		305371 => '1',
		305372 => '1',
		305373 => '1',
		305374 => '1',
		305375 => '1',
		305376 => '1',
		305377 => '1',
		305378 => '1',
		305379 => '1',
		305380 => '1',
		305381 => '1',
		305382 => '1',
		305383 => '1',
		305384 => '1',
		305385 => '1',
		305386 => '1',
		305387 => '1',
		305388 => '1',
		305389 => '1',
		305390 => '1',
		305391 => '1',
		305392 => '1',
		305393 => '1',
		305394 => '1',
		305395 => '1',
		305396 => '1',
		305397 => '1',
		305398 => '1',
		305399 => '1',
		305400 => '1',
		305401 => '1',
		305402 => '1',
		305403 => '1',
		305404 => '1',
		305405 => '1',
		305406 => '1',
		305407 => '1',
		305408 => '1',
		305409 => '1',
		305410 => '1',
		305411 => '1',
		305412 => '1',
		305413 => '1',
		305414 => '1',
		305415 => '1',
		305416 => '1',
		305417 => '1',
		305418 => '1',
		305419 => '1',
		305420 => '1',
		305421 => '1',
		305422 => '1',
		305423 => '1',
		305424 => '1',
		305425 => '1',
		305426 => '1',
		305427 => '1',
		305428 => '1',
		305429 => '1',
		305430 => '1',
		305431 => '1',
		305432 => '1',
		305433 => '1',
		305434 => '1',
		305435 => '1',
		305436 => '1',
		305437 => '1',
		305438 => '1',
		305439 => '1',
		305440 => '1',
		305441 => '1',
		305442 => '1',
		305443 => '1',
		305444 => '1',
		305445 => '1',
		305446 => '1',
		305447 => '1',
		305448 => '1',
		305449 => '1',
		305450 => '1',
		305451 => '1',
		305452 => '1',
		305453 => '1',
		305454 => '1',
		305455 => '1',
		305456 => '1',
		305457 => '1',
		305458 => '1',
		305459 => '1',
		305460 => '1',
		305461 => '1',
		305462 => '1',
		305463 => '1',
		305464 => '1',
		305465 => '1',
		305466 => '1',
		305467 => '1',
		305468 => '1',
		305469 => '1',
		305470 => '1',
		305471 => '1',
		305472 => '1',
		305473 => '1',
		305474 => '1',
		305475 => '1',
		305476 => '1',
		305477 => '1',
		305478 => '1',
		305479 => '1',
		305480 => '1',
		305481 => '1',
		305482 => '1',
		305483 => '1',
		305484 => '1',
		305485 => '1',
		305486 => '1',
		305487 => '1',
		305488 => '1',
		305489 => '1',
		305490 => '1',
		305491 => '1',
		305492 => '1',
		305493 => '1',
		305494 => '1',
		305495 => '1',
		305496 => '1',
		305497 => '1',
		305498 => '1',
		305499 => '1',
		305500 => '1',
		305501 => '1',
		305502 => '1',
		305503 => '1',
		305504 => '1',
		305505 => '1',
		305506 => '1',
		305507 => '1',
		305508 => '1',
		305509 => '1',
		305510 => '1',
		305511 => '1',
		305512 => '1',
		305513 => '1',
		305514 => '1',
		305515 => '1',
		305516 => '1',
		305517 => '1',
		305518 => '1',
		305519 => '1',
		305520 => '1',
		305521 => '1',
		305522 => '1',
		305523 => '1',
		305524 => '1',
		305525 => '1',
		305526 => '1',
		305527 => '1',
		305528 => '1',
		305529 => '1',
		305530 => '1',
		305531 => '1',
		305532 => '1',
		305533 => '1',
		305534 => '1',
		305535 => '1',
		305536 => '1',
		305537 => '1',
		305538 => '1',
		305539 => '1',
		305540 => '1',
		305541 => '1',
		305542 => '1',
		305543 => '1',
		305544 => '1',
		305545 => '1',
		305546 => '1',
		305547 => '1',
		305548 => '1',
		305549 => '1',
		305550 => '1',
		305551 => '1',
		305552 => '1',
		305553 => '1',
		305554 => '1',
		305555 => '1',
		305556 => '1',
		305557 => '1',
		305558 => '1',
		305559 => '1',
		305560 => '1',
		305561 => '1',
		305562 => '1',
		305563 => '1',
		305564 => '1',
		305565 => '1',
		305566 => '1',
		305567 => '1',
		305568 => '1',
		305569 => '1',
		305570 => '1',
		305571 => '1',
		305572 => '1',
		305573 => '1',
		305574 => '1',
		305575 => '1',
		305576 => '1',
		305577 => '1',
		305578 => '1',
		305579 => '1',
		305580 => '1',
		305581 => '1',
		305582 => '1',
		305583 => '1',
		305584 => '1',
		305585 => '1',
		305586 => '1',
		305587 => '1',
		305588 => '1',
		305589 => '1',
		305590 => '1',
		305591 => '1',
		305592 => '1',
		305593 => '1',
		305594 => '1',
		305595 => '1',
		305596 => '1',
		305597 => '1',
		305598 => '1',
		305599 => '1',
		305600 => '1',
		305601 => '1',
		305602 => '1',
		305603 => '1',
		305604 => '1',
		305605 => '1',
		305606 => '1',
		305607 => '1',
		305608 => '1',
		305609 => '1',
		305610 => '1',
		305611 => '1',
		305612 => '1',
		305613 => '1',
		305614 => '1',
		305615 => '1',
		305616 => '1',
		305617 => '1',
		305618 => '1',
		305619 => '1',
		305620 => '1',
		305621 => '1',
		305622 => '1',
		305623 => '1',
		305624 => '1',
		305625 => '1',
		305626 => '1',
		305627 => '1',
		305628 => '1',
		305629 => '1',
		305630 => '1',
		305631 => '1',
		305632 => '1',
		305633 => '1',
		305634 => '1',
		305635 => '1',
		305636 => '1',
		305637 => '1',
		305638 => '1',
		305639 => '1',
		305640 => '1',
		305641 => '1',
		305642 => '1',
		305643 => '1',
		305644 => '1',
		305645 => '1',
		305646 => '1',
		305647 => '1',
		305648 => '1',
		305649 => '1',
		305650 => '1',
		305651 => '1',
		305652 => '1',
		305653 => '1',
		305654 => '1',
		305655 => '1',
		305656 => '1',
		305657 => '1',
		305658 => '1',
		305659 => '1',
		306304 => '1',
		306305 => '1',
		306306 => '1',
		306307 => '1',
		306308 => '1',
		306309 => '1',
		306310 => '1',
		306311 => '1',
		306312 => '1',
		306313 => '1',
		306314 => '1',
		306315 => '1',
		306316 => '1',
		306317 => '1',
		306318 => '1',
		306319 => '1',
		306320 => '1',
		306321 => '1',
		306322 => '1',
		306323 => '1',
		306324 => '1',
		306325 => '1',
		306326 => '1',
		306327 => '1',
		306328 => '1',
		306329 => '1',
		306330 => '1',
		306331 => '1',
		306332 => '1',
		306333 => '1',
		306334 => '1',
		306335 => '1',
		306336 => '1',
		306337 => '1',
		306338 => '1',
		306339 => '1',
		306340 => '1',
		306341 => '1',
		306342 => '1',
		306343 => '1',
		306344 => '1',
		306345 => '1',
		306346 => '1',
		306347 => '1',
		306348 => '1',
		306349 => '1',
		306350 => '1',
		306351 => '1',
		306352 => '1',
		306353 => '1',
		306354 => '1',
		306355 => '1',
		306356 => '1',
		306357 => '1',
		306358 => '1',
		306359 => '1',
		306360 => '1',
		306361 => '1',
		306362 => '1',
		306363 => '1',
		306364 => '1',
		306365 => '1',
		306366 => '1',
		306367 => '1',
		306368 => '1',
		306369 => '1',
		306370 => '1',
		306371 => '1',
		306372 => '1',
		306373 => '1',
		306374 => '1',
		306375 => '1',
		306376 => '1',
		306377 => '1',
		306378 => '1',
		306379 => '1',
		306380 => '1',
		306381 => '1',
		306382 => '1',
		306383 => '1',
		306384 => '1',
		306385 => '1',
		306386 => '1',
		306387 => '1',
		306388 => '1',
		306389 => '1',
		306390 => '1',
		306391 => '1',
		306392 => '1',
		306393 => '1',
		306394 => '1',
		306395 => '1',
		306396 => '1',
		306397 => '1',
		306398 => '1',
		306399 => '1',
		306400 => '1',
		306401 => '1',
		306402 => '1',
		306403 => '1',
		306404 => '1',
		306405 => '1',
		306406 => '1',
		306407 => '1',
		306408 => '1',
		306409 => '1',
		306410 => '1',
		306411 => '1',
		306412 => '1',
		306413 => '1',
		306414 => '1',
		306415 => '1',
		306416 => '1',
		306417 => '1',
		306418 => '1',
		306419 => '1',
		306420 => '1',
		306421 => '1',
		306422 => '1',
		306423 => '1',
		306424 => '1',
		306425 => '1',
		306426 => '1',
		306427 => '1',
		306428 => '1',
		306429 => '1',
		306430 => '1',
		306431 => '1',
		306432 => '1',
		306433 => '1',
		306434 => '1',
		306435 => '1',
		306436 => '1',
		306437 => '1',
		306438 => '1',
		306439 => '1',
		306440 => '1',
		306441 => '1',
		306442 => '1',
		306443 => '1',
		306444 => '1',
		306445 => '1',
		306446 => '1',
		306447 => '1',
		306448 => '1',
		306449 => '1',
		306450 => '1',
		306451 => '1',
		306452 => '1',
		306453 => '1',
		306454 => '1',
		306455 => '1',
		306456 => '1',
		306457 => '1',
		306458 => '1',
		306459 => '1',
		306460 => '1',
		306461 => '1',
		306462 => '1',
		306463 => '1',
		306464 => '1',
		306465 => '1',
		306466 => '1',
		306467 => '1',
		306468 => '1',
		306469 => '1',
		306470 => '1',
		306471 => '1',
		306472 => '1',
		306473 => '1',
		306474 => '1',
		306475 => '1',
		306476 => '1',
		306477 => '1',
		306478 => '1',
		306479 => '1',
		306480 => '1',
		306481 => '1',
		306482 => '1',
		306483 => '1',
		306484 => '1',
		306485 => '1',
		306486 => '1',
		306487 => '1',
		306488 => '1',
		306489 => '1',
		306490 => '1',
		306491 => '1',
		306492 => '1',
		306493 => '1',
		306494 => '1',
		306495 => '1',
		306496 => '1',
		306497 => '1',
		306498 => '1',
		306499 => '1',
		306500 => '1',
		306501 => '1',
		306502 => '1',
		306503 => '1',
		306504 => '1',
		306505 => '1',
		306506 => '1',
		306507 => '1',
		306508 => '1',
		306509 => '1',
		306510 => '1',
		306511 => '1',
		306512 => '1',
		306513 => '1',
		306514 => '1',
		306515 => '1',
		306516 => '1',
		306517 => '1',
		306518 => '1',
		306519 => '1',
		306520 => '1',
		306521 => '1',
		306522 => '1',
		306523 => '1',
		306524 => '1',
		306525 => '1',
		306526 => '1',
		306527 => '1',
		306528 => '1',
		306529 => '1',
		306530 => '1',
		306531 => '1',
		306532 => '1',
		306533 => '1',
		306534 => '1',
		306535 => '1',
		306536 => '1',
		306537 => '1',
		306538 => '1',
		306539 => '1',
		306540 => '1',
		306541 => '1',
		306542 => '1',
		306543 => '1',
		306544 => '1',
		306545 => '1',
		306546 => '1',
		306547 => '1',
		306548 => '1',
		306549 => '1',
		306550 => '1',
		306551 => '1',
		306552 => '1',
		306553 => '1',
		306554 => '1',
		306555 => '1',
		306556 => '1',
		306557 => '1',
		306558 => '1',
		306559 => '1',
		306560 => '1',
		306561 => '1',
		306562 => '1',
		306563 => '1',
		306564 => '1',
		306565 => '1',
		306566 => '1',
		306567 => '1',
		306568 => '1',
		306569 => '1',
		306570 => '1',
		306571 => '1',
		306572 => '1',
		306573 => '1',
		306574 => '1',
		306575 => '1',
		306576 => '1',
		306577 => '1',
		306578 => '1',
		306579 => '1',
		306580 => '1',
		306581 => '1',
		306582 => '1',
		306583 => '1',
		306584 => '1',
		306585 => '1',
		306586 => '1',
		306587 => '1',
		306588 => '1',
		306589 => '1',
		306590 => '1',
		306591 => '1',
		306592 => '1',
		306593 => '1',
		306594 => '1',
		306595 => '1',
		306596 => '1',
		306597 => '1',
		306598 => '1',
		306599 => '1',
		306600 => '1',
		306601 => '1',
		306602 => '1',
		306603 => '1',
		306604 => '1',
		306605 => '1',
		306606 => '1',
		306607 => '1',
		306608 => '1',
		306609 => '1',
		306610 => '1',
		306611 => '1',
		306612 => '1',
		306613 => '1',
		306614 => '1',
		306615 => '1',
		306616 => '1',
		306617 => '1',
		306618 => '1',
		306619 => '1',
		306620 => '1',
		306621 => '1',
		306622 => '1',
		306623 => '1',
		306624 => '1',
		306625 => '1',
		306626 => '1',
		306627 => '1',
		306628 => '1',
		306629 => '1',
		306630 => '1',
		306631 => '1',
		306632 => '1',
		306633 => '1',
		306634 => '1',
		306635 => '1',
		306636 => '1',
		306637 => '1',
		306638 => '1',
		306639 => '1',
		306640 => '1',
		306641 => '1',
		306642 => '1',
		306643 => '1',
		306644 => '1',
		306645 => '1',
		306646 => '1',
		306647 => '1',
		306648 => '1',
		306649 => '1',
		306650 => '1',
		306651 => '1',
		306652 => '1',
		306653 => '1',
		306654 => '1',
		306655 => '1',
		306656 => '1',
		306657 => '1',
		306658 => '1',
		306659 => '1',
		306660 => '1',
		306661 => '1',
		306662 => '1',
		306663 => '1',
		306664 => '1',
		306665 => '1',
		306666 => '1',
		306667 => '1',
		306668 => '1',
		306669 => '1',
		306670 => '1',
		306671 => '1',
		306672 => '1',
		306673 => '1',
		306674 => '1',
		306675 => '1',
		306676 => '1',
		306677 => '1',
		306678 => '1',
		306679 => '1',
		306680 => '1',
		306681 => '1',
		306682 => '1',
		306683 => '1',
		307328 => '1',
		307329 => '1',
		307330 => '1',
		307331 => '1',
		307332 => '1',
		307333 => '1',
		307334 => '1',
		307335 => '1',
		307336 => '1',
		307337 => '1',
		307338 => '1',
		307339 => '1',
		307340 => '1',
		307341 => '1',
		307342 => '1',
		307343 => '1',
		307344 => '1',
		307345 => '1',
		307346 => '1',
		307347 => '1',
		307348 => '1',
		307349 => '1',
		307350 => '1',
		307351 => '1',
		307352 => '1',
		307353 => '1',
		307354 => '1',
		307355 => '1',
		307356 => '1',
		307357 => '1',
		307358 => '1',
		307359 => '1',
		307360 => '1',
		307361 => '1',
		307362 => '1',
		307363 => '1',
		307364 => '1',
		307365 => '1',
		307366 => '1',
		307367 => '1',
		307368 => '1',
		307369 => '1',
		307370 => '1',
		307371 => '1',
		307372 => '1',
		307373 => '1',
		307374 => '1',
		307375 => '1',
		307376 => '1',
		307377 => '1',
		307378 => '1',
		307379 => '1',
		307380 => '1',
		307381 => '1',
		307382 => '1',
		307383 => '1',
		307384 => '1',
		307385 => '1',
		307386 => '1',
		307387 => '1',
		307388 => '1',
		307389 => '1',
		307390 => '1',
		307391 => '1',
		307392 => '1',
		307393 => '1',
		307394 => '1',
		307395 => '1',
		307396 => '1',
		307397 => '1',
		307398 => '1',
		307399 => '1',
		307400 => '1',
		307401 => '1',
		307402 => '1',
		307403 => '1',
		307404 => '1',
		307405 => '1',
		307406 => '1',
		307407 => '1',
		307408 => '1',
		307409 => '1',
		307410 => '1',
		307411 => '1',
		307412 => '1',
		307413 => '1',
		307414 => '1',
		307415 => '1',
		307416 => '1',
		307417 => '1',
		307418 => '1',
		307419 => '1',
		307420 => '1',
		307421 => '1',
		307422 => '1',
		307423 => '1',
		307424 => '1',
		307425 => '1',
		307426 => '1',
		307427 => '1',
		307428 => '1',
		307429 => '1',
		307430 => '1',
		307431 => '1',
		307432 => '1',
		307433 => '1',
		307434 => '1',
		307435 => '1',
		307436 => '1',
		307437 => '1',
		307438 => '1',
		307439 => '1',
		307440 => '1',
		307441 => '1',
		307442 => '1',
		307443 => '1',
		307444 => '1',
		307445 => '1',
		307446 => '1',
		307447 => '1',
		307448 => '1',
		307449 => '1',
		307450 => '1',
		307451 => '1',
		307452 => '1',
		307453 => '1',
		307454 => '1',
		307455 => '1',
		307456 => '1',
		307457 => '1',
		307458 => '1',
		307459 => '1',
		307460 => '1',
		307461 => '1',
		307462 => '1',
		307463 => '1',
		307464 => '1',
		307465 => '1',
		307466 => '1',
		307467 => '1',
		307468 => '1',
		307469 => '1',
		307470 => '1',
		307471 => '1',
		307472 => '1',
		307473 => '1',
		307474 => '1',
		307475 => '1',
		307476 => '1',
		307477 => '1',
		307478 => '1',
		307479 => '1',
		307480 => '1',
		307481 => '1',
		307482 => '1',
		307483 => '1',
		307484 => '1',
		307485 => '1',
		307486 => '1',
		307487 => '1',
		307488 => '1',
		307489 => '1',
		307490 => '1',
		307491 => '1',
		307492 => '1',
		307493 => '1',
		307494 => '1',
		307495 => '1',
		307496 => '1',
		307497 => '1',
		307498 => '1',
		307499 => '1',
		307500 => '1',
		307501 => '1',
		307502 => '1',
		307503 => '1',
		307504 => '1',
		307505 => '1',
		307506 => '1',
		307507 => '1',
		307508 => '1',
		307509 => '1',
		307510 => '1',
		307511 => '1',
		307512 => '1',
		307513 => '1',
		307514 => '1',
		307515 => '1',
		307516 => '1',
		307517 => '1',
		307518 => '1',
		307519 => '1',
		307520 => '1',
		307521 => '1',
		307522 => '1',
		307523 => '1',
		307524 => '1',
		307525 => '1',
		307526 => '1',
		307527 => '1',
		307528 => '1',
		307529 => '1',
		307530 => '1',
		307531 => '1',
		307532 => '1',
		307533 => '1',
		307534 => '1',
		307535 => '1',
		307536 => '1',
		307537 => '1',
		307538 => '1',
		307539 => '1',
		307540 => '1',
		307541 => '1',
		307542 => '1',
		307543 => '1',
		307544 => '1',
		307545 => '1',
		307546 => '1',
		307547 => '1',
		307548 => '1',
		307549 => '1',
		307550 => '1',
		307551 => '1',
		307552 => '1',
		307553 => '1',
		307554 => '1',
		307555 => '1',
		307556 => '1',
		307557 => '1',
		307558 => '1',
		307559 => '1',
		307560 => '1',
		307561 => '1',
		307562 => '1',
		307563 => '1',
		307564 => '1',
		307565 => '1',
		307566 => '1',
		307567 => '1',
		307568 => '1',
		307569 => '1',
		307570 => '1',
		307571 => '1',
		307572 => '1',
		307573 => '1',
		307574 => '1',
		307575 => '1',
		307576 => '1',
		307577 => '1',
		307578 => '1',
		307579 => '1',
		307580 => '1',
		307581 => '1',
		307582 => '1',
		307583 => '1',
		307584 => '1',
		307585 => '1',
		307586 => '1',
		307587 => '1',
		307588 => '1',
		307589 => '1',
		307590 => '1',
		307591 => '1',
		307592 => '1',
		307593 => '1',
		307594 => '1',
		307595 => '1',
		307596 => '1',
		307597 => '1',
		307598 => '1',
		307599 => '1',
		307600 => '1',
		307601 => '1',
		307602 => '1',
		307603 => '1',
		307604 => '1',
		307605 => '1',
		307606 => '1',
		307607 => '1',
		307608 => '1',
		307609 => '1',
		307610 => '1',
		307611 => '1',
		307612 => '1',
		307613 => '1',
		307614 => '1',
		307615 => '1',
		307616 => '1',
		307617 => '1',
		307618 => '1',
		307619 => '1',
		307620 => '1',
		307621 => '1',
		307622 => '1',
		307623 => '1',
		307624 => '1',
		307625 => '1',
		307626 => '1',
		307627 => '1',
		307628 => '1',
		307629 => '1',
		307630 => '1',
		307631 => '1',
		307632 => '1',
		307633 => '1',
		307634 => '1',
		307635 => '1',
		307636 => '1',
		307637 => '1',
		307638 => '1',
		307639 => '1',
		307640 => '1',
		307641 => '1',
		307642 => '1',
		307643 => '1',
		307644 => '1',
		307645 => '1',
		307646 => '1',
		307647 => '1',
		307648 => '1',
		307649 => '1',
		307650 => '1',
		307651 => '1',
		307652 => '1',
		307653 => '1',
		307654 => '1',
		307655 => '1',
		307656 => '1',
		307657 => '1',
		307658 => '1',
		307659 => '1',
		307660 => '1',
		307661 => '1',
		307662 => '1',
		307663 => '1',
		307664 => '1',
		307665 => '1',
		307666 => '1',
		307667 => '1',
		307668 => '1',
		307669 => '1',
		307670 => '1',
		307671 => '1',
		307672 => '1',
		307673 => '1',
		307674 => '1',
		307675 => '1',
		307676 => '1',
		307677 => '1',
		307678 => '1',
		307679 => '1',
		307680 => '1',
		307681 => '1',
		307682 => '1',
		307683 => '1',
		307684 => '1',
		307685 => '1',
		307686 => '1',
		307687 => '1',
		307688 => '1',
		307689 => '1',
		307690 => '1',
		307691 => '1',
		307692 => '1',
		307693 => '1',
		307694 => '1',
		307695 => '1',
		307696 => '1',
		307697 => '1',
		307698 => '1',
		307699 => '1',
		307700 => '1',
		307701 => '1',
		307702 => '1',
		307703 => '1',
		307704 => '1',
		307705 => '1',
		307706 => '1',
		307707 => '1',
		308352 => '1',
		308353 => '1',
		308354 => '1',
		308355 => '1',
		308356 => '1',
		308357 => '1',
		308358 => '1',
		308359 => '1',
		308360 => '1',
		308361 => '1',
		308362 => '1',
		308363 => '1',
		308364 => '1',
		308365 => '1',
		308366 => '1',
		308367 => '1',
		308368 => '1',
		308369 => '1',
		308370 => '1',
		308371 => '1',
		308372 => '1',
		308373 => '1',
		308374 => '1',
		308375 => '1',
		308376 => '1',
		308377 => '1',
		308378 => '1',
		308379 => '1',
		308380 => '1',
		308381 => '1',
		308382 => '1',
		308383 => '1',
		308384 => '1',
		308385 => '1',
		308386 => '1',
		308387 => '1',
		308388 => '1',
		308389 => '1',
		308390 => '1',
		308391 => '1',
		308392 => '1',
		308393 => '1',
		308394 => '1',
		308395 => '1',
		308396 => '1',
		308397 => '1',
		308398 => '1',
		308399 => '1',
		308400 => '1',
		308401 => '1',
		308402 => '1',
		308403 => '1',
		308404 => '1',
		308405 => '1',
		308406 => '1',
		308407 => '1',
		308408 => '1',
		308409 => '1',
		308410 => '1',
		308411 => '1',
		308412 => '1',
		308413 => '1',
		308414 => '1',
		308415 => '1',
		308416 => '1',
		308417 => '1',
		308418 => '1',
		308419 => '1',
		308420 => '1',
		308421 => '1',
		308422 => '1',
		308423 => '1',
		308424 => '1',
		308425 => '1',
		308426 => '1',
		308427 => '1',
		308428 => '1',
		308429 => '1',
		308430 => '1',
		308431 => '1',
		308432 => '1',
		308433 => '1',
		308434 => '1',
		308435 => '1',
		308436 => '1',
		308437 => '1',
		308438 => '1',
		308439 => '1',
		308440 => '1',
		308441 => '1',
		308442 => '1',
		308443 => '1',
		308444 => '1',
		308445 => '1',
		308446 => '1',
		308447 => '1',
		308448 => '1',
		308449 => '1',
		308450 => '1',
		308451 => '1',
		308452 => '1',
		308453 => '1',
		308454 => '1',
		308455 => '1',
		308456 => '1',
		308457 => '1',
		308458 => '1',
		308459 => '1',
		308460 => '1',
		308461 => '1',
		308462 => '1',
		308463 => '1',
		308464 => '1',
		308465 => '1',
		308466 => '1',
		308467 => '1',
		308468 => '1',
		308469 => '1',
		308470 => '1',
		308471 => '1',
		308472 => '1',
		308473 => '1',
		308474 => '1',
		308475 => '1',
		308476 => '1',
		308477 => '1',
		308478 => '1',
		308479 => '1',
		308480 => '1',
		308481 => '1',
		308482 => '1',
		308483 => '1',
		308484 => '1',
		308485 => '1',
		308486 => '1',
		308487 => '1',
		308488 => '1',
		308489 => '1',
		308490 => '1',
		308491 => '1',
		308492 => '1',
		308493 => '1',
		308494 => '1',
		308495 => '1',
		308496 => '1',
		308497 => '1',
		308498 => '1',
		308499 => '1',
		308500 => '1',
		308501 => '1',
		308502 => '1',
		308503 => '1',
		308504 => '1',
		308505 => '1',
		308506 => '1',
		308507 => '1',
		308508 => '1',
		308509 => '1',
		308510 => '1',
		308511 => '1',
		308512 => '1',
		308513 => '1',
		308514 => '1',
		308515 => '1',
		308516 => '1',
		308517 => '1',
		308518 => '1',
		308519 => '1',
		308520 => '1',
		308521 => '1',
		308522 => '1',
		308523 => '1',
		308524 => '1',
		308525 => '1',
		308526 => '1',
		308527 => '1',
		308528 => '1',
		308529 => '1',
		308530 => '1',
		308531 => '1',
		308532 => '1',
		308533 => '1',
		308534 => '1',
		308535 => '1',
		308536 => '1',
		308537 => '1',
		308538 => '1',
		308539 => '1',
		308540 => '1',
		308541 => '1',
		308542 => '1',
		308543 => '1',
		308544 => '1',
		308545 => '1',
		308546 => '1',
		308547 => '1',
		308548 => '1',
		308549 => '1',
		308550 => '1',
		308551 => '1',
		308552 => '1',
		308553 => '1',
		308554 => '1',
		308555 => '1',
		308556 => '1',
		308557 => '1',
		308558 => '1',
		308559 => '1',
		308560 => '1',
		308561 => '1',
		308562 => '1',
		308563 => '1',
		308564 => '1',
		308565 => '1',
		308566 => '1',
		308567 => '1',
		308568 => '1',
		308569 => '1',
		308570 => '1',
		308571 => '1',
		308572 => '1',
		308573 => '1',
		308574 => '1',
		308575 => '1',
		308576 => '1',
		308577 => '1',
		308578 => '1',
		308579 => '1',
		308580 => '1',
		308581 => '1',
		308582 => '1',
		308583 => '1',
		308584 => '1',
		308585 => '1',
		308586 => '1',
		308587 => '1',
		308588 => '1',
		308589 => '1',
		308590 => '1',
		308591 => '1',
		308592 => '1',
		308593 => '1',
		308594 => '1',
		308595 => '1',
		308596 => '1',
		308597 => '1',
		308598 => '1',
		308599 => '1',
		308600 => '1',
		308601 => '1',
		308602 => '1',
		308603 => '1',
		308604 => '1',
		308605 => '1',
		308606 => '1',
		308607 => '1',
		308608 => '1',
		308609 => '1',
		308610 => '1',
		308611 => '1',
		308612 => '1',
		308613 => '1',
		308614 => '1',
		308615 => '1',
		308616 => '1',
		308617 => '1',
		308618 => '1',
		308619 => '1',
		308620 => '1',
		308621 => '1',
		308622 => '1',
		308623 => '1',
		308624 => '1',
		308625 => '1',
		308626 => '1',
		308627 => '1',
		308628 => '1',
		308629 => '1',
		308630 => '1',
		308631 => '1',
		308632 => '1',
		308633 => '1',
		308634 => '1',
		308635 => '1',
		308636 => '1',
		308637 => '1',
		308638 => '1',
		308639 => '1',
		308640 => '1',
		308641 => '1',
		308642 => '1',
		308643 => '1',
		308644 => '1',
		308645 => '1',
		308646 => '1',
		308647 => '1',
		308648 => '1',
		308649 => '1',
		308650 => '1',
		308651 => '1',
		308652 => '1',
		308653 => '1',
		308654 => '1',
		308655 => '1',
		308656 => '1',
		308657 => '1',
		308658 => '1',
		308659 => '1',
		308660 => '1',
		308661 => '1',
		308662 => '1',
		308663 => '1',
		308664 => '1',
		308665 => '1',
		308666 => '1',
		308667 => '1',
		308668 => '1',
		308669 => '1',
		308670 => '1',
		308671 => '1',
		308672 => '1',
		308673 => '1',
		308674 => '1',
		308675 => '1',
		308676 => '1',
		308677 => '1',
		308678 => '1',
		308679 => '1',
		308680 => '1',
		308681 => '1',
		308682 => '1',
		308683 => '1',
		308684 => '1',
		308685 => '1',
		308686 => '1',
		308687 => '1',
		308688 => '1',
		308689 => '1',
		308690 => '1',
		308691 => '1',
		308692 => '1',
		308693 => '1',
		308694 => '1',
		308695 => '1',
		308696 => '1',
		308697 => '1',
		308698 => '1',
		308699 => '1',
		308700 => '1',
		308701 => '1',
		308702 => '1',
		308703 => '1',
		308704 => '1',
		308705 => '1',
		308706 => '1',
		308707 => '1',
		308708 => '1',
		308709 => '1',
		308710 => '1',
		308711 => '1',
		308712 => '1',
		308713 => '1',
		308714 => '1',
		308715 => '1',
		308716 => '1',
		308717 => '1',
		308718 => '1',
		308719 => '1',
		308720 => '1',
		308721 => '1',
		308722 => '1',
		308723 => '1',
		308724 => '1',
		308725 => '1',
		308726 => '1',
		308727 => '1',
		308728 => '1',
		308729 => '1',
		308730 => '1',
		308731 => '1',
		309376 => '1',
		309377 => '1',
		309378 => '1',
		309379 => '1',
		309380 => '1',
		309381 => '1',
		309382 => '1',
		309383 => '1',
		309384 => '1',
		309385 => '1',
		309386 => '1',
		309387 => '1',
		309388 => '1',
		309389 => '1',
		309390 => '1',
		309391 => '1',
		309392 => '1',
		309393 => '1',
		309394 => '1',
		309395 => '1',
		309396 => '1',
		309397 => '1',
		309398 => '1',
		309399 => '1',
		309400 => '1',
		309401 => '1',
		309402 => '1',
		309403 => '1',
		309404 => '1',
		309405 => '1',
		309406 => '1',
		309407 => '1',
		309408 => '1',
		309409 => '1',
		309410 => '1',
		309411 => '1',
		309412 => '1',
		309413 => '1',
		309414 => '1',
		309415 => '1',
		309416 => '1',
		309417 => '1',
		309418 => '1',
		309419 => '1',
		309420 => '1',
		309421 => '1',
		309422 => '1',
		309423 => '1',
		309424 => '1',
		309425 => '1',
		309426 => '1',
		309427 => '1',
		309428 => '1',
		309429 => '1',
		309430 => '1',
		309431 => '1',
		309432 => '1',
		309433 => '1',
		309434 => '1',
		309435 => '1',
		309436 => '1',
		309437 => '1',
		309438 => '1',
		309439 => '1',
		309440 => '1',
		309441 => '1',
		309442 => '1',
		309443 => '1',
		309444 => '1',
		309445 => '1',
		309446 => '1',
		309447 => '1',
		309448 => '1',
		309449 => '1',
		309450 => '1',
		309451 => '1',
		309452 => '1',
		309453 => '1',
		309454 => '1',
		309455 => '1',
		309456 => '1',
		309457 => '1',
		309458 => '1',
		309459 => '1',
		309460 => '1',
		309461 => '1',
		309462 => '1',
		309463 => '1',
		309464 => '1',
		309465 => '1',
		309466 => '1',
		309467 => '1',
		309468 => '1',
		309469 => '1',
		309470 => '1',
		309471 => '1',
		309472 => '1',
		309473 => '1',
		309474 => '1',
		309475 => '1',
		309476 => '1',
		309477 => '1',
		309478 => '1',
		309479 => '1',
		309480 => '1',
		309481 => '1',
		309482 => '1',
		309483 => '1',
		309484 => '1',
		309485 => '1',
		309486 => '1',
		309487 => '1',
		309488 => '1',
		309489 => '1',
		309490 => '1',
		309491 => '1',
		309492 => '1',
		309493 => '1',
		309494 => '1',
		309495 => '1',
		309496 => '1',
		309497 => '1',
		309498 => '1',
		309499 => '1',
		309500 => '1',
		309501 => '1',
		309502 => '1',
		309503 => '1',
		309504 => '1',
		309505 => '1',
		309506 => '1',
		309507 => '1',
		309508 => '1',
		309509 => '1',
		309510 => '1',
		309511 => '1',
		309512 => '1',
		309513 => '1',
		309514 => '1',
		309515 => '1',
		309516 => '1',
		309517 => '1',
		309518 => '1',
		309519 => '1',
		309520 => '1',
		309521 => '1',
		309522 => '1',
		309523 => '1',
		309524 => '1',
		309525 => '1',
		309526 => '1',
		309527 => '1',
		309528 => '1',
		309529 => '1',
		309530 => '1',
		309531 => '1',
		309532 => '1',
		309533 => '1',
		309534 => '1',
		309535 => '1',
		309536 => '1',
		309537 => '1',
		309538 => '1',
		309539 => '1',
		309540 => '1',
		309541 => '1',
		309542 => '1',
		309543 => '1',
		309544 => '1',
		309545 => '1',
		309546 => '1',
		309547 => '1',
		309548 => '1',
		309549 => '1',
		309550 => '1',
		309551 => '1',
		309552 => '1',
		309553 => '1',
		309554 => '1',
		309555 => '1',
		309556 => '1',
		309557 => '1',
		309558 => '1',
		309559 => '1',
		309560 => '1',
		309561 => '1',
		309562 => '1',
		309563 => '1',
		309564 => '1',
		309565 => '1',
		309566 => '1',
		309567 => '1',
		309568 => '1',
		309569 => '1',
		309570 => '1',
		309571 => '1',
		309572 => '1',
		309573 => '1',
		309574 => '1',
		309575 => '1',
		309576 => '1',
		309577 => '1',
		309578 => '1',
		309579 => '1',
		309580 => '1',
		309581 => '1',
		309582 => '1',
		309583 => '1',
		309584 => '1',
		309585 => '1',
		309586 => '1',
		309587 => '1',
		309588 => '1',
		309589 => '1',
		309590 => '1',
		309591 => '1',
		309592 => '1',
		309593 => '1',
		309594 => '1',
		309595 => '1',
		309596 => '1',
		309597 => '1',
		309598 => '1',
		309599 => '1',
		309600 => '1',
		309601 => '1',
		309602 => '1',
		309603 => '1',
		309604 => '1',
		309605 => '1',
		309606 => '1',
		309607 => '1',
		309608 => '1',
		309609 => '1',
		309610 => '1',
		309611 => '1',
		309612 => '1',
		309613 => '1',
		309614 => '1',
		309615 => '1',
		309616 => '1',
		309617 => '1',
		309618 => '1',
		309619 => '1',
		309620 => '1',
		309621 => '1',
		309622 => '1',
		309623 => '1',
		309624 => '1',
		309625 => '1',
		309626 => '1',
		309627 => '1',
		309628 => '1',
		309629 => '1',
		309630 => '1',
		309631 => '1',
		309632 => '1',
		309633 => '1',
		309634 => '1',
		309635 => '1',
		309636 => '1',
		309637 => '1',
		309638 => '1',
		309639 => '1',
		309640 => '1',
		309641 => '1',
		309642 => '1',
		309643 => '1',
		309644 => '1',
		309645 => '1',
		309646 => '1',
		309647 => '1',
		309648 => '1',
		309649 => '1',
		309650 => '1',
		309651 => '1',
		309652 => '1',
		309653 => '1',
		309654 => '1',
		309655 => '1',
		309656 => '1',
		309657 => '1',
		309658 => '1',
		309659 => '1',
		309660 => '1',
		309661 => '1',
		309662 => '1',
		309663 => '1',
		309664 => '1',
		309665 => '1',
		309666 => '1',
		309667 => '1',
		309668 => '1',
		309669 => '1',
		309670 => '1',
		309671 => '1',
		309672 => '1',
		309673 => '1',
		309674 => '1',
		309675 => '1',
		309676 => '1',
		309677 => '1',
		309678 => '1',
		309679 => '1',
		309680 => '1',
		309681 => '1',
		309682 => '1',
		309683 => '1',
		309684 => '1',
		309685 => '1',
		309686 => '1',
		309687 => '1',
		309688 => '1',
		309689 => '1',
		309690 => '1',
		309691 => '1',
		309692 => '1',
		309693 => '1',
		309694 => '1',
		309695 => '1',
		309696 => '1',
		309697 => '1',
		309698 => '1',
		309699 => '1',
		309700 => '1',
		309701 => '1',
		309702 => '1',
		309703 => '1',
		309704 => '1',
		309705 => '1',
		309706 => '1',
		309707 => '1',
		309708 => '1',
		309709 => '1',
		309710 => '1',
		309711 => '1',
		309712 => '1',
		309713 => '1',
		309714 => '1',
		309715 => '1',
		309716 => '1',
		309717 => '1',
		309718 => '1',
		309719 => '1',
		309720 => '1',
		309721 => '1',
		309722 => '1',
		309723 => '1',
		309724 => '1',
		309725 => '1',
		309726 => '1',
		309727 => '1',
		309728 => '1',
		309729 => '1',
		309730 => '1',
		309731 => '1',
		309732 => '1',
		309733 => '1',
		309734 => '1',
		309735 => '1',
		309736 => '1',
		309737 => '1',
		309738 => '1',
		309739 => '1',
		309740 => '1',
		309741 => '1',
		309742 => '1',
		309743 => '1',
		309744 => '1',
		309745 => '1',
		309746 => '1',
		309747 => '1',
		309748 => '1',
		309749 => '1',
		309750 => '1',
		309751 => '1',
		309752 => '1',
		309753 => '1',
		309754 => '1',
		309755 => '1',
		310400 => '1',
		310401 => '1',
		310402 => '1',
		310403 => '1',
		310404 => '1',
		310525 => '1',
		310526 => '1',
		310527 => '1',
		310528 => '1',
		310529 => '1',
		310650 => '1',
		310651 => '1',
		310652 => '1',
		310653 => '1',
		310654 => '1',
		310775 => '1',
		310776 => '1',
		310777 => '1',
		310778 => '1',
		310779 => '1',
		311424 => '1',
		311425 => '1',
		311426 => '1',
		311427 => '1',
		311428 => '1',
		311549 => '1',
		311550 => '1',
		311551 => '1',
		311552 => '1',
		311553 => '1',
		311674 => '1',
		311675 => '1',
		311676 => '1',
		311677 => '1',
		311678 => '1',
		311799 => '1',
		311800 => '1',
		311801 => '1',
		311802 => '1',
		311803 => '1',
		312448 => '1',
		312449 => '1',
		312450 => '1',
		312451 => '1',
		312452 => '1',
		312573 => '1',
		312574 => '1',
		312575 => '1',
		312576 => '1',
		312577 => '1',
		312698 => '1',
		312699 => '1',
		312700 => '1',
		312701 => '1',
		312702 => '1',
		312823 => '1',
		312824 => '1',
		312825 => '1',
		312826 => '1',
		312827 => '1',
		313472 => '1',
		313473 => '1',
		313474 => '1',
		313475 => '1',
		313476 => '1',
		313597 => '1',
		313598 => '1',
		313599 => '1',
		313600 => '1',
		313601 => '1',
		313722 => '1',
		313723 => '1',
		313724 => '1',
		313725 => '1',
		313726 => '1',
		313847 => '1',
		313848 => '1',
		313849 => '1',
		313850 => '1',
		313851 => '1',
		314496 => '1',
		314497 => '1',
		314498 => '1',
		314499 => '1',
		314500 => '1',
		314621 => '1',
		314622 => '1',
		314623 => '1',
		314624 => '1',
		314625 => '1',
		314746 => '1',
		314747 => '1',
		314748 => '1',
		314749 => '1',
		314750 => '1',
		314871 => '1',
		314872 => '1',
		314873 => '1',
		314874 => '1',
		314875 => '1',
		315520 => '1',
		315521 => '1',
		315522 => '1',
		315523 => '1',
		315524 => '1',
		315645 => '1',
		315646 => '1',
		315647 => '1',
		315648 => '1',
		315649 => '1',
		315770 => '1',
		315771 => '1',
		315772 => '1',
		315773 => '1',
		315774 => '1',
		315895 => '1',
		315896 => '1',
		315897 => '1',
		315898 => '1',
		315899 => '1',
		316544 => '1',
		316545 => '1',
		316546 => '1',
		316547 => '1',
		316548 => '1',
		316669 => '1',
		316670 => '1',
		316671 => '1',
		316672 => '1',
		316673 => '1',
		316794 => '1',
		316795 => '1',
		316796 => '1',
		316797 => '1',
		316798 => '1',
		316919 => '1',
		316920 => '1',
		316921 => '1',
		316922 => '1',
		316923 => '1',
		317568 => '1',
		317569 => '1',
		317570 => '1',
		317571 => '1',
		317572 => '1',
		317693 => '1',
		317694 => '1',
		317695 => '1',
		317696 => '1',
		317697 => '1',
		317818 => '1',
		317819 => '1',
		317820 => '1',
		317821 => '1',
		317822 => '1',
		317943 => '1',
		317944 => '1',
		317945 => '1',
		317946 => '1',
		317947 => '1',
		318592 => '1',
		318593 => '1',
		318594 => '1',
		318595 => '1',
		318596 => '1',
		318717 => '1',
		318718 => '1',
		318719 => '1',
		318720 => '1',
		318721 => '1',
		318842 => '1',
		318843 => '1',
		318844 => '1',
		318845 => '1',
		318846 => '1',
		318967 => '1',
		318968 => '1',
		318969 => '1',
		318970 => '1',
		318971 => '1',
		319616 => '1',
		319617 => '1',
		319618 => '1',
		319619 => '1',
		319620 => '1',
		319741 => '1',
		319742 => '1',
		319743 => '1',
		319744 => '1',
		319745 => '1',
		319866 => '1',
		319867 => '1',
		319868 => '1',
		319869 => '1',
		319870 => '1',
		319991 => '1',
		319992 => '1',
		319993 => '1',
		319994 => '1',
		319995 => '1',
		320640 => '1',
		320641 => '1',
		320642 => '1',
		320643 => '1',
		320644 => '1',
		320765 => '1',
		320766 => '1',
		320767 => '1',
		320768 => '1',
		320769 => '1',
		320890 => '1',
		320891 => '1',
		320892 => '1',
		320893 => '1',
		320894 => '1',
		321015 => '1',
		321016 => '1',
		321017 => '1',
		321018 => '1',
		321019 => '1',
		321664 => '1',
		321665 => '1',
		321666 => '1',
		321667 => '1',
		321668 => '1',
		321789 => '1',
		321790 => '1',
		321791 => '1',
		321792 => '1',
		321793 => '1',
		321914 => '1',
		321915 => '1',
		321916 => '1',
		321917 => '1',
		321918 => '1',
		322039 => '1',
		322040 => '1',
		322041 => '1',
		322042 => '1',
		322043 => '1',
		322688 => '1',
		322689 => '1',
		322690 => '1',
		322691 => '1',
		322692 => '1',
		322813 => '1',
		322814 => '1',
		322815 => '1',
		322816 => '1',
		322817 => '1',
		322938 => '1',
		322939 => '1',
		322940 => '1',
		322941 => '1',
		322942 => '1',
		323063 => '1',
		323064 => '1',
		323065 => '1',
		323066 => '1',
		323067 => '1',
		323712 => '1',
		323713 => '1',
		323714 => '1',
		323715 => '1',
		323716 => '1',
		323837 => '1',
		323838 => '1',
		323839 => '1',
		323840 => '1',
		323841 => '1',
		323962 => '1',
		323963 => '1',
		323964 => '1',
		323965 => '1',
		323966 => '1',
		324087 => '1',
		324088 => '1',
		324089 => '1',
		324090 => '1',
		324091 => '1',
		324736 => '1',
		324737 => '1',
		324738 => '1',
		324739 => '1',
		324740 => '1',
		324861 => '1',
		324862 => '1',
		324863 => '1',
		324864 => '1',
		324865 => '1',
		324986 => '1',
		324987 => '1',
		324988 => '1',
		324989 => '1',
		324990 => '1',
		325111 => '1',
		325112 => '1',
		325113 => '1',
		325114 => '1',
		325115 => '1',
		325760 => '1',
		325761 => '1',
		325762 => '1',
		325763 => '1',
		325764 => '1',
		325885 => '1',
		325886 => '1',
		325887 => '1',
		325888 => '1',
		325889 => '1',
		326010 => '1',
		326011 => '1',
		326012 => '1',
		326013 => '1',
		326014 => '1',
		326135 => '1',
		326136 => '1',
		326137 => '1',
		326138 => '1',
		326139 => '1',
		326784 => '1',
		326785 => '1',
		326786 => '1',
		326787 => '1',
		326788 => '1',
		326909 => '1',
		326910 => '1',
		326911 => '1',
		326912 => '1',
		326913 => '1',
		327034 => '1',
		327035 => '1',
		327036 => '1',
		327037 => '1',
		327038 => '1',
		327159 => '1',
		327160 => '1',
		327161 => '1',
		327162 => '1',
		327163 => '1',
		327808 => '1',
		327809 => '1',
		327810 => '1',
		327811 => '1',
		327812 => '1',
		327933 => '1',
		327934 => '1',
		327935 => '1',
		327936 => '1',
		327937 => '1',
		328058 => '1',
		328059 => '1',
		328060 => '1',
		328061 => '1',
		328062 => '1',
		328183 => '1',
		328184 => '1',
		328185 => '1',
		328186 => '1',
		328187 => '1',
		328832 => '1',
		328833 => '1',
		328834 => '1',
		328835 => '1',
		328836 => '1',
		328957 => '1',
		328958 => '1',
		328959 => '1',
		328960 => '1',
		328961 => '1',
		329082 => '1',
		329083 => '1',
		329084 => '1',
		329085 => '1',
		329086 => '1',
		329207 => '1',
		329208 => '1',
		329209 => '1',
		329210 => '1',
		329211 => '1',
		329856 => '1',
		329857 => '1',
		329858 => '1',
		329859 => '1',
		329860 => '1',
		329981 => '1',
		329982 => '1',
		329983 => '1',
		329984 => '1',
		329985 => '1',
		330106 => '1',
		330107 => '1',
		330108 => '1',
		330109 => '1',
		330110 => '1',
		330231 => '1',
		330232 => '1',
		330233 => '1',
		330234 => '1',
		330235 => '1',
		330880 => '1',
		330881 => '1',
		330882 => '1',
		330883 => '1',
		330884 => '1',
		331005 => '1',
		331006 => '1',
		331007 => '1',
		331008 => '1',
		331009 => '1',
		331130 => '1',
		331131 => '1',
		331132 => '1',
		331133 => '1',
		331134 => '1',
		331255 => '1',
		331256 => '1',
		331257 => '1',
		331258 => '1',
		331259 => '1',
		331904 => '1',
		331905 => '1',
		331906 => '1',
		331907 => '1',
		331908 => '1',
		332029 => '1',
		332030 => '1',
		332031 => '1',
		332032 => '1',
		332033 => '1',
		332154 => '1',
		332155 => '1',
		332156 => '1',
		332157 => '1',
		332158 => '1',
		332279 => '1',
		332280 => '1',
		332281 => '1',
		332282 => '1',
		332283 => '1',
		332928 => '1',
		332929 => '1',
		332930 => '1',
		332931 => '1',
		332932 => '1',
		333053 => '1',
		333054 => '1',
		333055 => '1',
		333056 => '1',
		333057 => '1',
		333178 => '1',
		333179 => '1',
		333180 => '1',
		333181 => '1',
		333182 => '1',
		333303 => '1',
		333304 => '1',
		333305 => '1',
		333306 => '1',
		333307 => '1',
		333952 => '1',
		333953 => '1',
		333954 => '1',
		333955 => '1',
		333956 => '1',
		334077 => '1',
		334078 => '1',
		334079 => '1',
		334080 => '1',
		334081 => '1',
		334202 => '1',
		334203 => '1',
		334204 => '1',
		334205 => '1',
		334206 => '1',
		334327 => '1',
		334328 => '1',
		334329 => '1',
		334330 => '1',
		334331 => '1',
		334976 => '1',
		334977 => '1',
		334978 => '1',
		334979 => '1',
		334980 => '1',
		335101 => '1',
		335102 => '1',
		335103 => '1',
		335104 => '1',
		335105 => '1',
		335226 => '1',
		335227 => '1',
		335228 => '1',
		335229 => '1',
		335230 => '1',
		335351 => '1',
		335352 => '1',
		335353 => '1',
		335354 => '1',
		335355 => '1',
		336000 => '1',
		336001 => '1',
		336002 => '1',
		336003 => '1',
		336004 => '1',
		336125 => '1',
		336126 => '1',
		336127 => '1',
		336128 => '1',
		336129 => '1',
		336250 => '1',
		336251 => '1',
		336252 => '1',
		336253 => '1',
		336254 => '1',
		336375 => '1',
		336376 => '1',
		336377 => '1',
		336378 => '1',
		336379 => '1',
		337024 => '1',
		337025 => '1',
		337026 => '1',
		337027 => '1',
		337028 => '1',
		337149 => '1',
		337150 => '1',
		337151 => '1',
		337152 => '1',
		337153 => '1',
		337274 => '1',
		337275 => '1',
		337276 => '1',
		337277 => '1',
		337278 => '1',
		337399 => '1',
		337400 => '1',
		337401 => '1',
		337402 => '1',
		337403 => '1',
		338048 => '1',
		338049 => '1',
		338050 => '1',
		338051 => '1',
		338052 => '1',
		338173 => '1',
		338174 => '1',
		338175 => '1',
		338176 => '1',
		338177 => '1',
		338298 => '1',
		338299 => '1',
		338300 => '1',
		338301 => '1',
		338302 => '1',
		338423 => '1',
		338424 => '1',
		338425 => '1',
		338426 => '1',
		338427 => '1',
		339072 => '1',
		339073 => '1',
		339074 => '1',
		339075 => '1',
		339076 => '1',
		339197 => '1',
		339198 => '1',
		339199 => '1',
		339200 => '1',
		339201 => '1',
		339322 => '1',
		339323 => '1',
		339324 => '1',
		339325 => '1',
		339326 => '1',
		339447 => '1',
		339448 => '1',
		339449 => '1',
		339450 => '1',
		339451 => '1',
		340096 => '1',
		340097 => '1',
		340098 => '1',
		340099 => '1',
		340100 => '1',
		340221 => '1',
		340222 => '1',
		340223 => '1',
		340224 => '1',
		340225 => '1',
		340346 => '1',
		340347 => '1',
		340348 => '1',
		340349 => '1',
		340350 => '1',
		340471 => '1',
		340472 => '1',
		340473 => '1',
		340474 => '1',
		340475 => '1',
		341120 => '1',
		341121 => '1',
		341122 => '1',
		341123 => '1',
		341124 => '1',
		341245 => '1',
		341246 => '1',
		341247 => '1',
		341248 => '1',
		341249 => '1',
		341370 => '1',
		341371 => '1',
		341372 => '1',
		341373 => '1',
		341374 => '1',
		341495 => '1',
		341496 => '1',
		341497 => '1',
		341498 => '1',
		341499 => '1',
		342144 => '1',
		342145 => '1',
		342146 => '1',
		342147 => '1',
		342148 => '1',
		342269 => '1',
		342270 => '1',
		342271 => '1',
		342272 => '1',
		342273 => '1',
		342394 => '1',
		342395 => '1',
		342396 => '1',
		342397 => '1',
		342398 => '1',
		342519 => '1',
		342520 => '1',
		342521 => '1',
		342522 => '1',
		342523 => '1',
		343168 => '1',
		343169 => '1',
		343170 => '1',
		343171 => '1',
		343172 => '1',
		343293 => '1',
		343294 => '1',
		343295 => '1',
		343296 => '1',
		343297 => '1',
		343418 => '1',
		343419 => '1',
		343420 => '1',
		343421 => '1',
		343422 => '1',
		343543 => '1',
		343544 => '1',
		343545 => '1',
		343546 => '1',
		343547 => '1',
		344192 => '1',
		344193 => '1',
		344194 => '1',
		344195 => '1',
		344196 => '1',
		344317 => '1',
		344318 => '1',
		344319 => '1',
		344320 => '1',
		344321 => '1',
		344442 => '1',
		344443 => '1',
		344444 => '1',
		344445 => '1',
		344446 => '1',
		344567 => '1',
		344568 => '1',
		344569 => '1',
		344570 => '1',
		344571 => '1',
		345216 => '1',
		345217 => '1',
		345218 => '1',
		345219 => '1',
		345220 => '1',
		345341 => '1',
		345342 => '1',
		345343 => '1',
		345344 => '1',
		345345 => '1',
		345466 => '1',
		345467 => '1',
		345468 => '1',
		345469 => '1',
		345470 => '1',
		345591 => '1',
		345592 => '1',
		345593 => '1',
		345594 => '1',
		345595 => '1',
		346240 => '1',
		346241 => '1',
		346242 => '1',
		346243 => '1',
		346244 => '1',
		346365 => '1',
		346366 => '1',
		346367 => '1',
		346368 => '1',
		346369 => '1',
		346490 => '1',
		346491 => '1',
		346492 => '1',
		346493 => '1',
		346494 => '1',
		346615 => '1',
		346616 => '1',
		346617 => '1',
		346618 => '1',
		346619 => '1',
		347264 => '1',
		347265 => '1',
		347266 => '1',
		347267 => '1',
		347268 => '1',
		347389 => '1',
		347390 => '1',
		347391 => '1',
		347392 => '1',
		347393 => '1',
		347514 => '1',
		347515 => '1',
		347516 => '1',
		347517 => '1',
		347518 => '1',
		347639 => '1',
		347640 => '1',
		347641 => '1',
		347642 => '1',
		347643 => '1',
		348288 => '1',
		348289 => '1',
		348290 => '1',
		348291 => '1',
		348292 => '1',
		348413 => '1',
		348414 => '1',
		348415 => '1',
		348416 => '1',
		348417 => '1',
		348538 => '1',
		348539 => '1',
		348540 => '1',
		348541 => '1',
		348542 => '1',
		348663 => '1',
		348664 => '1',
		348665 => '1',
		348666 => '1',
		348667 => '1',
		349312 => '1',
		349313 => '1',
		349314 => '1',
		349315 => '1',
		349316 => '1',
		349437 => '1',
		349438 => '1',
		349439 => '1',
		349440 => '1',
		349441 => '1',
		349562 => '1',
		349563 => '1',
		349564 => '1',
		349565 => '1',
		349566 => '1',
		349687 => '1',
		349688 => '1',
		349689 => '1',
		349690 => '1',
		349691 => '1',
		350336 => '1',
		350337 => '1',
		350338 => '1',
		350339 => '1',
		350340 => '1',
		350461 => '1',
		350462 => '1',
		350463 => '1',
		350464 => '1',
		350465 => '1',
		350586 => '1',
		350587 => '1',
		350588 => '1',
		350589 => '1',
		350590 => '1',
		350711 => '1',
		350712 => '1',
		350713 => '1',
		350714 => '1',
		350715 => '1',
		351360 => '1',
		351361 => '1',
		351362 => '1',
		351363 => '1',
		351364 => '1',
		351485 => '1',
		351486 => '1',
		351487 => '1',
		351488 => '1',
		351489 => '1',
		351610 => '1',
		351611 => '1',
		351612 => '1',
		351613 => '1',
		351614 => '1',
		351735 => '1',
		351736 => '1',
		351737 => '1',
		351738 => '1',
		351739 => '1',
		352384 => '1',
		352385 => '1',
		352386 => '1',
		352387 => '1',
		352388 => '1',
		352509 => '1',
		352510 => '1',
		352511 => '1',
		352512 => '1',
		352513 => '1',
		352634 => '1',
		352635 => '1',
		352636 => '1',
		352637 => '1',
		352638 => '1',
		352759 => '1',
		352760 => '1',
		352761 => '1',
		352762 => '1',
		352763 => '1',
		353408 => '1',
		353409 => '1',
		353410 => '1',
		353411 => '1',
		353412 => '1',
		353533 => '1',
		353534 => '1',
		353535 => '1',
		353536 => '1',
		353537 => '1',
		353658 => '1',
		353659 => '1',
		353660 => '1',
		353661 => '1',
		353662 => '1',
		353783 => '1',
		353784 => '1',
		353785 => '1',
		353786 => '1',
		353787 => '1',
		354432 => '1',
		354433 => '1',
		354434 => '1',
		354435 => '1',
		354436 => '1',
		354557 => '1',
		354558 => '1',
		354559 => '1',
		354560 => '1',
		354561 => '1',
		354682 => '1',
		354683 => '1',
		354684 => '1',
		354685 => '1',
		354686 => '1',
		354807 => '1',
		354808 => '1',
		354809 => '1',
		354810 => '1',
		354811 => '1',
		355456 => '1',
		355457 => '1',
		355458 => '1',
		355459 => '1',
		355460 => '1',
		355581 => '1',
		355582 => '1',
		355583 => '1',
		355584 => '1',
		355585 => '1',
		355706 => '1',
		355707 => '1',
		355708 => '1',
		355709 => '1',
		355710 => '1',
		355831 => '1',
		355832 => '1',
		355833 => '1',
		355834 => '1',
		355835 => '1',
		356480 => '1',
		356481 => '1',
		356482 => '1',
		356483 => '1',
		356484 => '1',
		356605 => '1',
		356606 => '1',
		356607 => '1',
		356608 => '1',
		356609 => '1',
		356730 => '1',
		356731 => '1',
		356732 => '1',
		356733 => '1',
		356734 => '1',
		356855 => '1',
		356856 => '1',
		356857 => '1',
		356858 => '1',
		356859 => '1',
		357504 => '1',
		357505 => '1',
		357506 => '1',
		357507 => '1',
		357508 => '1',
		357629 => '1',
		357630 => '1',
		357631 => '1',
		357632 => '1',
		357633 => '1',
		357754 => '1',
		357755 => '1',
		357756 => '1',
		357757 => '1',
		357758 => '1',
		357879 => '1',
		357880 => '1',
		357881 => '1',
		357882 => '1',
		357883 => '1',
		358528 => '1',
		358529 => '1',
		358530 => '1',
		358531 => '1',
		358532 => '1',
		358653 => '1',
		358654 => '1',
		358655 => '1',
		358656 => '1',
		358657 => '1',
		358778 => '1',
		358779 => '1',
		358780 => '1',
		358781 => '1',
		358782 => '1',
		358903 => '1',
		358904 => '1',
		358905 => '1',
		358906 => '1',
		358907 => '1',
		359552 => '1',
		359553 => '1',
		359554 => '1',
		359555 => '1',
		359556 => '1',
		359677 => '1',
		359678 => '1',
		359679 => '1',
		359680 => '1',
		359681 => '1',
		359802 => '1',
		359803 => '1',
		359804 => '1',
		359805 => '1',
		359806 => '1',
		359927 => '1',
		359928 => '1',
		359929 => '1',
		359930 => '1',
		359931 => '1',
		360576 => '1',
		360577 => '1',
		360578 => '1',
		360579 => '1',
		360580 => '1',
		360701 => '1',
		360702 => '1',
		360703 => '1',
		360704 => '1',
		360705 => '1',
		360826 => '1',
		360827 => '1',
		360828 => '1',
		360829 => '1',
		360830 => '1',
		360951 => '1',
		360952 => '1',
		360953 => '1',
		360954 => '1',
		360955 => '1',
		361600 => '1',
		361601 => '1',
		361602 => '1',
		361603 => '1',
		361604 => '1',
		361725 => '1',
		361726 => '1',
		361727 => '1',
		361728 => '1',
		361729 => '1',
		361850 => '1',
		361851 => '1',
		361852 => '1',
		361853 => '1',
		361854 => '1',
		361975 => '1',
		361976 => '1',
		361977 => '1',
		361978 => '1',
		361979 => '1',
		362624 => '1',
		362625 => '1',
		362626 => '1',
		362627 => '1',
		362628 => '1',
		362749 => '1',
		362750 => '1',
		362751 => '1',
		362752 => '1',
		362753 => '1',
		362874 => '1',
		362875 => '1',
		362876 => '1',
		362877 => '1',
		362878 => '1',
		362999 => '1',
		363000 => '1',
		363001 => '1',
		363002 => '1',
		363003 => '1',
		363648 => '1',
		363649 => '1',
		363650 => '1',
		363651 => '1',
		363652 => '1',
		363773 => '1',
		363774 => '1',
		363775 => '1',
		363776 => '1',
		363777 => '1',
		363898 => '1',
		363899 => '1',
		363900 => '1',
		363901 => '1',
		363902 => '1',
		364023 => '1',
		364024 => '1',
		364025 => '1',
		364026 => '1',
		364027 => '1',
		364672 => '1',
		364673 => '1',
		364674 => '1',
		364675 => '1',
		364676 => '1',
		364797 => '1',
		364798 => '1',
		364799 => '1',
		364800 => '1',
		364801 => '1',
		364922 => '1',
		364923 => '1',
		364924 => '1',
		364925 => '1',
		364926 => '1',
		365047 => '1',
		365048 => '1',
		365049 => '1',
		365050 => '1',
		365051 => '1',
		365696 => '1',
		365697 => '1',
		365698 => '1',
		365699 => '1',
		365700 => '1',
		365821 => '1',
		365822 => '1',
		365823 => '1',
		365824 => '1',
		365825 => '1',
		365946 => '1',
		365947 => '1',
		365948 => '1',
		365949 => '1',
		365950 => '1',
		366071 => '1',
		366072 => '1',
		366073 => '1',
		366074 => '1',
		366075 => '1',
		366720 => '1',
		366721 => '1',
		366722 => '1',
		366723 => '1',
		366724 => '1',
		366845 => '1',
		366846 => '1',
		366847 => '1',
		366848 => '1',
		366849 => '1',
		366970 => '1',
		366971 => '1',
		366972 => '1',
		366973 => '1',
		366974 => '1',
		367095 => '1',
		367096 => '1',
		367097 => '1',
		367098 => '1',
		367099 => '1',
		367744 => '1',
		367745 => '1',
		367746 => '1',
		367747 => '1',
		367748 => '1',
		367869 => '1',
		367870 => '1',
		367871 => '1',
		367872 => '1',
		367873 => '1',
		367994 => '1',
		367995 => '1',
		367996 => '1',
		367997 => '1',
		367998 => '1',
		368119 => '1',
		368120 => '1',
		368121 => '1',
		368122 => '1',
		368123 => '1',
		368768 => '1',
		368769 => '1',
		368770 => '1',
		368771 => '1',
		368772 => '1',
		368893 => '1',
		368894 => '1',
		368895 => '1',
		368896 => '1',
		368897 => '1',
		369018 => '1',
		369019 => '1',
		369020 => '1',
		369021 => '1',
		369022 => '1',
		369143 => '1',
		369144 => '1',
		369145 => '1',
		369146 => '1',
		369147 => '1',
		369792 => '1',
		369793 => '1',
		369794 => '1',
		369795 => '1',
		369796 => '1',
		369917 => '1',
		369918 => '1',
		369919 => '1',
		369920 => '1',
		369921 => '1',
		370042 => '1',
		370043 => '1',
		370044 => '1',
		370045 => '1',
		370046 => '1',
		370167 => '1',
		370168 => '1',
		370169 => '1',
		370170 => '1',
		370171 => '1',
		370816 => '1',
		370817 => '1',
		370818 => '1',
		370819 => '1',
		370820 => '1',
		370941 => '1',
		370942 => '1',
		370943 => '1',
		370944 => '1',
		370945 => '1',
		371066 => '1',
		371067 => '1',
		371068 => '1',
		371069 => '1',
		371070 => '1',
		371191 => '1',
		371192 => '1',
		371193 => '1',
		371194 => '1',
		371195 => '1',
		371840 => '1',
		371841 => '1',
		371842 => '1',
		371843 => '1',
		371844 => '1',
		371965 => '1',
		371966 => '1',
		371967 => '1',
		371968 => '1',
		371969 => '1',
		372090 => '1',
		372091 => '1',
		372092 => '1',
		372093 => '1',
		372094 => '1',
		372215 => '1',
		372216 => '1',
		372217 => '1',
		372218 => '1',
		372219 => '1',
		372864 => '1',
		372865 => '1',
		372866 => '1',
		372867 => '1',
		372868 => '1',
		372989 => '1',
		372990 => '1',
		372991 => '1',
		372992 => '1',
		372993 => '1',
		373114 => '1',
		373115 => '1',
		373116 => '1',
		373117 => '1',
		373118 => '1',
		373239 => '1',
		373240 => '1',
		373241 => '1',
		373242 => '1',
		373243 => '1',
		373888 => '1',
		373889 => '1',
		373890 => '1',
		373891 => '1',
		373892 => '1',
		374013 => '1',
		374014 => '1',
		374015 => '1',
		374016 => '1',
		374017 => '1',
		374138 => '1',
		374139 => '1',
		374140 => '1',
		374141 => '1',
		374142 => '1',
		374263 => '1',
		374264 => '1',
		374265 => '1',
		374266 => '1',
		374267 => '1',
		374912 => '1',
		374913 => '1',
		374914 => '1',
		374915 => '1',
		374916 => '1',
		375037 => '1',
		375038 => '1',
		375039 => '1',
		375040 => '1',
		375041 => '1',
		375162 => '1',
		375163 => '1',
		375164 => '1',
		375165 => '1',
		375166 => '1',
		375287 => '1',
		375288 => '1',
		375289 => '1',
		375290 => '1',
		375291 => '1',
		375936 => '1',
		375937 => '1',
		375938 => '1',
		375939 => '1',
		375940 => '1',
		376061 => '1',
		376062 => '1',
		376063 => '1',
		376064 => '1',
		376065 => '1',
		376186 => '1',
		376187 => '1',
		376188 => '1',
		376189 => '1',
		376190 => '1',
		376311 => '1',
		376312 => '1',
		376313 => '1',
		376314 => '1',
		376315 => '1',
		376960 => '1',
		376961 => '1',
		376962 => '1',
		376963 => '1',
		376964 => '1',
		377085 => '1',
		377086 => '1',
		377087 => '1',
		377088 => '1',
		377089 => '1',
		377210 => '1',
		377211 => '1',
		377212 => '1',
		377213 => '1',
		377214 => '1',
		377335 => '1',
		377336 => '1',
		377337 => '1',
		377338 => '1',
		377339 => '1',
		377984 => '1',
		377985 => '1',
		377986 => '1',
		377987 => '1',
		377988 => '1',
		378109 => '1',
		378110 => '1',
		378111 => '1',
		378112 => '1',
		378113 => '1',
		378234 => '1',
		378235 => '1',
		378236 => '1',
		378237 => '1',
		378238 => '1',
		378359 => '1',
		378360 => '1',
		378361 => '1',
		378362 => '1',
		378363 => '1',
		379008 => '1',
		379009 => '1',
		379010 => '1',
		379011 => '1',
		379012 => '1',
		379133 => '1',
		379134 => '1',
		379135 => '1',
		379136 => '1',
		379137 => '1',
		379258 => '1',
		379259 => '1',
		379260 => '1',
		379261 => '1',
		379262 => '1',
		379383 => '1',
		379384 => '1',
		379385 => '1',
		379386 => '1',
		379387 => '1',
		380032 => '1',
		380033 => '1',
		380034 => '1',
		380035 => '1',
		380036 => '1',
		380157 => '1',
		380158 => '1',
		380159 => '1',
		380160 => '1',
		380161 => '1',
		380282 => '1',
		380283 => '1',
		380284 => '1',
		380285 => '1',
		380286 => '1',
		380407 => '1',
		380408 => '1',
		380409 => '1',
		380410 => '1',
		380411 => '1',
		381056 => '1',
		381057 => '1',
		381058 => '1',
		381059 => '1',
		381060 => '1',
		381181 => '1',
		381182 => '1',
		381183 => '1',
		381184 => '1',
		381185 => '1',
		381306 => '1',
		381307 => '1',
		381308 => '1',
		381309 => '1',
		381310 => '1',
		381431 => '1',
		381432 => '1',
		381433 => '1',
		381434 => '1',
		381435 => '1',
		382080 => '1',
		382081 => '1',
		382082 => '1',
		382083 => '1',
		382084 => '1',
		382205 => '1',
		382206 => '1',
		382207 => '1',
		382208 => '1',
		382209 => '1',
		382330 => '1',
		382331 => '1',
		382332 => '1',
		382333 => '1',
		382334 => '1',
		382455 => '1',
		382456 => '1',
		382457 => '1',
		382458 => '1',
		382459 => '1',
		383104 => '1',
		383105 => '1',
		383106 => '1',
		383107 => '1',
		383108 => '1',
		383229 => '1',
		383230 => '1',
		383231 => '1',
		383232 => '1',
		383233 => '1',
		383354 => '1',
		383355 => '1',
		383356 => '1',
		383357 => '1',
		383358 => '1',
		383479 => '1',
		383480 => '1',
		383481 => '1',
		383482 => '1',
		383483 => '1',
		384128 => '1',
		384129 => '1',
		384130 => '1',
		384131 => '1',
		384132 => '1',
		384253 => '1',
		384254 => '1',
		384255 => '1',
		384256 => '1',
		384257 => '1',
		384378 => '1',
		384379 => '1',
		384380 => '1',
		384381 => '1',
		384382 => '1',
		384503 => '1',
		384504 => '1',
		384505 => '1',
		384506 => '1',
		384507 => '1',
		385152 => '1',
		385153 => '1',
		385154 => '1',
		385155 => '1',
		385156 => '1',
		385277 => '1',
		385278 => '1',
		385279 => '1',
		385280 => '1',
		385281 => '1',
		385402 => '1',
		385403 => '1',
		385404 => '1',
		385405 => '1',
		385406 => '1',
		385527 => '1',
		385528 => '1',
		385529 => '1',
		385530 => '1',
		385531 => '1',
		386176 => '1',
		386177 => '1',
		386178 => '1',
		386179 => '1',
		386180 => '1',
		386301 => '1',
		386302 => '1',
		386303 => '1',
		386304 => '1',
		386305 => '1',
		386426 => '1',
		386427 => '1',
		386428 => '1',
		386429 => '1',
		386430 => '1',
		386551 => '1',
		386552 => '1',
		386553 => '1',
		386554 => '1',
		386555 => '1',
		387200 => '1',
		387201 => '1',
		387202 => '1',
		387203 => '1',
		387204 => '1',
		387325 => '1',
		387326 => '1',
		387327 => '1',
		387328 => '1',
		387329 => '1',
		387450 => '1',
		387451 => '1',
		387452 => '1',
		387453 => '1',
		387454 => '1',
		387575 => '1',
		387576 => '1',
		387577 => '1',
		387578 => '1',
		387579 => '1',
		388224 => '1',
		388225 => '1',
		388226 => '1',
		388227 => '1',
		388228 => '1',
		388349 => '1',
		388350 => '1',
		388351 => '1',
		388352 => '1',
		388353 => '1',
		388474 => '1',
		388475 => '1',
		388476 => '1',
		388477 => '1',
		388478 => '1',
		388599 => '1',
		388600 => '1',
		388601 => '1',
		388602 => '1',
		388603 => '1',
		389248 => '1',
		389249 => '1',
		389250 => '1',
		389251 => '1',
		389252 => '1',
		389373 => '1',
		389374 => '1',
		389375 => '1',
		389376 => '1',
		389377 => '1',
		389498 => '1',
		389499 => '1',
		389500 => '1',
		389501 => '1',
		389502 => '1',
		389623 => '1',
		389624 => '1',
		389625 => '1',
		389626 => '1',
		389627 => '1',
		390272 => '1',
		390273 => '1',
		390274 => '1',
		390275 => '1',
		390276 => '1',
		390397 => '1',
		390398 => '1',
		390399 => '1',
		390400 => '1',
		390401 => '1',
		390522 => '1',
		390523 => '1',
		390524 => '1',
		390525 => '1',
		390526 => '1',
		390647 => '1',
		390648 => '1',
		390649 => '1',
		390650 => '1',
		390651 => '1',
		391296 => '1',
		391297 => '1',
		391298 => '1',
		391299 => '1',
		391300 => '1',
		391421 => '1',
		391422 => '1',
		391423 => '1',
		391424 => '1',
		391425 => '1',
		391546 => '1',
		391547 => '1',
		391548 => '1',
		391549 => '1',
		391550 => '1',
		391671 => '1',
		391672 => '1',
		391673 => '1',
		391674 => '1',
		391675 => '1',
		392320 => '1',
		392321 => '1',
		392322 => '1',
		392323 => '1',
		392324 => '1',
		392445 => '1',
		392446 => '1',
		392447 => '1',
		392448 => '1',
		392449 => '1',
		392570 => '1',
		392571 => '1',
		392572 => '1',
		392573 => '1',
		392574 => '1',
		392695 => '1',
		392696 => '1',
		392697 => '1',
		392698 => '1',
		392699 => '1',
		393344 => '1',
		393345 => '1',
		393346 => '1',
		393347 => '1',
		393348 => '1',
		393469 => '1',
		393470 => '1',
		393471 => '1',
		393472 => '1',
		393473 => '1',
		393594 => '1',
		393595 => '1',
		393596 => '1',
		393597 => '1',
		393598 => '1',
		393719 => '1',
		393720 => '1',
		393721 => '1',
		393722 => '1',
		393723 => '1',
		394368 => '1',
		394369 => '1',
		394370 => '1',
		394371 => '1',
		394372 => '1',
		394493 => '1',
		394494 => '1',
		394495 => '1',
		394496 => '1',
		394497 => '1',
		394618 => '1',
		394619 => '1',
		394620 => '1',
		394621 => '1',
		394622 => '1',
		394743 => '1',
		394744 => '1',
		394745 => '1',
		394746 => '1',
		394747 => '1',
		395392 => '1',
		395393 => '1',
		395394 => '1',
		395395 => '1',
		395396 => '1',
		395517 => '1',
		395518 => '1',
		395519 => '1',
		395520 => '1',
		395521 => '1',
		395642 => '1',
		395643 => '1',
		395644 => '1',
		395645 => '1',
		395646 => '1',
		395767 => '1',
		395768 => '1',
		395769 => '1',
		395770 => '1',
		395771 => '1',
		396416 => '1',
		396417 => '1',
		396418 => '1',
		396419 => '1',
		396420 => '1',
		396541 => '1',
		396542 => '1',
		396543 => '1',
		396544 => '1',
		396545 => '1',
		396666 => '1',
		396667 => '1',
		396668 => '1',
		396669 => '1',
		396670 => '1',
		396791 => '1',
		396792 => '1',
		396793 => '1',
		396794 => '1',
		396795 => '1',
		397440 => '1',
		397441 => '1',
		397442 => '1',
		397443 => '1',
		397444 => '1',
		397565 => '1',
		397566 => '1',
		397567 => '1',
		397568 => '1',
		397569 => '1',
		397690 => '1',
		397691 => '1',
		397692 => '1',
		397693 => '1',
		397694 => '1',
		397815 => '1',
		397816 => '1',
		397817 => '1',
		397818 => '1',
		397819 => '1',
		398464 => '1',
		398465 => '1',
		398466 => '1',
		398467 => '1',
		398468 => '1',
		398589 => '1',
		398590 => '1',
		398591 => '1',
		398592 => '1',
		398593 => '1',
		398714 => '1',
		398715 => '1',
		398716 => '1',
		398717 => '1',
		398718 => '1',
		398839 => '1',
		398840 => '1',
		398841 => '1',
		398842 => '1',
		398843 => '1',
		399488 => '1',
		399489 => '1',
		399490 => '1',
		399491 => '1',
		399492 => '1',
		399613 => '1',
		399614 => '1',
		399615 => '1',
		399616 => '1',
		399617 => '1',
		399738 => '1',
		399739 => '1',
		399740 => '1',
		399741 => '1',
		399742 => '1',
		399863 => '1',
		399864 => '1',
		399865 => '1',
		399866 => '1',
		399867 => '1',
		400512 => '1',
		400513 => '1',
		400514 => '1',
		400515 => '1',
		400516 => '1',
		400637 => '1',
		400638 => '1',
		400639 => '1',
		400640 => '1',
		400641 => '1',
		400762 => '1',
		400763 => '1',
		400764 => '1',
		400765 => '1',
		400766 => '1',
		400887 => '1',
		400888 => '1',
		400889 => '1',
		400890 => '1',
		400891 => '1',
		401536 => '1',
		401537 => '1',
		401538 => '1',
		401539 => '1',
		401540 => '1',
		401661 => '1',
		401662 => '1',
		401663 => '1',
		401664 => '1',
		401665 => '1',
		401786 => '1',
		401787 => '1',
		401788 => '1',
		401789 => '1',
		401790 => '1',
		401911 => '1',
		401912 => '1',
		401913 => '1',
		401914 => '1',
		401915 => '1',
		402560 => '1',
		402561 => '1',
		402562 => '1',
		402563 => '1',
		402564 => '1',
		402685 => '1',
		402686 => '1',
		402687 => '1',
		402688 => '1',
		402689 => '1',
		402810 => '1',
		402811 => '1',
		402812 => '1',
		402813 => '1',
		402814 => '1',
		402935 => '1',
		402936 => '1',
		402937 => '1',
		402938 => '1',
		402939 => '1',
		403584 => '1',
		403585 => '1',
		403586 => '1',
		403587 => '1',
		403588 => '1',
		403709 => '1',
		403710 => '1',
		403711 => '1',
		403712 => '1',
		403713 => '1',
		403834 => '1',
		403835 => '1',
		403836 => '1',
		403837 => '1',
		403838 => '1',
		403959 => '1',
		403960 => '1',
		403961 => '1',
		403962 => '1',
		403963 => '1',
		404608 => '1',
		404609 => '1',
		404610 => '1',
		404611 => '1',
		404612 => '1',
		404733 => '1',
		404734 => '1',
		404735 => '1',
		404736 => '1',
		404737 => '1',
		404858 => '1',
		404859 => '1',
		404860 => '1',
		404861 => '1',
		404862 => '1',
		404983 => '1',
		404984 => '1',
		404985 => '1',
		404986 => '1',
		404987 => '1',
		405632 => '1',
		405633 => '1',
		405634 => '1',
		405635 => '1',
		405636 => '1',
		405757 => '1',
		405758 => '1',
		405759 => '1',
		405760 => '1',
		405761 => '1',
		405882 => '1',
		405883 => '1',
		405884 => '1',
		405885 => '1',
		405886 => '1',
		406007 => '1',
		406008 => '1',
		406009 => '1',
		406010 => '1',
		406011 => '1',
		406656 => '1',
		406657 => '1',
		406658 => '1',
		406659 => '1',
		406660 => '1',
		406781 => '1',
		406782 => '1',
		406783 => '1',
		406784 => '1',
		406785 => '1',
		406906 => '1',
		406907 => '1',
		406908 => '1',
		406909 => '1',
		406910 => '1',
		407031 => '1',
		407032 => '1',
		407033 => '1',
		407034 => '1',
		407035 => '1',
		407680 => '1',
		407681 => '1',
		407682 => '1',
		407683 => '1',
		407684 => '1',
		407805 => '1',
		407806 => '1',
		407807 => '1',
		407808 => '1',
		407809 => '1',
		407930 => '1',
		407931 => '1',
		407932 => '1',
		407933 => '1',
		407934 => '1',
		408055 => '1',
		408056 => '1',
		408057 => '1',
		408058 => '1',
		408059 => '1',
		408704 => '1',
		408705 => '1',
		408706 => '1',
		408707 => '1',
		408708 => '1',
		408829 => '1',
		408830 => '1',
		408831 => '1',
		408832 => '1',
		408833 => '1',
		408954 => '1',
		408955 => '1',
		408956 => '1',
		408957 => '1',
		408958 => '1',
		409079 => '1',
		409080 => '1',
		409081 => '1',
		409082 => '1',
		409083 => '1',
		409728 => '1',
		409729 => '1',
		409730 => '1',
		409731 => '1',
		409732 => '1',
		409853 => '1',
		409854 => '1',
		409855 => '1',
		409856 => '1',
		409857 => '1',
		409978 => '1',
		409979 => '1',
		409980 => '1',
		409981 => '1',
		409982 => '1',
		410103 => '1',
		410104 => '1',
		410105 => '1',
		410106 => '1',
		410107 => '1',
		410752 => '1',
		410753 => '1',
		410754 => '1',
		410755 => '1',
		410756 => '1',
		410877 => '1',
		410878 => '1',
		410879 => '1',
		410880 => '1',
		410881 => '1',
		411002 => '1',
		411003 => '1',
		411004 => '1',
		411005 => '1',
		411006 => '1',
		411127 => '1',
		411128 => '1',
		411129 => '1',
		411130 => '1',
		411131 => '1',
		411776 => '1',
		411777 => '1',
		411778 => '1',
		411779 => '1',
		411780 => '1',
		411901 => '1',
		411902 => '1',
		411903 => '1',
		411904 => '1',
		411905 => '1',
		412026 => '1',
		412027 => '1',
		412028 => '1',
		412029 => '1',
		412030 => '1',
		412151 => '1',
		412152 => '1',
		412153 => '1',
		412154 => '1',
		412155 => '1',
		412800 => '1',
		412801 => '1',
		412802 => '1',
		412803 => '1',
		412804 => '1',
		412925 => '1',
		412926 => '1',
		412927 => '1',
		412928 => '1',
		412929 => '1',
		413050 => '1',
		413051 => '1',
		413052 => '1',
		413053 => '1',
		413054 => '1',
		413175 => '1',
		413176 => '1',
		413177 => '1',
		413178 => '1',
		413179 => '1',
		413824 => '1',
		413825 => '1',
		413826 => '1',
		413827 => '1',
		413828 => '1',
		413949 => '1',
		413950 => '1',
		413951 => '1',
		413952 => '1',
		413953 => '1',
		414074 => '1',
		414075 => '1',
		414076 => '1',
		414077 => '1',
		414078 => '1',
		414199 => '1',
		414200 => '1',
		414201 => '1',
		414202 => '1',
		414203 => '1',
		414848 => '1',
		414849 => '1',
		414850 => '1',
		414851 => '1',
		414852 => '1',
		414973 => '1',
		414974 => '1',
		414975 => '1',
		414976 => '1',
		414977 => '1',
		415098 => '1',
		415099 => '1',
		415100 => '1',
		415101 => '1',
		415102 => '1',
		415223 => '1',
		415224 => '1',
		415225 => '1',
		415226 => '1',
		415227 => '1',
		415872 => '1',
		415873 => '1',
		415874 => '1',
		415875 => '1',
		415876 => '1',
		415997 => '1',
		415998 => '1',
		415999 => '1',
		416000 => '1',
		416001 => '1',
		416122 => '1',
		416123 => '1',
		416124 => '1',
		416125 => '1',
		416126 => '1',
		416247 => '1',
		416248 => '1',
		416249 => '1',
		416250 => '1',
		416251 => '1',
		416896 => '1',
		416897 => '1',
		416898 => '1',
		416899 => '1',
		416900 => '1',
		417021 => '1',
		417022 => '1',
		417023 => '1',
		417024 => '1',
		417025 => '1',
		417146 => '1',
		417147 => '1',
		417148 => '1',
		417149 => '1',
		417150 => '1',
		417271 => '1',
		417272 => '1',
		417273 => '1',
		417274 => '1',
		417275 => '1',
		417920 => '1',
		417921 => '1',
		417922 => '1',
		417923 => '1',
		417924 => '1',
		418045 => '1',
		418046 => '1',
		418047 => '1',
		418048 => '1',
		418049 => '1',
		418170 => '1',
		418171 => '1',
		418172 => '1',
		418173 => '1',
		418174 => '1',
		418295 => '1',
		418296 => '1',
		418297 => '1',
		418298 => '1',
		418299 => '1',
		418944 => '1',
		418945 => '1',
		418946 => '1',
		418947 => '1',
		418948 => '1',
		419069 => '1',
		419070 => '1',
		419071 => '1',
		419072 => '1',
		419073 => '1',
		419194 => '1',
		419195 => '1',
		419196 => '1',
		419197 => '1',
		419198 => '1',
		419319 => '1',
		419320 => '1',
		419321 => '1',
		419322 => '1',
		419323 => '1',
		419968 => '1',
		419969 => '1',
		419970 => '1',
		419971 => '1',
		419972 => '1',
		420093 => '1',
		420094 => '1',
		420095 => '1',
		420096 => '1',
		420097 => '1',
		420218 => '1',
		420219 => '1',
		420220 => '1',
		420221 => '1',
		420222 => '1',
		420343 => '1',
		420344 => '1',
		420345 => '1',
		420346 => '1',
		420347 => '1',
		420992 => '1',
		420993 => '1',
		420994 => '1',
		420995 => '1',
		420996 => '1',
		421117 => '1',
		421118 => '1',
		421119 => '1',
		421120 => '1',
		421121 => '1',
		421242 => '1',
		421243 => '1',
		421244 => '1',
		421245 => '1',
		421246 => '1',
		421367 => '1',
		421368 => '1',
		421369 => '1',
		421370 => '1',
		421371 => '1',
		422016 => '1',
		422017 => '1',
		422018 => '1',
		422019 => '1',
		422020 => '1',
		422141 => '1',
		422142 => '1',
		422143 => '1',
		422144 => '1',
		422145 => '1',
		422266 => '1',
		422267 => '1',
		422268 => '1',
		422269 => '1',
		422270 => '1',
		422391 => '1',
		422392 => '1',
		422393 => '1',
		422394 => '1',
		422395 => '1',
		423040 => '1',
		423041 => '1',
		423042 => '1',
		423043 => '1',
		423044 => '1',
		423165 => '1',
		423166 => '1',
		423167 => '1',
		423168 => '1',
		423169 => '1',
		423290 => '1',
		423291 => '1',
		423292 => '1',
		423293 => '1',
		423294 => '1',
		423415 => '1',
		423416 => '1',
		423417 => '1',
		423418 => '1',
		423419 => '1',
		424064 => '1',
		424065 => '1',
		424066 => '1',
		424067 => '1',
		424068 => '1',
		424189 => '1',
		424190 => '1',
		424191 => '1',
		424192 => '1',
		424193 => '1',
		424314 => '1',
		424315 => '1',
		424316 => '1',
		424317 => '1',
		424318 => '1',
		424439 => '1',
		424440 => '1',
		424441 => '1',
		424442 => '1',
		424443 => '1',
		425088 => '1',
		425089 => '1',
		425090 => '1',
		425091 => '1',
		425092 => '1',
		425213 => '1',
		425214 => '1',
		425215 => '1',
		425216 => '1',
		425217 => '1',
		425338 => '1',
		425339 => '1',
		425340 => '1',
		425341 => '1',
		425342 => '1',
		425463 => '1',
		425464 => '1',
		425465 => '1',
		425466 => '1',
		425467 => '1',
		426112 => '1',
		426113 => '1',
		426114 => '1',
		426115 => '1',
		426116 => '1',
		426237 => '1',
		426238 => '1',
		426239 => '1',
		426240 => '1',
		426241 => '1',
		426362 => '1',
		426363 => '1',
		426364 => '1',
		426365 => '1',
		426366 => '1',
		426487 => '1',
		426488 => '1',
		426489 => '1',
		426490 => '1',
		426491 => '1',
		427136 => '1',
		427137 => '1',
		427138 => '1',
		427139 => '1',
		427140 => '1',
		427261 => '1',
		427262 => '1',
		427263 => '1',
		427264 => '1',
		427265 => '1',
		427386 => '1',
		427387 => '1',
		427388 => '1',
		427389 => '1',
		427390 => '1',
		427511 => '1',
		427512 => '1',
		427513 => '1',
		427514 => '1',
		427515 => '1',
		428160 => '1',
		428161 => '1',
		428162 => '1',
		428163 => '1',
		428164 => '1',
		428285 => '1',
		428286 => '1',
		428287 => '1',
		428288 => '1',
		428289 => '1',
		428410 => '1',
		428411 => '1',
		428412 => '1',
		428413 => '1',
		428414 => '1',
		428535 => '1',
		428536 => '1',
		428537 => '1',
		428538 => '1',
		428539 => '1',
		429184 => '1',
		429185 => '1',
		429186 => '1',
		429187 => '1',
		429188 => '1',
		429309 => '1',
		429310 => '1',
		429311 => '1',
		429312 => '1',
		429313 => '1',
		429434 => '1',
		429435 => '1',
		429436 => '1',
		429437 => '1',
		429438 => '1',
		429559 => '1',
		429560 => '1',
		429561 => '1',
		429562 => '1',
		429563 => '1',
		430208 => '1',
		430209 => '1',
		430210 => '1',
		430211 => '1',
		430212 => '1',
		430333 => '1',
		430334 => '1',
		430335 => '1',
		430336 => '1',
		430337 => '1',
		430458 => '1',
		430459 => '1',
		430460 => '1',
		430461 => '1',
		430462 => '1',
		430583 => '1',
		430584 => '1',
		430585 => '1',
		430586 => '1',
		430587 => '1',
		431232 => '1',
		431233 => '1',
		431234 => '1',
		431235 => '1',
		431236 => '1',
		431357 => '1',
		431358 => '1',
		431359 => '1',
		431360 => '1',
		431361 => '1',
		431482 => '1',
		431483 => '1',
		431484 => '1',
		431485 => '1',
		431486 => '1',
		431607 => '1',
		431608 => '1',
		431609 => '1',
		431610 => '1',
		431611 => '1',
		432256 => '1',
		432257 => '1',
		432258 => '1',
		432259 => '1',
		432260 => '1',
		432381 => '1',
		432382 => '1',
		432383 => '1',
		432384 => '1',
		432385 => '1',
		432506 => '1',
		432507 => '1',
		432508 => '1',
		432509 => '1',
		432510 => '1',
		432631 => '1',
		432632 => '1',
		432633 => '1',
		432634 => '1',
		432635 => '1',
		433280 => '1',
		433281 => '1',
		433282 => '1',
		433283 => '1',
		433284 => '1',
		433285 => '1',
		433286 => '1',
		433287 => '1',
		433288 => '1',
		433289 => '1',
		433290 => '1',
		433291 => '1',
		433292 => '1',
		433293 => '1',
		433294 => '1',
		433295 => '1',
		433296 => '1',
		433297 => '1',
		433298 => '1',
		433299 => '1',
		433300 => '1',
		433301 => '1',
		433302 => '1',
		433303 => '1',
		433304 => '1',
		433305 => '1',
		433306 => '1',
		433307 => '1',
		433308 => '1',
		433309 => '1',
		433310 => '1',
		433311 => '1',
		433312 => '1',
		433313 => '1',
		433314 => '1',
		433315 => '1',
		433316 => '1',
		433317 => '1',
		433318 => '1',
		433319 => '1',
		433320 => '1',
		433321 => '1',
		433322 => '1',
		433323 => '1',
		433324 => '1',
		433325 => '1',
		433326 => '1',
		433327 => '1',
		433328 => '1',
		433329 => '1',
		433330 => '1',
		433331 => '1',
		433332 => '1',
		433333 => '1',
		433334 => '1',
		433335 => '1',
		433336 => '1',
		433337 => '1',
		433338 => '1',
		433339 => '1',
		433340 => '1',
		433341 => '1',
		433342 => '1',
		433343 => '1',
		433344 => '1',
		433345 => '1',
		433346 => '1',
		433347 => '1',
		433348 => '1',
		433349 => '1',
		433350 => '1',
		433351 => '1',
		433352 => '1',
		433353 => '1',
		433354 => '1',
		433355 => '1',
		433356 => '1',
		433357 => '1',
		433358 => '1',
		433359 => '1',
		433360 => '1',
		433361 => '1',
		433362 => '1',
		433363 => '1',
		433364 => '1',
		433365 => '1',
		433366 => '1',
		433367 => '1',
		433368 => '1',
		433369 => '1',
		433370 => '1',
		433371 => '1',
		433372 => '1',
		433373 => '1',
		433374 => '1',
		433375 => '1',
		433376 => '1',
		433377 => '1',
		433378 => '1',
		433379 => '1',
		433380 => '1',
		433381 => '1',
		433382 => '1',
		433383 => '1',
		433384 => '1',
		433385 => '1',
		433386 => '1',
		433387 => '1',
		433388 => '1',
		433389 => '1',
		433390 => '1',
		433391 => '1',
		433392 => '1',
		433393 => '1',
		433394 => '1',
		433395 => '1',
		433396 => '1',
		433397 => '1',
		433398 => '1',
		433399 => '1',
		433400 => '1',
		433401 => '1',
		433402 => '1',
		433403 => '1',
		433404 => '1',
		433405 => '1',
		433406 => '1',
		433407 => '1',
		433408 => '1',
		433409 => '1',
		433410 => '1',
		433411 => '1',
		433412 => '1',
		433413 => '1',
		433414 => '1',
		433415 => '1',
		433416 => '1',
		433417 => '1',
		433418 => '1',
		433419 => '1',
		433420 => '1',
		433421 => '1',
		433422 => '1',
		433423 => '1',
		433424 => '1',
		433425 => '1',
		433426 => '1',
		433427 => '1',
		433428 => '1',
		433429 => '1',
		433430 => '1',
		433431 => '1',
		433432 => '1',
		433433 => '1',
		433434 => '1',
		433435 => '1',
		433436 => '1',
		433437 => '1',
		433438 => '1',
		433439 => '1',
		433440 => '1',
		433441 => '1',
		433442 => '1',
		433443 => '1',
		433444 => '1',
		433445 => '1',
		433446 => '1',
		433447 => '1',
		433448 => '1',
		433449 => '1',
		433450 => '1',
		433451 => '1',
		433452 => '1',
		433453 => '1',
		433454 => '1',
		433455 => '1',
		433456 => '1',
		433457 => '1',
		433458 => '1',
		433459 => '1',
		433460 => '1',
		433461 => '1',
		433462 => '1',
		433463 => '1',
		433464 => '1',
		433465 => '1',
		433466 => '1',
		433467 => '1',
		433468 => '1',
		433469 => '1',
		433470 => '1',
		433471 => '1',
		433472 => '1',
		433473 => '1',
		433474 => '1',
		433475 => '1',
		433476 => '1',
		433477 => '1',
		433478 => '1',
		433479 => '1',
		433480 => '1',
		433481 => '1',
		433482 => '1',
		433483 => '1',
		433484 => '1',
		433485 => '1',
		433486 => '1',
		433487 => '1',
		433488 => '1',
		433489 => '1',
		433490 => '1',
		433491 => '1',
		433492 => '1',
		433493 => '1',
		433494 => '1',
		433495 => '1',
		433496 => '1',
		433497 => '1',
		433498 => '1',
		433499 => '1',
		433500 => '1',
		433501 => '1',
		433502 => '1',
		433503 => '1',
		433504 => '1',
		433505 => '1',
		433506 => '1',
		433507 => '1',
		433508 => '1',
		433509 => '1',
		433510 => '1',
		433511 => '1',
		433512 => '1',
		433513 => '1',
		433514 => '1',
		433515 => '1',
		433516 => '1',
		433517 => '1',
		433518 => '1',
		433519 => '1',
		433520 => '1',
		433521 => '1',
		433522 => '1',
		433523 => '1',
		433524 => '1',
		433525 => '1',
		433526 => '1',
		433527 => '1',
		433528 => '1',
		433529 => '1',
		433530 => '1',
		433531 => '1',
		433532 => '1',
		433533 => '1',
		433534 => '1',
		433535 => '1',
		433536 => '1',
		433537 => '1',
		433538 => '1',
		433539 => '1',
		433540 => '1',
		433541 => '1',
		433542 => '1',
		433543 => '1',
		433544 => '1',
		433545 => '1',
		433546 => '1',
		433547 => '1',
		433548 => '1',
		433549 => '1',
		433550 => '1',
		433551 => '1',
		433552 => '1',
		433553 => '1',
		433554 => '1',
		433555 => '1',
		433556 => '1',
		433557 => '1',
		433558 => '1',
		433559 => '1',
		433560 => '1',
		433561 => '1',
		433562 => '1',
		433563 => '1',
		433564 => '1',
		433565 => '1',
		433566 => '1',
		433567 => '1',
		433568 => '1',
		433569 => '1',
		433570 => '1',
		433571 => '1',
		433572 => '1',
		433573 => '1',
		433574 => '1',
		433575 => '1',
		433576 => '1',
		433577 => '1',
		433578 => '1',
		433579 => '1',
		433580 => '1',
		433581 => '1',
		433582 => '1',
		433583 => '1',
		433584 => '1',
		433585 => '1',
		433586 => '1',
		433587 => '1',
		433588 => '1',
		433589 => '1',
		433590 => '1',
		433591 => '1',
		433592 => '1',
		433593 => '1',
		433594 => '1',
		433595 => '1',
		433596 => '1',
		433597 => '1',
		433598 => '1',
		433599 => '1',
		433600 => '1',
		433601 => '1',
		433602 => '1',
		433603 => '1',
		433604 => '1',
		433605 => '1',
		433606 => '1',
		433607 => '1',
		433608 => '1',
		433609 => '1',
		433610 => '1',
		433611 => '1',
		433612 => '1',
		433613 => '1',
		433614 => '1',
		433615 => '1',
		433616 => '1',
		433617 => '1',
		433618 => '1',
		433619 => '1',
		433620 => '1',
		433621 => '1',
		433622 => '1',
		433623 => '1',
		433624 => '1',
		433625 => '1',
		433626 => '1',
		433627 => '1',
		433628 => '1',
		433629 => '1',
		433630 => '1',
		433631 => '1',
		433632 => '1',
		433633 => '1',
		433634 => '1',
		433635 => '1',
		433636 => '1',
		433637 => '1',
		433638 => '1',
		433639 => '1',
		433640 => '1',
		433641 => '1',
		433642 => '1',
		433643 => '1',
		433644 => '1',
		433645 => '1',
		433646 => '1',
		433647 => '1',
		433648 => '1',
		433649 => '1',
		433650 => '1',
		433651 => '1',
		433652 => '1',
		433653 => '1',
		433654 => '1',
		433655 => '1',
		433656 => '1',
		433657 => '1',
		433658 => '1',
		433659 => '1',
		434304 => '1',
		434305 => '1',
		434306 => '1',
		434307 => '1',
		434308 => '1',
		434309 => '1',
		434310 => '1',
		434311 => '1',
		434312 => '1',
		434313 => '1',
		434314 => '1',
		434315 => '1',
		434316 => '1',
		434317 => '1',
		434318 => '1',
		434319 => '1',
		434320 => '1',
		434321 => '1',
		434322 => '1',
		434323 => '1',
		434324 => '1',
		434325 => '1',
		434326 => '1',
		434327 => '1',
		434328 => '1',
		434329 => '1',
		434330 => '1',
		434331 => '1',
		434332 => '1',
		434333 => '1',
		434334 => '1',
		434335 => '1',
		434336 => '1',
		434337 => '1',
		434338 => '1',
		434339 => '1',
		434340 => '1',
		434341 => '1',
		434342 => '1',
		434343 => '1',
		434344 => '1',
		434345 => '1',
		434346 => '1',
		434347 => '1',
		434348 => '1',
		434349 => '1',
		434350 => '1',
		434351 => '1',
		434352 => '1',
		434353 => '1',
		434354 => '1',
		434355 => '1',
		434356 => '1',
		434357 => '1',
		434358 => '1',
		434359 => '1',
		434360 => '1',
		434361 => '1',
		434362 => '1',
		434363 => '1',
		434364 => '1',
		434365 => '1',
		434366 => '1',
		434367 => '1',
		434368 => '1',
		434369 => '1',
		434370 => '1',
		434371 => '1',
		434372 => '1',
		434373 => '1',
		434374 => '1',
		434375 => '1',
		434376 => '1',
		434377 => '1',
		434378 => '1',
		434379 => '1',
		434380 => '1',
		434381 => '1',
		434382 => '1',
		434383 => '1',
		434384 => '1',
		434385 => '1',
		434386 => '1',
		434387 => '1',
		434388 => '1',
		434389 => '1',
		434390 => '1',
		434391 => '1',
		434392 => '1',
		434393 => '1',
		434394 => '1',
		434395 => '1',
		434396 => '1',
		434397 => '1',
		434398 => '1',
		434399 => '1',
		434400 => '1',
		434401 => '1',
		434402 => '1',
		434403 => '1',
		434404 => '1',
		434405 => '1',
		434406 => '1',
		434407 => '1',
		434408 => '1',
		434409 => '1',
		434410 => '1',
		434411 => '1',
		434412 => '1',
		434413 => '1',
		434414 => '1',
		434415 => '1',
		434416 => '1',
		434417 => '1',
		434418 => '1',
		434419 => '1',
		434420 => '1',
		434421 => '1',
		434422 => '1',
		434423 => '1',
		434424 => '1',
		434425 => '1',
		434426 => '1',
		434427 => '1',
		434428 => '1',
		434429 => '1',
		434430 => '1',
		434431 => '1',
		434432 => '1',
		434433 => '1',
		434434 => '1',
		434435 => '1',
		434436 => '1',
		434437 => '1',
		434438 => '1',
		434439 => '1',
		434440 => '1',
		434441 => '1',
		434442 => '1',
		434443 => '1',
		434444 => '1',
		434445 => '1',
		434446 => '1',
		434447 => '1',
		434448 => '1',
		434449 => '1',
		434450 => '1',
		434451 => '1',
		434452 => '1',
		434453 => '1',
		434454 => '1',
		434455 => '1',
		434456 => '1',
		434457 => '1',
		434458 => '1',
		434459 => '1',
		434460 => '1',
		434461 => '1',
		434462 => '1',
		434463 => '1',
		434464 => '1',
		434465 => '1',
		434466 => '1',
		434467 => '1',
		434468 => '1',
		434469 => '1',
		434470 => '1',
		434471 => '1',
		434472 => '1',
		434473 => '1',
		434474 => '1',
		434475 => '1',
		434476 => '1',
		434477 => '1',
		434478 => '1',
		434479 => '1',
		434480 => '1',
		434481 => '1',
		434482 => '1',
		434483 => '1',
		434484 => '1',
		434485 => '1',
		434486 => '1',
		434487 => '1',
		434488 => '1',
		434489 => '1',
		434490 => '1',
		434491 => '1',
		434492 => '1',
		434493 => '1',
		434494 => '1',
		434495 => '1',
		434496 => '1',
		434497 => '1',
		434498 => '1',
		434499 => '1',
		434500 => '1',
		434501 => '1',
		434502 => '1',
		434503 => '1',
		434504 => '1',
		434505 => '1',
		434506 => '1',
		434507 => '1',
		434508 => '1',
		434509 => '1',
		434510 => '1',
		434511 => '1',
		434512 => '1',
		434513 => '1',
		434514 => '1',
		434515 => '1',
		434516 => '1',
		434517 => '1',
		434518 => '1',
		434519 => '1',
		434520 => '1',
		434521 => '1',
		434522 => '1',
		434523 => '1',
		434524 => '1',
		434525 => '1',
		434526 => '1',
		434527 => '1',
		434528 => '1',
		434529 => '1',
		434530 => '1',
		434531 => '1',
		434532 => '1',
		434533 => '1',
		434534 => '1',
		434535 => '1',
		434536 => '1',
		434537 => '1',
		434538 => '1',
		434539 => '1',
		434540 => '1',
		434541 => '1',
		434542 => '1',
		434543 => '1',
		434544 => '1',
		434545 => '1',
		434546 => '1',
		434547 => '1',
		434548 => '1',
		434549 => '1',
		434550 => '1',
		434551 => '1',
		434552 => '1',
		434553 => '1',
		434554 => '1',
		434555 => '1',
		434556 => '1',
		434557 => '1',
		434558 => '1',
		434559 => '1',
		434560 => '1',
		434561 => '1',
		434562 => '1',
		434563 => '1',
		434564 => '1',
		434565 => '1',
		434566 => '1',
		434567 => '1',
		434568 => '1',
		434569 => '1',
		434570 => '1',
		434571 => '1',
		434572 => '1',
		434573 => '1',
		434574 => '1',
		434575 => '1',
		434576 => '1',
		434577 => '1',
		434578 => '1',
		434579 => '1',
		434580 => '1',
		434581 => '1',
		434582 => '1',
		434583 => '1',
		434584 => '1',
		434585 => '1',
		434586 => '1',
		434587 => '1',
		434588 => '1',
		434589 => '1',
		434590 => '1',
		434591 => '1',
		434592 => '1',
		434593 => '1',
		434594 => '1',
		434595 => '1',
		434596 => '1',
		434597 => '1',
		434598 => '1',
		434599 => '1',
		434600 => '1',
		434601 => '1',
		434602 => '1',
		434603 => '1',
		434604 => '1',
		434605 => '1',
		434606 => '1',
		434607 => '1',
		434608 => '1',
		434609 => '1',
		434610 => '1',
		434611 => '1',
		434612 => '1',
		434613 => '1',
		434614 => '1',
		434615 => '1',
		434616 => '1',
		434617 => '1',
		434618 => '1',
		434619 => '1',
		434620 => '1',
		434621 => '1',
		434622 => '1',
		434623 => '1',
		434624 => '1',
		434625 => '1',
		434626 => '1',
		434627 => '1',
		434628 => '1',
		434629 => '1',
		434630 => '1',
		434631 => '1',
		434632 => '1',
		434633 => '1',
		434634 => '1',
		434635 => '1',
		434636 => '1',
		434637 => '1',
		434638 => '1',
		434639 => '1',
		434640 => '1',
		434641 => '1',
		434642 => '1',
		434643 => '1',
		434644 => '1',
		434645 => '1',
		434646 => '1',
		434647 => '1',
		434648 => '1',
		434649 => '1',
		434650 => '1',
		434651 => '1',
		434652 => '1',
		434653 => '1',
		434654 => '1',
		434655 => '1',
		434656 => '1',
		434657 => '1',
		434658 => '1',
		434659 => '1',
		434660 => '1',
		434661 => '1',
		434662 => '1',
		434663 => '1',
		434664 => '1',
		434665 => '1',
		434666 => '1',
		434667 => '1',
		434668 => '1',
		434669 => '1',
		434670 => '1',
		434671 => '1',
		434672 => '1',
		434673 => '1',
		434674 => '1',
		434675 => '1',
		434676 => '1',
		434677 => '1',
		434678 => '1',
		434679 => '1',
		434680 => '1',
		434681 => '1',
		434682 => '1',
		434683 => '1',
		435328 => '1',
		435329 => '1',
		435330 => '1',
		435331 => '1',
		435332 => '1',
		435333 => '1',
		435334 => '1',
		435335 => '1',
		435336 => '1',
		435337 => '1',
		435338 => '1',
		435339 => '1',
		435340 => '1',
		435341 => '1',
		435342 => '1',
		435343 => '1',
		435344 => '1',
		435345 => '1',
		435346 => '1',
		435347 => '1',
		435348 => '1',
		435349 => '1',
		435350 => '1',
		435351 => '1',
		435352 => '1',
		435353 => '1',
		435354 => '1',
		435355 => '1',
		435356 => '1',
		435357 => '1',
		435358 => '1',
		435359 => '1',
		435360 => '1',
		435361 => '1',
		435362 => '1',
		435363 => '1',
		435364 => '1',
		435365 => '1',
		435366 => '1',
		435367 => '1',
		435368 => '1',
		435369 => '1',
		435370 => '1',
		435371 => '1',
		435372 => '1',
		435373 => '1',
		435374 => '1',
		435375 => '1',
		435376 => '1',
		435377 => '1',
		435378 => '1',
		435379 => '1',
		435380 => '1',
		435381 => '1',
		435382 => '1',
		435383 => '1',
		435384 => '1',
		435385 => '1',
		435386 => '1',
		435387 => '1',
		435388 => '1',
		435389 => '1',
		435390 => '1',
		435391 => '1',
		435392 => '1',
		435393 => '1',
		435394 => '1',
		435395 => '1',
		435396 => '1',
		435397 => '1',
		435398 => '1',
		435399 => '1',
		435400 => '1',
		435401 => '1',
		435402 => '1',
		435403 => '1',
		435404 => '1',
		435405 => '1',
		435406 => '1',
		435407 => '1',
		435408 => '1',
		435409 => '1',
		435410 => '1',
		435411 => '1',
		435412 => '1',
		435413 => '1',
		435414 => '1',
		435415 => '1',
		435416 => '1',
		435417 => '1',
		435418 => '1',
		435419 => '1',
		435420 => '1',
		435421 => '1',
		435422 => '1',
		435423 => '1',
		435424 => '1',
		435425 => '1',
		435426 => '1',
		435427 => '1',
		435428 => '1',
		435429 => '1',
		435430 => '1',
		435431 => '1',
		435432 => '1',
		435433 => '1',
		435434 => '1',
		435435 => '1',
		435436 => '1',
		435437 => '1',
		435438 => '1',
		435439 => '1',
		435440 => '1',
		435441 => '1',
		435442 => '1',
		435443 => '1',
		435444 => '1',
		435445 => '1',
		435446 => '1',
		435447 => '1',
		435448 => '1',
		435449 => '1',
		435450 => '1',
		435451 => '1',
		435452 => '1',
		435453 => '1',
		435454 => '1',
		435455 => '1',
		435456 => '1',
		435457 => '1',
		435458 => '1',
		435459 => '1',
		435460 => '1',
		435461 => '1',
		435462 => '1',
		435463 => '1',
		435464 => '1',
		435465 => '1',
		435466 => '1',
		435467 => '1',
		435468 => '1',
		435469 => '1',
		435470 => '1',
		435471 => '1',
		435472 => '1',
		435473 => '1',
		435474 => '1',
		435475 => '1',
		435476 => '1',
		435477 => '1',
		435478 => '1',
		435479 => '1',
		435480 => '1',
		435481 => '1',
		435482 => '1',
		435483 => '1',
		435484 => '1',
		435485 => '1',
		435486 => '1',
		435487 => '1',
		435488 => '1',
		435489 => '1',
		435490 => '1',
		435491 => '1',
		435492 => '1',
		435493 => '1',
		435494 => '1',
		435495 => '1',
		435496 => '1',
		435497 => '1',
		435498 => '1',
		435499 => '1',
		435500 => '1',
		435501 => '1',
		435502 => '1',
		435503 => '1',
		435504 => '1',
		435505 => '1',
		435506 => '1',
		435507 => '1',
		435508 => '1',
		435509 => '1',
		435510 => '1',
		435511 => '1',
		435512 => '1',
		435513 => '1',
		435514 => '1',
		435515 => '1',
		435516 => '1',
		435517 => '1',
		435518 => '1',
		435519 => '1',
		435520 => '1',
		435521 => '1',
		435522 => '1',
		435523 => '1',
		435524 => '1',
		435525 => '1',
		435526 => '1',
		435527 => '1',
		435528 => '1',
		435529 => '1',
		435530 => '1',
		435531 => '1',
		435532 => '1',
		435533 => '1',
		435534 => '1',
		435535 => '1',
		435536 => '1',
		435537 => '1',
		435538 => '1',
		435539 => '1',
		435540 => '1',
		435541 => '1',
		435542 => '1',
		435543 => '1',
		435544 => '1',
		435545 => '1',
		435546 => '1',
		435547 => '1',
		435548 => '1',
		435549 => '1',
		435550 => '1',
		435551 => '1',
		435552 => '1',
		435553 => '1',
		435554 => '1',
		435555 => '1',
		435556 => '1',
		435557 => '1',
		435558 => '1',
		435559 => '1',
		435560 => '1',
		435561 => '1',
		435562 => '1',
		435563 => '1',
		435564 => '1',
		435565 => '1',
		435566 => '1',
		435567 => '1',
		435568 => '1',
		435569 => '1',
		435570 => '1',
		435571 => '1',
		435572 => '1',
		435573 => '1',
		435574 => '1',
		435575 => '1',
		435576 => '1',
		435577 => '1',
		435578 => '1',
		435579 => '1',
		435580 => '1',
		435581 => '1',
		435582 => '1',
		435583 => '1',
		435584 => '1',
		435585 => '1',
		435586 => '1',
		435587 => '1',
		435588 => '1',
		435589 => '1',
		435590 => '1',
		435591 => '1',
		435592 => '1',
		435593 => '1',
		435594 => '1',
		435595 => '1',
		435596 => '1',
		435597 => '1',
		435598 => '1',
		435599 => '1',
		435600 => '1',
		435601 => '1',
		435602 => '1',
		435603 => '1',
		435604 => '1',
		435605 => '1',
		435606 => '1',
		435607 => '1',
		435608 => '1',
		435609 => '1',
		435610 => '1',
		435611 => '1',
		435612 => '1',
		435613 => '1',
		435614 => '1',
		435615 => '1',
		435616 => '1',
		435617 => '1',
		435618 => '1',
		435619 => '1',
		435620 => '1',
		435621 => '1',
		435622 => '1',
		435623 => '1',
		435624 => '1',
		435625 => '1',
		435626 => '1',
		435627 => '1',
		435628 => '1',
		435629 => '1',
		435630 => '1',
		435631 => '1',
		435632 => '1',
		435633 => '1',
		435634 => '1',
		435635 => '1',
		435636 => '1',
		435637 => '1',
		435638 => '1',
		435639 => '1',
		435640 => '1',
		435641 => '1',
		435642 => '1',
		435643 => '1',
		435644 => '1',
		435645 => '1',
		435646 => '1',
		435647 => '1',
		435648 => '1',
		435649 => '1',
		435650 => '1',
		435651 => '1',
		435652 => '1',
		435653 => '1',
		435654 => '1',
		435655 => '1',
		435656 => '1',
		435657 => '1',
		435658 => '1',
		435659 => '1',
		435660 => '1',
		435661 => '1',
		435662 => '1',
		435663 => '1',
		435664 => '1',
		435665 => '1',
		435666 => '1',
		435667 => '1',
		435668 => '1',
		435669 => '1',
		435670 => '1',
		435671 => '1',
		435672 => '1',
		435673 => '1',
		435674 => '1',
		435675 => '1',
		435676 => '1',
		435677 => '1',
		435678 => '1',
		435679 => '1',
		435680 => '1',
		435681 => '1',
		435682 => '1',
		435683 => '1',
		435684 => '1',
		435685 => '1',
		435686 => '1',
		435687 => '1',
		435688 => '1',
		435689 => '1',
		435690 => '1',
		435691 => '1',
		435692 => '1',
		435693 => '1',
		435694 => '1',
		435695 => '1',
		435696 => '1',
		435697 => '1',
		435698 => '1',
		435699 => '1',
		435700 => '1',
		435701 => '1',
		435702 => '1',
		435703 => '1',
		435704 => '1',
		435705 => '1',
		435706 => '1',
		435707 => '1',
		436352 => '1',
		436353 => '1',
		436354 => '1',
		436355 => '1',
		436356 => '1',
		436357 => '1',
		436358 => '1',
		436359 => '1',
		436360 => '1',
		436361 => '1',
		436362 => '1',
		436363 => '1',
		436364 => '1',
		436365 => '1',
		436366 => '1',
		436367 => '1',
		436368 => '1',
		436369 => '1',
		436370 => '1',
		436371 => '1',
		436372 => '1',
		436373 => '1',
		436374 => '1',
		436375 => '1',
		436376 => '1',
		436377 => '1',
		436378 => '1',
		436379 => '1',
		436380 => '1',
		436381 => '1',
		436382 => '1',
		436383 => '1',
		436384 => '1',
		436385 => '1',
		436386 => '1',
		436387 => '1',
		436388 => '1',
		436389 => '1',
		436390 => '1',
		436391 => '1',
		436392 => '1',
		436393 => '1',
		436394 => '1',
		436395 => '1',
		436396 => '1',
		436397 => '1',
		436398 => '1',
		436399 => '1',
		436400 => '1',
		436401 => '1',
		436402 => '1',
		436403 => '1',
		436404 => '1',
		436405 => '1',
		436406 => '1',
		436407 => '1',
		436408 => '1',
		436409 => '1',
		436410 => '1',
		436411 => '1',
		436412 => '1',
		436413 => '1',
		436414 => '1',
		436415 => '1',
		436416 => '1',
		436417 => '1',
		436418 => '1',
		436419 => '1',
		436420 => '1',
		436421 => '1',
		436422 => '1',
		436423 => '1',
		436424 => '1',
		436425 => '1',
		436426 => '1',
		436427 => '1',
		436428 => '1',
		436429 => '1',
		436430 => '1',
		436431 => '1',
		436432 => '1',
		436433 => '1',
		436434 => '1',
		436435 => '1',
		436436 => '1',
		436437 => '1',
		436438 => '1',
		436439 => '1',
		436440 => '1',
		436441 => '1',
		436442 => '1',
		436443 => '1',
		436444 => '1',
		436445 => '1',
		436446 => '1',
		436447 => '1',
		436448 => '1',
		436449 => '1',
		436450 => '1',
		436451 => '1',
		436452 => '1',
		436453 => '1',
		436454 => '1',
		436455 => '1',
		436456 => '1',
		436457 => '1',
		436458 => '1',
		436459 => '1',
		436460 => '1',
		436461 => '1',
		436462 => '1',
		436463 => '1',
		436464 => '1',
		436465 => '1',
		436466 => '1',
		436467 => '1',
		436468 => '1',
		436469 => '1',
		436470 => '1',
		436471 => '1',
		436472 => '1',
		436473 => '1',
		436474 => '1',
		436475 => '1',
		436476 => '1',
		436477 => '1',
		436478 => '1',
		436479 => '1',
		436480 => '1',
		436481 => '1',
		436482 => '1',
		436483 => '1',
		436484 => '1',
		436485 => '1',
		436486 => '1',
		436487 => '1',
		436488 => '1',
		436489 => '1',
		436490 => '1',
		436491 => '1',
		436492 => '1',
		436493 => '1',
		436494 => '1',
		436495 => '1',
		436496 => '1',
		436497 => '1',
		436498 => '1',
		436499 => '1',
		436500 => '1',
		436501 => '1',
		436502 => '1',
		436503 => '1',
		436504 => '1',
		436505 => '1',
		436506 => '1',
		436507 => '1',
		436508 => '1',
		436509 => '1',
		436510 => '1',
		436511 => '1',
		436512 => '1',
		436513 => '1',
		436514 => '1',
		436515 => '1',
		436516 => '1',
		436517 => '1',
		436518 => '1',
		436519 => '1',
		436520 => '1',
		436521 => '1',
		436522 => '1',
		436523 => '1',
		436524 => '1',
		436525 => '1',
		436526 => '1',
		436527 => '1',
		436528 => '1',
		436529 => '1',
		436530 => '1',
		436531 => '1',
		436532 => '1',
		436533 => '1',
		436534 => '1',
		436535 => '1',
		436536 => '1',
		436537 => '1',
		436538 => '1',
		436539 => '1',
		436540 => '1',
		436541 => '1',
		436542 => '1',
		436543 => '1',
		436544 => '1',
		436545 => '1',
		436546 => '1',
		436547 => '1',
		436548 => '1',
		436549 => '1',
		436550 => '1',
		436551 => '1',
		436552 => '1',
		436553 => '1',
		436554 => '1',
		436555 => '1',
		436556 => '1',
		436557 => '1',
		436558 => '1',
		436559 => '1',
		436560 => '1',
		436561 => '1',
		436562 => '1',
		436563 => '1',
		436564 => '1',
		436565 => '1',
		436566 => '1',
		436567 => '1',
		436568 => '1',
		436569 => '1',
		436570 => '1',
		436571 => '1',
		436572 => '1',
		436573 => '1',
		436574 => '1',
		436575 => '1',
		436576 => '1',
		436577 => '1',
		436578 => '1',
		436579 => '1',
		436580 => '1',
		436581 => '1',
		436582 => '1',
		436583 => '1',
		436584 => '1',
		436585 => '1',
		436586 => '1',
		436587 => '1',
		436588 => '1',
		436589 => '1',
		436590 => '1',
		436591 => '1',
		436592 => '1',
		436593 => '1',
		436594 => '1',
		436595 => '1',
		436596 => '1',
		436597 => '1',
		436598 => '1',
		436599 => '1',
		436600 => '1',
		436601 => '1',
		436602 => '1',
		436603 => '1',
		436604 => '1',
		436605 => '1',
		436606 => '1',
		436607 => '1',
		436608 => '1',
		436609 => '1',
		436610 => '1',
		436611 => '1',
		436612 => '1',
		436613 => '1',
		436614 => '1',
		436615 => '1',
		436616 => '1',
		436617 => '1',
		436618 => '1',
		436619 => '1',
		436620 => '1',
		436621 => '1',
		436622 => '1',
		436623 => '1',
		436624 => '1',
		436625 => '1',
		436626 => '1',
		436627 => '1',
		436628 => '1',
		436629 => '1',
		436630 => '1',
		436631 => '1',
		436632 => '1',
		436633 => '1',
		436634 => '1',
		436635 => '1',
		436636 => '1',
		436637 => '1',
		436638 => '1',
		436639 => '1',
		436640 => '1',
		436641 => '1',
		436642 => '1',
		436643 => '1',
		436644 => '1',
		436645 => '1',
		436646 => '1',
		436647 => '1',
		436648 => '1',
		436649 => '1',
		436650 => '1',
		436651 => '1',
		436652 => '1',
		436653 => '1',
		436654 => '1',
		436655 => '1',
		436656 => '1',
		436657 => '1',
		436658 => '1',
		436659 => '1',
		436660 => '1',
		436661 => '1',
		436662 => '1',
		436663 => '1',
		436664 => '1',
		436665 => '1',
		436666 => '1',
		436667 => '1',
		436668 => '1',
		436669 => '1',
		436670 => '1',
		436671 => '1',
		436672 => '1',
		436673 => '1',
		436674 => '1',
		436675 => '1',
		436676 => '1',
		436677 => '1',
		436678 => '1',
		436679 => '1',
		436680 => '1',
		436681 => '1',
		436682 => '1',
		436683 => '1',
		436684 => '1',
		436685 => '1',
		436686 => '1',
		436687 => '1',
		436688 => '1',
		436689 => '1',
		436690 => '1',
		436691 => '1',
		436692 => '1',
		436693 => '1',
		436694 => '1',
		436695 => '1',
		436696 => '1',
		436697 => '1',
		436698 => '1',
		436699 => '1',
		436700 => '1',
		436701 => '1',
		436702 => '1',
		436703 => '1',
		436704 => '1',
		436705 => '1',
		436706 => '1',
		436707 => '1',
		436708 => '1',
		436709 => '1',
		436710 => '1',
		436711 => '1',
		436712 => '1',
		436713 => '1',
		436714 => '1',
		436715 => '1',
		436716 => '1',
		436717 => '1',
		436718 => '1',
		436719 => '1',
		436720 => '1',
		436721 => '1',
		436722 => '1',
		436723 => '1',
		436724 => '1',
		436725 => '1',
		436726 => '1',
		436727 => '1',
		436728 => '1',
		436729 => '1',
		436730 => '1',
		436731 => '1',
		437376 => '1',
		437377 => '1',
		437378 => '1',
		437379 => '1',
		437380 => '1',
		437381 => '1',
		437382 => '1',
		437383 => '1',
		437384 => '1',
		437385 => '1',
		437386 => '1',
		437387 => '1',
		437388 => '1',
		437389 => '1',
		437390 => '1',
		437391 => '1',
		437392 => '1',
		437393 => '1',
		437394 => '1',
		437395 => '1',
		437396 => '1',
		437397 => '1',
		437398 => '1',
		437399 => '1',
		437400 => '1',
		437401 => '1',
		437402 => '1',
		437403 => '1',
		437404 => '1',
		437405 => '1',
		437406 => '1',
		437407 => '1',
		437408 => '1',
		437409 => '1',
		437410 => '1',
		437411 => '1',
		437412 => '1',
		437413 => '1',
		437414 => '1',
		437415 => '1',
		437416 => '1',
		437417 => '1',
		437418 => '1',
		437419 => '1',
		437420 => '1',
		437421 => '1',
		437422 => '1',
		437423 => '1',
		437424 => '1',
		437425 => '1',
		437426 => '1',
		437427 => '1',
		437428 => '1',
		437429 => '1',
		437430 => '1',
		437431 => '1',
		437432 => '1',
		437433 => '1',
		437434 => '1',
		437435 => '1',
		437436 => '1',
		437437 => '1',
		437438 => '1',
		437439 => '1',
		437440 => '1',
		437441 => '1',
		437442 => '1',
		437443 => '1',
		437444 => '1',
		437445 => '1',
		437446 => '1',
		437447 => '1',
		437448 => '1',
		437449 => '1',
		437450 => '1',
		437451 => '1',
		437452 => '1',
		437453 => '1',
		437454 => '1',
		437455 => '1',
		437456 => '1',
		437457 => '1',
		437458 => '1',
		437459 => '1',
		437460 => '1',
		437461 => '1',
		437462 => '1',
		437463 => '1',
		437464 => '1',
		437465 => '1',
		437466 => '1',
		437467 => '1',
		437468 => '1',
		437469 => '1',
		437470 => '1',
		437471 => '1',
		437472 => '1',
		437473 => '1',
		437474 => '1',
		437475 => '1',
		437476 => '1',
		437477 => '1',
		437478 => '1',
		437479 => '1',
		437480 => '1',
		437481 => '1',
		437482 => '1',
		437483 => '1',
		437484 => '1',
		437485 => '1',
		437486 => '1',
		437487 => '1',
		437488 => '1',
		437489 => '1',
		437490 => '1',
		437491 => '1',
		437492 => '1',
		437493 => '1',
		437494 => '1',
		437495 => '1',
		437496 => '1',
		437497 => '1',
		437498 => '1',
		437499 => '1',
		437500 => '1',
		437501 => '1',
		437502 => '1',
		437503 => '1',
		437504 => '1',
		437505 => '1',
		437506 => '1',
		437507 => '1',
		437508 => '1',
		437509 => '1',
		437510 => '1',
		437511 => '1',
		437512 => '1',
		437513 => '1',
		437514 => '1',
		437515 => '1',
		437516 => '1',
		437517 => '1',
		437518 => '1',
		437519 => '1',
		437520 => '1',
		437521 => '1',
		437522 => '1',
		437523 => '1',
		437524 => '1',
		437525 => '1',
		437526 => '1',
		437527 => '1',
		437528 => '1',
		437529 => '1',
		437530 => '1',
		437531 => '1',
		437532 => '1',
		437533 => '1',
		437534 => '1',
		437535 => '1',
		437536 => '1',
		437537 => '1',
		437538 => '1',
		437539 => '1',
		437540 => '1',
		437541 => '1',
		437542 => '1',
		437543 => '1',
		437544 => '1',
		437545 => '1',
		437546 => '1',
		437547 => '1',
		437548 => '1',
		437549 => '1',
		437550 => '1',
		437551 => '1',
		437552 => '1',
		437553 => '1',
		437554 => '1',
		437555 => '1',
		437556 => '1',
		437557 => '1',
		437558 => '1',
		437559 => '1',
		437560 => '1',
		437561 => '1',
		437562 => '1',
		437563 => '1',
		437564 => '1',
		437565 => '1',
		437566 => '1',
		437567 => '1',
		437568 => '1',
		437569 => '1',
		437570 => '1',
		437571 => '1',
		437572 => '1',
		437573 => '1',
		437574 => '1',
		437575 => '1',
		437576 => '1',
		437577 => '1',
		437578 => '1',
		437579 => '1',
		437580 => '1',
		437581 => '1',
		437582 => '1',
		437583 => '1',
		437584 => '1',
		437585 => '1',
		437586 => '1',
		437587 => '1',
		437588 => '1',
		437589 => '1',
		437590 => '1',
		437591 => '1',
		437592 => '1',
		437593 => '1',
		437594 => '1',
		437595 => '1',
		437596 => '1',
		437597 => '1',
		437598 => '1',
		437599 => '1',
		437600 => '1',
		437601 => '1',
		437602 => '1',
		437603 => '1',
		437604 => '1',
		437605 => '1',
		437606 => '1',
		437607 => '1',
		437608 => '1',
		437609 => '1',
		437610 => '1',
		437611 => '1',
		437612 => '1',
		437613 => '1',
		437614 => '1',
		437615 => '1',
		437616 => '1',
		437617 => '1',
		437618 => '1',
		437619 => '1',
		437620 => '1',
		437621 => '1',
		437622 => '1',
		437623 => '1',
		437624 => '1',
		437625 => '1',
		437626 => '1',
		437627 => '1',
		437628 => '1',
		437629 => '1',
		437630 => '1',
		437631 => '1',
		437632 => '1',
		437633 => '1',
		437634 => '1',
		437635 => '1',
		437636 => '1',
		437637 => '1',
		437638 => '1',
		437639 => '1',
		437640 => '1',
		437641 => '1',
		437642 => '1',
		437643 => '1',
		437644 => '1',
		437645 => '1',
		437646 => '1',
		437647 => '1',
		437648 => '1',
		437649 => '1',
		437650 => '1',
		437651 => '1',
		437652 => '1',
		437653 => '1',
		437654 => '1',
		437655 => '1',
		437656 => '1',
		437657 => '1',
		437658 => '1',
		437659 => '1',
		437660 => '1',
		437661 => '1',
		437662 => '1',
		437663 => '1',
		437664 => '1',
		437665 => '1',
		437666 => '1',
		437667 => '1',
		437668 => '1',
		437669 => '1',
		437670 => '1',
		437671 => '1',
		437672 => '1',
		437673 => '1',
		437674 => '1',
		437675 => '1',
		437676 => '1',
		437677 => '1',
		437678 => '1',
		437679 => '1',
		437680 => '1',
		437681 => '1',
		437682 => '1',
		437683 => '1',
		437684 => '1',
		437685 => '1',
		437686 => '1',
		437687 => '1',
		437688 => '1',
		437689 => '1',
		437690 => '1',
		437691 => '1',
		437692 => '1',
		437693 => '1',
		437694 => '1',
		437695 => '1',
		437696 => '1',
		437697 => '1',
		437698 => '1',
		437699 => '1',
		437700 => '1',
		437701 => '1',
		437702 => '1',
		437703 => '1',
		437704 => '1',
		437705 => '1',
		437706 => '1',
		437707 => '1',
		437708 => '1',
		437709 => '1',
		437710 => '1',
		437711 => '1',
		437712 => '1',
		437713 => '1',
		437714 => '1',
		437715 => '1',
		437716 => '1',
		437717 => '1',
		437718 => '1',
		437719 => '1',
		437720 => '1',
		437721 => '1',
		437722 => '1',
		437723 => '1',
		437724 => '1',
		437725 => '1',
		437726 => '1',
		437727 => '1',
		437728 => '1',
		437729 => '1',
		437730 => '1',
		437731 => '1',
		437732 => '1',
		437733 => '1',
		437734 => '1',
		437735 => '1',
		437736 => '1',
		437737 => '1',
		437738 => '1',
		437739 => '1',
		437740 => '1',
		437741 => '1',
		437742 => '1',
		437743 => '1',
		437744 => '1',
		437745 => '1',
		437746 => '1',
		437747 => '1',
		437748 => '1',
		437749 => '1',
		437750 => '1',
		437751 => '1',
		437752 => '1',
		437753 => '1',
		437754 => '1',
		437755 => '1',
