library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM_vide_sel is
	port (CLK : in std_logic;
		  EN : in std_logic;
		  ADDR : in std_logic_vector(11 downto 0);
		  DATA : out std_logic_vector(7 downto 0));
end ROM_vide_sel;

architecture Behavioral of ROM_vide_sel is

type zone_memoire is array ((2**12)-1 downto 0) of std_logic_vector (7 downto 0);
constant ROM: zone_memoire := (
	0 => "11111111",
	1 => "11111111",
	2 => "11111111",
	3 => "11111111",
	4 => "11111111",
	5 => "11111111",
	6 => "11111111",
	7 => "11111111",
	8 => "11111111",
	9 => "11111111",
	10 => "11111111",
	11 => "11111111",
	12 => "11111111",
	13 => "11111111",
	14 => "11111111",
	15 => "11111111",
	16 => "11111111",
	17 => "11111111",
	18 => "11111111",
	19 => "11111111",
	20 => "11111111",
	21 => "11111111",
	22 => "11111111",
	23 => "11111111",
	24 => "11111111",
	25 => "11111111",
	26 => "11111111",
	27 => "11111111",
	28 => "11111111",
	29 => "11111111",
	30 => "11111111",
	31 => "11111111",
	32 => "11111111",
	33 => "11111111",
	34 => "11111111",
	35 => "11111111",
	36 => "11111111",
	37 => "11111111",
	38 => "11111111",
	39 => "11111111",
	40 => "11111111",
	41 => "11111111",
	42 => "11111111",
	43 => "11111111",
	44 => "11111111",
	45 => "11111111",
	46 => "11111111",
	47 => "11111111",
	48 => "11111111",
	49 => "11111111",
	50 => "11111111",
	51 => "11111111",
	52 => "11111111",
	53 => "11111111",
	54 => "11111111",
	55 => "11111111",
	56 => "11111111",
	57 => "11111111",
	58 => "11111111",
	59 => "11111111",
	64 => "11111111",
	65 => "11111111",
	66 => "11111111",
	67 => "11111111",
	68 => "11111111",
	69 => "11111111",
	70 => "11111111",
	71 => "11111111",
	72 => "11111111",
	73 => "11111111",
	74 => "11111111",
	75 => "11111111",
	76 => "11111111",
	77 => "11111111",
	78 => "11111111",
	79 => "11111111",
	80 => "11111111",
	81 => "11111111",
	82 => "11111111",
	83 => "11111111",
	84 => "11111111",
	85 => "11111111",
	86 => "11111111",
	87 => "11111111",
	88 => "11111111",
	89 => "11111111",
	90 => "11111111",
	91 => "11111111",
	92 => "11111111",
	93 => "11111111",
	94 => "11111111",
	95 => "11111111",
	96 => "11111111",
	97 => "11111111",
	98 => "11111111",
	99 => "11111111",
	100 => "11111111",
	101 => "11111111",
	102 => "11111111",
	103 => "11111111",
	104 => "11111111",
	105 => "11111111",
	106 => "11111111",
	107 => "11111111",
	108 => "11111111",
	109 => "11111111",
	110 => "11111111",
	111 => "11111111",
	112 => "11111111",
	113 => "11111111",
	114 => "11111111",
	115 => "11111111",
	116 => "11111111",
	117 => "11111111",
	118 => "11111111",
	119 => "11111111",
	120 => "11111111",
	121 => "11111111",
	122 => "11111111",
	123 => "11111111",
	128 => "11111111",
	129 => "11111111",
	130 => "11111111",
	131 => "11111111",
	132 => "11111111",
	133 => "11111111",
	134 => "11111111",
	135 => "11111111",
	136 => "11111111",
	137 => "11111111",
	138 => "11111111",
	139 => "11111111",
	140 => "11111111",
	141 => "11111111",
	142 => "11111111",
	143 => "11111111",
	144 => "11111111",
	145 => "11111111",
	146 => "11111111",
	147 => "11111111",
	148 => "11111111",
	149 => "11111111",
	150 => "11111111",
	151 => "11111111",
	152 => "11111111",
	153 => "11111111",
	154 => "11111111",
	155 => "11111111",
	156 => "11111111",
	157 => "11111111",
	158 => "11111111",
	159 => "11111111",
	160 => "11111111",
	161 => "11111111",
	162 => "11111111",
	163 => "11111111",
	164 => "11111111",
	165 => "11111111",
	166 => "11111111",
	167 => "11111111",
	168 => "11111111",
	169 => "11111111",
	170 => "11111111",
	171 => "11111111",
	172 => "11111111",
	173 => "11111111",
	174 => "11111111",
	175 => "11111111",
	176 => "11111111",
	177 => "11111111",
	178 => "11111111",
	179 => "11111111",
	180 => "11111111",
	181 => "11111111",
	182 => "11111111",
	183 => "11111111",
	184 => "11111111",
	185 => "11111111",
	186 => "11111111",
	187 => "11111111",
	192 => "11111111",
	193 => "11111111",
	194 => "11111111",
	195 => "11111111",
	196 => "11111111",
	197 => "11111111",
	198 => "11111111",
	199 => "11111111",
	200 => "11111111",
	201 => "11111111",
	202 => "11111111",
	203 => "11111111",
	204 => "11111111",
	205 => "11111111",
	206 => "11111111",
	207 => "11111111",
	208 => "11111111",
	209 => "11111111",
	210 => "11111111",
	211 => "11111111",
	212 => "11111111",
	213 => "11111111",
	214 => "11111111",
	215 => "11111111",
	216 => "11111111",
	217 => "11111111",
	218 => "11111111",
	219 => "11111111",
	220 => "11111111",
	221 => "11111111",
	222 => "11111111",
	223 => "11111111",
	224 => "11111111",
	225 => "11111111",
	226 => "11111111",
	227 => "11111111",
	228 => "11111111",
	229 => "11111111",
	230 => "11111111",
	231 => "11111111",
	232 => "11111111",
	233 => "11111111",
	234 => "11111111",
	235 => "11111111",
	236 => "11111111",
	237 => "11111111",
	238 => "11111111",
	239 => "11111111",
	240 => "11111111",
	241 => "11111111",
	242 => "11111111",
	243 => "11111111",
	244 => "11111111",
	245 => "11111111",
	246 => "11111111",
	247 => "11111111",
	248 => "11111111",
	249 => "11111111",
	250 => "11111111",
	251 => "11111111",
	256 => "11111111",
	257 => "11111111",
	258 => "11111111",
	259 => "11111111",
	260 => "11111111",
	261 => "11111111",
	262 => "11111111",
	263 => "11111111",
	264 => "11111111",
	265 => "11111111",
	266 => "11111111",
	267 => "11111111",
	268 => "11111111",
	269 => "11111111",
	270 => "11111111",
	271 => "11111111",
	272 => "11111111",
	273 => "11111111",
	274 => "11111111",
	275 => "11111111",
	276 => "11111111",
	277 => "11111111",
	278 => "11111111",
	279 => "11111111",
	280 => "11111111",
	281 => "11111111",
	282 => "11111111",
	283 => "11111111",
	284 => "11111111",
	285 => "11111111",
	286 => "11111111",
	287 => "11111111",
	288 => "11111111",
	289 => "11111111",
	290 => "11111111",
	291 => "11111111",
	292 => "11111111",
	293 => "11111111",
	294 => "11111111",
	295 => "11111111",
	296 => "11111111",
	297 => "11111111",
	298 => "11111111",
	299 => "11111111",
	300 => "11111111",
	301 => "11111111",
	302 => "11111111",
	303 => "11111111",
	304 => "11111111",
	305 => "11111111",
	306 => "11111111",
	307 => "11111111",
	308 => "11111111",
	309 => "11111111",
	310 => "11111111",
	311 => "11111111",
	312 => "11111111",
	313 => "11111111",
	314 => "11111111",
	315 => "11111111",
	320 => "11111111",
	321 => "11111111",
	322 => "11111111",
	323 => "11111111",
	324 => "11111111",
	325 => "11111111",
	326 => "11111111",
	327 => "11111111",
	328 => "11111111",
	329 => "11111111",
	330 => "11111111",
	331 => "11111111",
	332 => "11111111",
	333 => "11111111",
	334 => "11111111",
	335 => "11111111",
	336 => "11111111",
	337 => "11111111",
	338 => "11111111",
	339 => "11111111",
	340 => "11111111",
	341 => "11111111",
	342 => "11111111",
	343 => "11111111",
	344 => "11111111",
	345 => "11111111",
	346 => "11111111",
	347 => "11111111",
	348 => "11111111",
	349 => "11111111",
	350 => "11111111",
	351 => "11111111",
	352 => "11111111",
	353 => "11111111",
	354 => "11111111",
	355 => "11111111",
	356 => "11111111",
	357 => "11111111",
	358 => "11111111",
	359 => "11111111",
	360 => "11111111",
	361 => "11111111",
	362 => "11111111",
	363 => "11111111",
	364 => "11111111",
	365 => "11111111",
	366 => "11111111",
	367 => "11111111",
	368 => "11111111",
	369 => "11111111",
	370 => "11111111",
	371 => "11111111",
	372 => "11111111",
	373 => "11111111",
	374 => "11111111",
	375 => "11111111",
	376 => "11111111",
	377 => "11111111",
	378 => "11111111",
	379 => "11111111",
	384 => "11111111",
	385 => "11111111",
	386 => "11111111",
	387 => "11111111",
	388 => "11111111",
	389 => "11111111",
	390 => "11111111",
	391 => "11111111",
	392 => "11111111",
	393 => "11111111",
	394 => "11111111",
	395 => "11111111",
	396 => "11111111",
	397 => "11111111",
	398 => "11111111",
	399 => "11111111",
	400 => "11111111",
	401 => "11111111",
	402 => "11111111",
	403 => "11111111",
	404 => "11111111",
	405 => "11111111",
	406 => "11111111",
	407 => "11111111",
	408 => "11111111",
	409 => "11111111",
	410 => "11111111",
	411 => "11111111",
	412 => "11111111",
	413 => "11111111",
	414 => "11111111",
	415 => "11111111",
	416 => "11111111",
	417 => "11111111",
	418 => "11111111",
	419 => "11111111",
	420 => "11111111",
	421 => "11111111",
	422 => "11111111",
	423 => "11111111",
	424 => "11111111",
	425 => "11111111",
	426 => "11111111",
	427 => "11111111",
	428 => "11111111",
	429 => "11111111",
	430 => "11111111",
	431 => "11111111",
	432 => "11111111",
	433 => "11111111",
	434 => "11111111",
	435 => "11111111",
	436 => "11111111",
	437 => "11111111",
	438 => "11111111",
	439 => "11111111",
	440 => "11111111",
	441 => "11111111",
	442 => "11111111",
	443 => "11111111",
	448 => "11111111",
	449 => "11111111",
	450 => "11111111",
	451 => "11111111",
	452 => "11111111",
	453 => "11111111",
	454 => "11111111",
	455 => "11111111",
	456 => "11111111",
	457 => "11111111",
	458 => "11111111",
	459 => "11111111",
	460 => "11111111",
	461 => "11111111",
	462 => "11111111",
	463 => "11111111",
	464 => "11111111",
	465 => "11111111",
	466 => "11111111",
	467 => "11111111",
	468 => "11111111",
	469 => "11111111",
	470 => "11111111",
	471 => "11111111",
	472 => "11111111",
	473 => "11111111",
	474 => "11111111",
	475 => "11111111",
	476 => "11111111",
	477 => "11111111",
	478 => "11111111",
	479 => "11111111",
	480 => "11111111",
	481 => "11111111",
	482 => "11111111",
	483 => "11111111",
	484 => "11111111",
	485 => "11111111",
	486 => "11111111",
	487 => "11111111",
	488 => "11111111",
	489 => "11111111",
	490 => "11111111",
	491 => "11111111",
	492 => "11111111",
	493 => "11111111",
	494 => "11111111",
	495 => "11111111",
	496 => "11111111",
	497 => "11111111",
	498 => "11111111",
	499 => "11111111",
	500 => "11111111",
	501 => "11111111",
	502 => "11111111",
	503 => "11111111",
	504 => "11111111",
	505 => "11111111",
	506 => "11111111",
	507 => "11111111",
	512 => "11111111",
	513 => "11111111",
	514 => "11111111",
	515 => "11111111",
	516 => "11111111",
	517 => "11111111",
	518 => "11111111",
	519 => "11111111",
	520 => "11111111",
	521 => "11111111",
	522 => "11111111",
	523 => "11111111",
	524 => "11111111",
	525 => "11111111",
	526 => "11111111",
	527 => "11111111",
	528 => "11111111",
	529 => "11111111",
	530 => "11111111",
	531 => "11111111",
	532 => "11111111",
	533 => "11111111",
	534 => "11111111",
	535 => "11111111",
	536 => "11111111",
	537 => "11111111",
	538 => "11111111",
	539 => "11111111",
	540 => "11111111",
	541 => "11111111",
	542 => "11111111",
	543 => "11111111",
	544 => "11111111",
	545 => "11111111",
	546 => "11111111",
	547 => "11111111",
	548 => "11111111",
	549 => "11111111",
	550 => "11111111",
	551 => "11111111",
	552 => "11111111",
	553 => "11111111",
	554 => "11111111",
	555 => "11111111",
	556 => "11111111",
	557 => "11111111",
	558 => "11111111",
	559 => "11111111",
	560 => "11111111",
	561 => "11111111",
	562 => "11111111",
	563 => "11111111",
	564 => "11111111",
	565 => "11111111",
	566 => "11111111",
	567 => "11111111",
	568 => "11111111",
	569 => "11111111",
	570 => "11111111",
	571 => "11111111",
	576 => "11111111",
	577 => "11111111",
	578 => "11111111",
	579 => "11111111",
	580 => "11111111",
	581 => "11111111",
	582 => "11111111",
	583 => "11111111",
	584 => "11111111",
	585 => "11111111",
	586 => "11111111",
	587 => "11111111",
	588 => "11111111",
	589 => "11111111",
	590 => "11111111",
	591 => "11111111",
	592 => "11111111",
	593 => "11111111",
	594 => "11111111",
	595 => "11111111",
	596 => "11111111",
	597 => "11111111",
	598 => "11111111",
	599 => "11111111",
	600 => "11111111",
	601 => "11111111",
	602 => "11111111",
	603 => "11111111",
	604 => "11111111",
	605 => "11111111",
	606 => "11111111",
	607 => "11111111",
	608 => "11111111",
	609 => "11111111",
	610 => "11111111",
	611 => "11111111",
	612 => "11111111",
	613 => "11111111",
	614 => "11111111",
	615 => "11111111",
	616 => "11111111",
	617 => "11111111",
	618 => "11111111",
	619 => "11111111",
	620 => "11111111",
	621 => "11111111",
	622 => "11111111",
	623 => "11111111",
	624 => "11111111",
	625 => "11111111",
	626 => "11111111",
	627 => "11111111",
	628 => "11111111",
	629 => "11111111",
	630 => "11111111",
	631 => "11111111",
	632 => "11111111",
	633 => "11111111",
	634 => "11111111",
	635 => "11111111",
	640 => "11111111",
	641 => "11111111",
	642 => "11111111",
	643 => "11111111",
	644 => "11111111",
	645 => "11111111",
	646 => "11111111",
	647 => "11111111",
	648 => "11111111",
	649 => "11111111",
	650 => "11111111",
	651 => "11111111",
	652 => "11111111",
	653 => "11111111",
	654 => "11111111",
	655 => "11111111",
	656 => "11111111",
	657 => "11111111",
	658 => "11111111",
	659 => "11111111",
	660 => "11111111",
	661 => "11111111",
	662 => "11111111",
	663 => "11111111",
	664 => "11111111",
	665 => "11111111",
	666 => "11111111",
	667 => "11111111",
	668 => "11111111",
	669 => "11111111",
	670 => "11111111",
	671 => "11111111",
	672 => "11111111",
	673 => "11111111",
	674 => "11111111",
	675 => "11111111",
	676 => "11111111",
	677 => "11111111",
	678 => "11111111",
	679 => "11111111",
	680 => "11111111",
	681 => "11111111",
	682 => "11111111",
	683 => "11111111",
	684 => "11111111",
	685 => "11111111",
	686 => "11111111",
	687 => "11111111",
	688 => "11111111",
	689 => "11111111",
	690 => "11111111",
	691 => "11111111",
	692 => "11111111",
	693 => "11111111",
	694 => "11111111",
	695 => "11111111",
	696 => "11111111",
	697 => "11111111",
	698 => "11111111",
	699 => "11111111",
	704 => "11111111",
	705 => "11111111",
	706 => "11111111",
	707 => "11111111",
	708 => "11111111",
	709 => "11111111",
	710 => "11111111",
	711 => "11111111",
	712 => "11111111",
	713 => "11111111",
	714 => "11111111",
	715 => "11111111",
	716 => "11111111",
	717 => "11111111",
	718 => "11111111",
	719 => "11111111",
	720 => "11111111",
	721 => "11111111",
	722 => "11111111",
	723 => "11111111",
	724 => "11111111",
	725 => "11111111",
	726 => "11111111",
	727 => "11111111",
	728 => "11111111",
	729 => "11111111",
	730 => "11111111",
	731 => "11111111",
	732 => "11111111",
	733 => "11111111",
	734 => "11111111",
	735 => "11111111",
	736 => "11111111",
	737 => "11111111",
	738 => "11111111",
	739 => "11111111",
	740 => "11111111",
	741 => "11111111",
	742 => "11111111",
	743 => "11111111",
	744 => "11111111",
	745 => "11111111",
	746 => "11111111",
	747 => "11111111",
	748 => "11111111",
	749 => "11111111",
	750 => "11111111",
	751 => "11111111",
	752 => "11111111",
	753 => "11111111",
	754 => "11111111",
	755 => "11111111",
	756 => "11111111",
	757 => "11111111",
	758 => "11111111",
	759 => "11111111",
	760 => "11111111",
	761 => "11111111",
	762 => "11111111",
	763 => "11111111",
	768 => "11111111",
	769 => "11111111",
	770 => "11111111",
	771 => "11111111",
	772 => "11111111",
	773 => "11111111",
	774 => "11111111",
	775 => "11111111",
	776 => "11111111",
	777 => "11111111",
	778 => "11111111",
	779 => "11111111",
	780 => "11111111",
	781 => "11111111",
	782 => "11111111",
	783 => "11111111",
	784 => "11111111",
	785 => "11111111",
	786 => "11111111",
	787 => "11111111",
	788 => "11111111",
	789 => "11111111",
	790 => "11111111",
	791 => "11111111",
	792 => "11111111",
	793 => "11111111",
	794 => "11111111",
	795 => "11111111",
	796 => "11111111",
	797 => "11111111",
	798 => "11111111",
	799 => "11111111",
	800 => "11111111",
	801 => "11111111",
	802 => "11111111",
	803 => "11111111",
	804 => "11111111",
	805 => "11111111",
	806 => "11111111",
	807 => "11111111",
	808 => "11111111",
	809 => "11111111",
	810 => "11111111",
	811 => "11111111",
	812 => "11111111",
	813 => "11111111",
	814 => "11111111",
	815 => "11111111",
	816 => "11111111",
	817 => "11111111",
	818 => "11111111",
	819 => "11111111",
	820 => "11111111",
	821 => "11111111",
	822 => "11111111",
	823 => "11111111",
	824 => "11111111",
	825 => "11111111",
	826 => "11111111",
	827 => "11111111",
	832 => "11111111",
	833 => "11111111",
	834 => "11111111",
	835 => "11111111",
	836 => "11111111",
	837 => "11111111",
	838 => "11111111",
	839 => "11111111",
	840 => "11111111",
	841 => "11111111",
	842 => "11111111",
	843 => "11111111",
	844 => "11111111",
	845 => "11111111",
	846 => "11111111",
	847 => "11111111",
	848 => "11111111",
	849 => "11111111",
	850 => "11111111",
	851 => "11111111",
	852 => "11111111",
	853 => "11111111",
	854 => "11111111",
	855 => "11111111",
	856 => "11111111",
	857 => "11111111",
	858 => "11111111",
	859 => "11111111",
	860 => "11111111",
	861 => "11111111",
	862 => "11111111",
	863 => "11111111",
	864 => "11111111",
	865 => "11111111",
	866 => "11111111",
	867 => "11111111",
	868 => "11111111",
	869 => "11111111",
	870 => "11111111",
	871 => "11111111",
	872 => "11111111",
	873 => "11111111",
	874 => "11111111",
	875 => "11111111",
	876 => "11111111",
	877 => "11111111",
	878 => "11111111",
	879 => "11111111",
	880 => "11111111",
	881 => "11111111",
	882 => "11111111",
	883 => "11111111",
	884 => "11111111",
	885 => "11111111",
	886 => "11111111",
	887 => "11111111",
	888 => "11111111",
	889 => "11111111",
	890 => "11111111",
	891 => "11111111",
	896 => "11111111",
	897 => "11111111",
	898 => "11111111",
	899 => "11111111",
	900 => "11111111",
	901 => "11111111",
	902 => "11111111",
	903 => "11111111",
	904 => "11111111",
	905 => "11111111",
	906 => "11111111",
	907 => "11111111",
	908 => "11111111",
	909 => "11111111",
	910 => "11111111",
	911 => "11111111",
	912 => "11111111",
	913 => "11111111",
	914 => "11111111",
	915 => "11111111",
	916 => "11111111",
	917 => "11111111",
	918 => "11111111",
	919 => "11111111",
	920 => "11111111",
	921 => "11111111",
	922 => "11111111",
	923 => "11111111",
	924 => "11111111",
	925 => "11111111",
	926 => "11111111",
	927 => "11111111",
	928 => "11111111",
	929 => "11111111",
	930 => "11111111",
	931 => "11111111",
	932 => "11111111",
	933 => "11111111",
	934 => "11111111",
	935 => "11111111",
	936 => "11111111",
	937 => "11111111",
	938 => "11111111",
	939 => "11111111",
	940 => "11111111",
	941 => "11111111",
	942 => "11111111",
	943 => "11111111",
	944 => "11111111",
	945 => "11111111",
	946 => "11111111",
	947 => "11111111",
	948 => "11111111",
	949 => "11111111",
	950 => "11111111",
	951 => "11111111",
	952 => "11111111",
	953 => "11111111",
	954 => "11111111",
	955 => "11111111",
	960 => "11111111",
	961 => "11111111",
	962 => "11111111",
	963 => "11111111",
	964 => "11111111",
	965 => "11111111",
	966 => "11111111",
	967 => "11111111",
	968 => "11111111",
	969 => "11111111",
	970 => "11111111",
	971 => "11111111",
	972 => "11111111",
	973 => "11111111",
	974 => "11111111",
	975 => "11111111",
	976 => "11111111",
	977 => "11111111",
	978 => "11111111",
	979 => "11111111",
	980 => "11111111",
	981 => "11111111",
	982 => "11111111",
	983 => "11111111",
	984 => "11111111",
	985 => "11111111",
	986 => "11111111",
	987 => "11111111",
	988 => "11111111",
	989 => "11111111",
	990 => "11111111",
	991 => "11111111",
	992 => "11111111",
	993 => "11111111",
	994 => "11111111",
	995 => "11111111",
	996 => "11111111",
	997 => "11111111",
	998 => "11111111",
	999 => "11111111",
	1000 => "11111111",
	1001 => "11111111",
	1002 => "11111111",
	1003 => "11111111",
	1004 => "11111111",
	1005 => "11111111",
	1006 => "11111111",
	1007 => "11111111",
	1008 => "11111111",
	1009 => "11111111",
	1010 => "11111111",
	1011 => "11111111",
	1012 => "11111111",
	1013 => "11111111",
	1014 => "11111111",
	1015 => "11111111",
	1016 => "11111111",
	1017 => "11111111",
	1018 => "11111111",
	1019 => "11111111",
	1024 => "11111111",
	1025 => "11111111",
	1026 => "11111111",
	1027 => "11111111",
	1028 => "11111111",
	1029 => "11111111",
	1030 => "11111111",
	1031 => "11111111",
	1032 => "11111111",
	1033 => "11111111",
	1034 => "11111111",
	1035 => "11111111",
	1036 => "11111111",
	1037 => "11111111",
	1038 => "11111111",
	1039 => "11111111",
	1040 => "11111111",
	1041 => "11111111",
	1042 => "11111111",
	1043 => "11111111",
	1044 => "11111111",
	1045 => "11111111",
	1046 => "11111111",
	1047 => "11111111",
	1048 => "11111111",
	1049 => "11111111",
	1050 => "11111111",
	1051 => "11111111",
	1052 => "11111111",
	1053 => "11111111",
	1054 => "11111111",
	1055 => "11111111",
	1056 => "11111111",
	1057 => "11111111",
	1058 => "11111111",
	1059 => "11111111",
	1060 => "11111111",
	1061 => "11111111",
	1062 => "11111111",
	1063 => "11111111",
	1064 => "11111111",
	1065 => "11111111",
	1066 => "11111111",
	1067 => "11111111",
	1068 => "11111111",
	1069 => "11111111",
	1070 => "11111111",
	1071 => "11111111",
	1072 => "11111111",
	1073 => "11111111",
	1074 => "11111111",
	1075 => "11111111",
	1076 => "11111111",
	1077 => "11111111",
	1078 => "11111111",
	1079 => "11111111",
	1080 => "11111111",
	1081 => "11111111",
	1082 => "11111111",
	1083 => "11111111",
	1088 => "11111111",
	1089 => "11111111",
	1090 => "11111111",
	1091 => "11111111",
	1092 => "11111111",
	1093 => "11111111",
	1094 => "11111111",
	1095 => "11111111",
	1096 => "11111111",
	1097 => "11111111",
	1098 => "11111111",
	1099 => "11111111",
	1100 => "11111111",
	1101 => "11111111",
	1102 => "11111111",
	1103 => "11111111",
	1104 => "11111111",
	1105 => "11111111",
	1106 => "11111111",
	1107 => "11111111",
	1108 => "11111111",
	1109 => "11111111",
	1110 => "11111111",
	1111 => "11111111",
	1112 => "11111111",
	1113 => "11111111",
	1114 => "11111111",
	1115 => "11111111",
	1116 => "11111111",
	1117 => "11111111",
	1118 => "11111111",
	1119 => "11111111",
	1120 => "11111111",
	1121 => "11111111",
	1122 => "11111111",
	1123 => "11111111",
	1124 => "11111111",
	1125 => "11111111",
	1126 => "11111111",
	1127 => "11111111",
	1128 => "11111111",
	1129 => "11111111",
	1130 => "11111111",
	1131 => "11111111",
	1132 => "11111111",
	1133 => "11111111",
	1134 => "11111111",
	1135 => "11111111",
	1136 => "11111111",
	1137 => "11111111",
	1138 => "11111111",
	1139 => "11111111",
	1140 => "11111111",
	1141 => "11111111",
	1142 => "11111111",
	1143 => "11111111",
	1144 => "11111111",
	1145 => "11111111",
	1146 => "11111111",
	1147 => "11111111",
	1152 => "11111111",
	1153 => "11111111",
	1154 => "11111111",
	1155 => "11111111",
	1156 => "11111111",
	1157 => "11111111",
	1158 => "11111111",
	1159 => "11111111",
	1160 => "11111111",
	1161 => "11111111",
	1162 => "11111111",
	1163 => "11111111",
	1164 => "11111111",
	1165 => "11111111",
	1166 => "11111111",
	1167 => "11111111",
	1168 => "11111111",
	1169 => "11111111",
	1170 => "11111111",
	1171 => "11111111",
	1172 => "11111111",
	1173 => "11111111",
	1174 => "11111111",
	1175 => "11111111",
	1176 => "11111111",
	1177 => "11111111",
	1178 => "11111111",
	1179 => "11111111",
	1180 => "11111111",
	1181 => "11111111",
	1182 => "11111111",
	1183 => "11111111",
	1184 => "11111111",
	1185 => "11111111",
	1186 => "11111111",
	1187 => "11111111",
	1188 => "11111111",
	1189 => "11111111",
	1190 => "11111111",
	1191 => "11111111",
	1192 => "11111111",
	1193 => "11111111",
	1194 => "11111111",
	1195 => "11111111",
	1196 => "11111111",
	1197 => "11111111",
	1198 => "11111111",
	1199 => "11111111",
	1200 => "11111111",
	1201 => "11111111",
	1202 => "11111111",
	1203 => "11111111",
	1204 => "11111111",
	1205 => "11111111",
	1206 => "11111111",
	1207 => "11111111",
	1208 => "11111111",
	1209 => "11111111",
	1210 => "11111111",
	1211 => "11111111",
	1216 => "11111111",
	1217 => "11111111",
	1218 => "11111111",
	1219 => "11111111",
	1220 => "11111111",
	1221 => "11111111",
	1222 => "11111111",
	1223 => "11111111",
	1224 => "11111111",
	1225 => "11111111",
	1226 => "11111111",
	1227 => "11111111",
	1228 => "11111111",
	1229 => "11111111",
	1230 => "11111111",
	1231 => "11111111",
	1232 => "11111111",
	1233 => "11111111",
	1234 => "11111111",
	1235 => "11111111",
	1236 => "11111111",
	1237 => "11111111",
	1238 => "11111111",
	1239 => "11111111",
	1240 => "11111111",
	1241 => "11111111",
	1242 => "11111111",
	1243 => "11111111",
	1244 => "11111111",
	1245 => "11111111",
	1246 => "11111111",
	1247 => "11111111",
	1248 => "11111111",
	1249 => "11111111",
	1250 => "11111111",
	1251 => "11111111",
	1252 => "11111111",
	1253 => "11111111",
	1254 => "11111111",
	1255 => "11111111",
	1256 => "11111111",
	1257 => "11111111",
	1258 => "11111111",
	1259 => "11111111",
	1260 => "11111111",
	1261 => "11111111",
	1262 => "11111111",
	1263 => "11111111",
	1264 => "11111111",
	1265 => "11111111",
	1266 => "11111111",
	1267 => "11111111",
	1268 => "11111111",
	1269 => "11111111",
	1270 => "11111111",
	1271 => "11111111",
	1272 => "11111111",
	1273 => "11111111",
	1274 => "11111111",
	1275 => "11111111",
	1280 => "11111111",
	1281 => "11111111",
	1282 => "11111111",
	1283 => "11111111",
	1284 => "11111111",
	1285 => "11111111",
	1286 => "11111111",
	1287 => "11111111",
	1288 => "11111111",
	1289 => "11111111",
	1290 => "11111111",
	1291 => "11111111",
	1292 => "11111111",
	1293 => "11111111",
	1294 => "11111111",
	1295 => "11111111",
	1296 => "11111111",
	1297 => "11111111",
	1298 => "11111111",
	1299 => "11111111",
	1300 => "11111111",
	1301 => "11111111",
	1302 => "11111111",
	1303 => "11111111",
	1304 => "11111111",
	1305 => "11111111",
	1306 => "11111111",
	1307 => "11111111",
	1308 => "11111111",
	1309 => "11111111",
	1310 => "11111111",
	1311 => "11111111",
	1312 => "11111111",
	1313 => "11111111",
	1314 => "11111111",
	1315 => "11111111",
	1316 => "11111111",
	1317 => "11111111",
	1318 => "11111111",
	1319 => "11111111",
	1320 => "11111111",
	1321 => "11111111",
	1322 => "11111111",
	1323 => "11111111",
	1324 => "11111111",
	1325 => "11111111",
	1326 => "11111111",
	1327 => "11111111",
	1328 => "11111111",
	1329 => "11111111",
	1330 => "11111111",
	1331 => "11111111",
	1332 => "11111111",
	1333 => "11111111",
	1334 => "11111111",
	1335 => "11111111",
	1336 => "11111111",
	1337 => "11111111",
	1338 => "11111111",
	1339 => "11111111",
	1344 => "11111111",
	1345 => "11111111",
	1346 => "11111111",
	1347 => "11111111",
	1348 => "11111111",
	1349 => "11111111",
	1350 => "11111111",
	1351 => "11111111",
	1352 => "11111111",
	1353 => "11111111",
	1354 => "11111111",
	1355 => "11111111",
	1356 => "11111111",
	1357 => "11111111",
	1358 => "11111111",
	1359 => "11111111",
	1360 => "11111111",
	1361 => "11111111",
	1362 => "11111111",
	1363 => "11111111",
	1364 => "11111111",
	1365 => "11111111",
	1366 => "11111111",
	1367 => "11111111",
	1368 => "11111111",
	1369 => "11111111",
	1370 => "11111111",
	1371 => "11111111",
	1372 => "11111111",
	1373 => "11111111",
	1374 => "11111111",
	1375 => "11111111",
	1376 => "11111111",
	1377 => "11111111",
	1378 => "11111111",
	1379 => "11111111",
	1380 => "11111111",
	1381 => "11111111",
	1382 => "11111111",
	1383 => "11111111",
	1384 => "11111111",
	1385 => "11111111",
	1386 => "11111111",
	1387 => "11111111",
	1388 => "11111111",
	1389 => "11111111",
	1390 => "11111111",
	1391 => "11111111",
	1392 => "11111111",
	1393 => "11111111",
	1394 => "11111111",
	1395 => "11111111",
	1396 => "11111111",
	1397 => "11111111",
	1398 => "11111111",
	1399 => "11111111",
	1400 => "11111111",
	1401 => "11111111",
	1402 => "11111111",
	1403 => "11111111",
	1408 => "11111111",
	1409 => "11111111",
	1410 => "11111111",
	1411 => "11111111",
	1412 => "11111111",
	1413 => "11111111",
	1414 => "11111111",
	1415 => "11111111",
	1416 => "11111111",
	1417 => "11111111",
	1418 => "11111111",
	1419 => "11111111",
	1420 => "11111111",
	1421 => "11111111",
	1422 => "11111111",
	1423 => "11111111",
	1424 => "11111111",
	1425 => "11111111",
	1426 => "11111111",
	1427 => "11111111",
	1428 => "11111111",
	1429 => "11111111",
	1430 => "11111111",
	1431 => "11111111",
	1432 => "11111111",
	1433 => "11111111",
	1434 => "11111111",
	1435 => "11111111",
	1436 => "11111111",
	1437 => "11111111",
	1438 => "11111111",
	1439 => "11111111",
	1440 => "11111111",
	1441 => "11111111",
	1442 => "11111111",
	1443 => "11111111",
	1444 => "11111111",
	1445 => "11111111",
	1446 => "11111111",
	1447 => "11111111",
	1448 => "11111111",
	1449 => "11111111",
	1450 => "11111111",
	1451 => "11111111",
	1452 => "11111111",
	1453 => "11111111",
	1454 => "11111111",
	1455 => "11111111",
	1456 => "11111111",
	1457 => "11111111",
	1458 => "11111111",
	1459 => "11111111",
	1460 => "11111111",
	1461 => "11111111",
	1462 => "11111111",
	1463 => "11111111",
	1464 => "11111111",
	1465 => "11111111",
	1466 => "11111111",
	1467 => "11111111",
	1472 => "11111111",
	1473 => "11111111",
	1474 => "11111111",
	1475 => "11111111",
	1476 => "11111111",
	1477 => "11111111",
	1478 => "11111111",
	1479 => "11111111",
	1480 => "11111111",
	1481 => "11111111",
	1482 => "11111111",
	1483 => "11111111",
	1484 => "11111111",
	1485 => "11111111",
	1486 => "11111111",
	1487 => "11111111",
	1488 => "11111111",
	1489 => "11111111",
	1490 => "11111111",
	1491 => "11111111",
	1492 => "11111111",
	1493 => "11111111",
	1494 => "11111111",
	1495 => "11111111",
	1496 => "11111111",
	1497 => "11111111",
	1498 => "11111111",
	1499 => "11111111",
	1500 => "11111111",
	1501 => "11111111",
	1502 => "11111111",
	1503 => "11111111",
	1504 => "11111111",
	1505 => "11111111",
	1506 => "11111111",
	1507 => "11111111",
	1508 => "11111111",
	1509 => "11111111",
	1510 => "11111111",
	1511 => "11111111",
	1512 => "11111111",
	1513 => "11111111",
	1514 => "11111111",
	1515 => "11111111",
	1516 => "11111111",
	1517 => "11111111",
	1518 => "11111111",
	1519 => "11111111",
	1520 => "11111111",
	1521 => "11111111",
	1522 => "11111111",
	1523 => "11111111",
	1524 => "11111111",
	1525 => "11111111",
	1526 => "11111111",
	1527 => "11111111",
	1528 => "11111111",
	1529 => "11111111",
	1530 => "11111111",
	1531 => "11111111",
	1536 => "11111111",
	1537 => "11111111",
	1538 => "11111111",
	1539 => "11111111",
	1540 => "11111111",
	1541 => "11111111",
	1542 => "11111111",
	1543 => "11111111",
	1544 => "11111111",
	1545 => "11111111",
	1546 => "11111111",
	1547 => "11111111",
	1548 => "11111111",
	1549 => "11111111",
	1550 => "11111111",
	1551 => "11111111",
	1552 => "11111111",
	1553 => "11111111",
	1554 => "11111111",
	1555 => "11111111",
	1556 => "11111111",
	1557 => "11111111",
	1558 => "11111111",
	1559 => "11111111",
	1560 => "11111111",
	1561 => "11111111",
	1562 => "11111111",
	1563 => "11111111",
	1564 => "11111111",
	1565 => "11111111",
	1566 => "11111111",
	1567 => "11111111",
	1568 => "11111111",
	1569 => "11111111",
	1570 => "11111111",
	1571 => "11111111",
	1572 => "11111111",
	1573 => "11111111",
	1574 => "11111111",
	1575 => "11111111",
	1576 => "11111111",
	1577 => "11111111",
	1578 => "11111111",
	1579 => "11111111",
	1580 => "11111111",
	1581 => "11111111",
	1582 => "11111111",
	1583 => "11111111",
	1584 => "11111111",
	1585 => "11111111",
	1586 => "11111111",
	1587 => "11111111",
	1588 => "11111111",
	1589 => "11111111",
	1590 => "11111111",
	1591 => "11111111",
	1592 => "11111111",
	1593 => "11111111",
	1594 => "11111111",
	1595 => "11111111",
	1600 => "11111111",
	1601 => "11111111",
	1602 => "11111111",
	1603 => "11111111",
	1604 => "11111111",
	1605 => "11111111",
	1606 => "11111111",
	1607 => "11111111",
	1608 => "11111111",
	1609 => "11111111",
	1610 => "11111111",
	1611 => "11111111",
	1612 => "11111111",
	1613 => "11111111",
	1614 => "11111111",
	1615 => "11111111",
	1616 => "11111111",
	1617 => "11111111",
	1618 => "11111111",
	1619 => "11111111",
	1620 => "11111111",
	1621 => "11111111",
	1622 => "11111111",
	1623 => "11111111",
	1624 => "11111111",
	1625 => "11111111",
	1626 => "11111111",
	1627 => "11111111",
	1628 => "11111111",
	1629 => "11111111",
	1630 => "11111111",
	1631 => "11111111",
	1632 => "11111111",
	1633 => "11111111",
	1634 => "11111111",
	1635 => "11111111",
	1636 => "11111111",
	1637 => "11111111",
	1638 => "11111111",
	1639 => "11111111",
	1640 => "11111111",
	1641 => "11111111",
	1642 => "11111111",
	1643 => "11111111",
	1644 => "11111111",
	1645 => "11111111",
	1646 => "11111111",
	1647 => "11111111",
	1648 => "11111111",
	1649 => "11111111",
	1650 => "11111111",
	1651 => "11111111",
	1652 => "11111111",
	1653 => "11111111",
	1654 => "11111111",
	1655 => "11111111",
	1656 => "11111111",
	1657 => "11111111",
	1658 => "11111111",
	1659 => "11111111",
	1664 => "11111111",
	1665 => "11111111",
	1666 => "11111111",
	1667 => "11111111",
	1668 => "11111111",
	1669 => "11111111",
	1670 => "11111111",
	1671 => "11111111",
	1672 => "11111111",
	1673 => "11111111",
	1674 => "11111111",
	1675 => "11111111",
	1676 => "11111111",
	1677 => "11111111",
	1678 => "11111111",
	1679 => "11111111",
	1680 => "11111111",
	1681 => "11111111",
	1682 => "11111111",
	1683 => "11111111",
	1684 => "11111111",
	1685 => "11111111",
	1686 => "11111111",
	1687 => "11111111",
	1688 => "11111111",
	1689 => "11111111",
	1690 => "11111111",
	1691 => "11111111",
	1692 => "11111111",
	1693 => "11111111",
	1694 => "11111111",
	1695 => "11111111",
	1696 => "11111111",
	1697 => "11111111",
	1698 => "11111111",
	1699 => "11111111",
	1700 => "11111111",
	1701 => "11111111",
	1702 => "11111111",
	1703 => "11111111",
	1704 => "11111111",
	1705 => "11111111",
	1706 => "11111111",
	1707 => "11111111",
	1708 => "11111111",
	1709 => "11111111",
	1710 => "11111111",
	1711 => "11111111",
	1712 => "11111111",
	1713 => "11111111",
	1714 => "11111111",
	1715 => "11111111",
	1716 => "11111111",
	1717 => "11111111",
	1718 => "11111111",
	1719 => "11111111",
	1720 => "11111111",
	1721 => "11111111",
	1722 => "11111111",
	1723 => "11111111",
	1728 => "11111111",
	1729 => "11111111",
	1730 => "11111111",
	1731 => "11111111",
	1732 => "11111111",
	1733 => "11111111",
	1734 => "11111111",
	1735 => "11111111",
	1736 => "11111111",
	1737 => "11111111",
	1738 => "11111111",
	1739 => "11111111",
	1740 => "11111111",
	1741 => "11111111",
	1742 => "11111111",
	1743 => "11111111",
	1744 => "11111111",
	1745 => "11111111",
	1746 => "11111111",
	1747 => "11111111",
	1748 => "11111111",
	1749 => "11111111",
	1750 => "11111111",
	1751 => "11111111",
	1752 => "11111111",
	1753 => "11111111",
	1754 => "11111111",
	1755 => "11111111",
	1756 => "11111111",
	1757 => "11111111",
	1758 => "11111111",
	1759 => "11111111",
	1760 => "11111111",
	1761 => "11111111",
	1762 => "11111111",
	1763 => "11111111",
	1764 => "11111111",
	1765 => "11111111",
	1766 => "11111111",
	1767 => "11111111",
	1768 => "11111111",
	1769 => "11111111",
	1770 => "11111111",
	1771 => "11111111",
	1772 => "11111111",
	1773 => "11111111",
	1774 => "11111111",
	1775 => "11111111",
	1776 => "11111111",
	1777 => "11111111",
	1778 => "11111111",
	1779 => "11111111",
	1780 => "11111111",
	1781 => "11111111",
	1782 => "11111111",
	1783 => "11111111",
	1784 => "11111111",
	1785 => "11111111",
	1786 => "11111111",
	1787 => "11111111",
	1792 => "11111111",
	1793 => "11111111",
	1794 => "11111111",
	1795 => "11111111",
	1796 => "11111111",
	1797 => "11111111",
	1798 => "11111111",
	1799 => "11111111",
	1800 => "11111111",
	1801 => "11111111",
	1802 => "11111111",
	1803 => "11111111",
	1804 => "11111111",
	1805 => "11111111",
	1806 => "11111111",
	1807 => "11111111",
	1808 => "11111111",
	1809 => "11111111",
	1810 => "11111111",
	1811 => "11111111",
	1812 => "11111111",
	1813 => "11111111",
	1814 => "11111111",
	1815 => "11111111",
	1816 => "11111111",
	1817 => "11111111",
	1818 => "11111111",
	1819 => "11111111",
	1820 => "11111111",
	1821 => "11111111",
	1822 => "11111111",
	1823 => "11111111",
	1824 => "11111111",
	1825 => "11111111",
	1826 => "11111111",
	1827 => "11111111",
	1828 => "11111111",
	1829 => "11111111",
	1830 => "11111111",
	1831 => "11111111",
	1832 => "11111111",
	1833 => "11111111",
	1834 => "11111111",
	1835 => "11111111",
	1836 => "11111111",
	1837 => "11111111",
	1838 => "11111111",
	1839 => "11111111",
	1840 => "11111111",
	1841 => "11111111",
	1842 => "11111111",
	1843 => "11111111",
	1844 => "11111111",
	1845 => "11111111",
	1846 => "11111111",
	1847 => "11111111",
	1848 => "11111111",
	1849 => "11111111",
	1850 => "11111111",
	1851 => "11111111",
	1856 => "11111111",
	1857 => "11111111",
	1858 => "11111111",
	1859 => "11111111",
	1860 => "11111111",
	1861 => "11111111",
	1862 => "11111111",
	1863 => "11111111",
	1864 => "11111111",
	1865 => "11111111",
	1866 => "11111111",
	1867 => "11111111",
	1868 => "11111111",
	1869 => "11111111",
	1870 => "11111111",
	1871 => "11111111",
	1872 => "11111111",
	1873 => "11111111",
	1874 => "11111111",
	1875 => "11111111",
	1876 => "11111111",
	1877 => "11111111",
	1878 => "11111111",
	1879 => "11111111",
	1880 => "11111111",
	1881 => "11111111",
	1882 => "11111111",
	1883 => "11111111",
	1884 => "11111111",
	1885 => "11111111",
	1886 => "11111111",
	1887 => "11111111",
	1888 => "11111111",
	1889 => "11111111",
	1890 => "11111111",
	1891 => "11111111",
	1892 => "11111111",
	1893 => "11111111",
	1894 => "11111111",
	1895 => "11111111",
	1896 => "11111111",
	1897 => "11111111",
	1898 => "11111111",
	1899 => "11111111",
	1900 => "11111111",
	1901 => "11111111",
	1902 => "11111111",
	1903 => "11111111",
	1904 => "11111111",
	1905 => "11111111",
	1906 => "11111111",
	1907 => "11111111",
	1908 => "11111111",
	1909 => "11111111",
	1910 => "11111111",
	1911 => "11111111",
	1912 => "11111111",
	1913 => "11111111",
	1914 => "11111111",
	1915 => "11111111",
	1920 => "11111111",
	1921 => "11111111",
	1922 => "11111111",
	1923 => "11111111",
	1924 => "11111111",
	1925 => "11111111",
	1926 => "11111111",
	1927 => "11111111",
	1928 => "11111111",
	1929 => "11111111",
	1930 => "11111111",
	1931 => "11111111",
	1932 => "11111111",
	1933 => "11111111",
	1934 => "11111111",
	1935 => "11111111",
	1936 => "11111111",
	1937 => "11111111",
	1938 => "11111111",
	1939 => "11111111",
	1940 => "11111111",
	1941 => "11111111",
	1942 => "11111111",
	1943 => "11111111",
	1944 => "11111111",
	1945 => "11111111",
	1946 => "11111111",
	1947 => "11111111",
	1948 => "11111111",
	1949 => "11111111",
	1950 => "11111111",
	1951 => "11111111",
	1952 => "11111111",
	1953 => "11111111",
	1954 => "11111111",
	1955 => "11111111",
	1956 => "11111111",
	1957 => "11111111",
	1958 => "11111111",
	1959 => "11111111",
	1960 => "11111111",
	1961 => "11111111",
	1962 => "11111111",
	1963 => "11111111",
	1964 => "11111111",
	1965 => "11111111",
	1966 => "11111111",
	1967 => "11111111",
	1968 => "11111111",
	1969 => "11111111",
	1970 => "11111111",
	1971 => "11111111",
	1972 => "11111111",
	1973 => "11111111",
	1974 => "11111111",
	1975 => "11111111",
	1976 => "11111111",
	1977 => "11111111",
	1978 => "11111111",
	1979 => "11111111",
	1984 => "11111111",
	1985 => "11111111",
	1986 => "11111111",
	1987 => "11111111",
	1988 => "11111111",
	1989 => "11111111",
	1990 => "11111111",
	1991 => "11111111",
	1992 => "11111111",
	1993 => "11111111",
	1994 => "11111111",
	1995 => "11111111",
	1996 => "11111111",
	1997 => "11111111",
	1998 => "11111111",
	1999 => "11111111",
	2000 => "11111111",
	2001 => "11111111",
	2002 => "11111111",
	2003 => "11111111",
	2004 => "11111111",
	2005 => "11111111",
	2006 => "11111111",
	2007 => "11111111",
	2008 => "11111111",
	2009 => "11111111",
	2010 => "11111111",
	2011 => "11111111",
	2012 => "11111111",
	2013 => "11111111",
	2014 => "11111111",
	2015 => "11111111",
	2016 => "11111111",
	2017 => "11111111",
	2018 => "11111111",
	2019 => "11111111",
	2020 => "11111111",
	2021 => "11111111",
	2022 => "11111111",
	2023 => "11111111",
	2024 => "11111111",
	2025 => "11111111",
	2026 => "11111111",
	2027 => "11111111",
	2028 => "11111111",
	2029 => "11111111",
	2030 => "11111111",
	2031 => "11111111",
	2032 => "11111111",
	2033 => "11111111",
	2034 => "11111111",
	2035 => "11111111",
	2036 => "11111111",
	2037 => "11111111",
	2038 => "11111111",
	2039 => "11111111",
	2040 => "11111111",
	2041 => "11111111",
	2042 => "11111111",
	2043 => "11111111",
	2048 => "11111111",
	2049 => "11111111",
	2050 => "11111111",
	2051 => "11111111",
	2052 => "11111111",
	2053 => "11111111",
	2054 => "11111111",
	2055 => "11111111",
	2056 => "11111111",
	2057 => "11111111",
	2058 => "11111111",
	2059 => "11111111",
	2060 => "11111111",
	2061 => "11111111",
	2062 => "11111111",
	2063 => "11111111",
	2064 => "11111111",
	2065 => "11111111",
	2066 => "11111111",
	2067 => "11111111",
	2068 => "11111111",
	2069 => "11111111",
	2070 => "11111111",
	2071 => "11111111",
	2072 => "11111111",
	2073 => "11111111",
	2074 => "11111111",
	2075 => "11111111",
	2076 => "11111111",
	2077 => "11111111",
	2078 => "11111111",
	2079 => "11111111",
	2080 => "11111111",
	2081 => "11111111",
	2082 => "11111111",
	2083 => "11111111",
	2084 => "11111111",
	2085 => "11111111",
	2086 => "11111111",
	2087 => "11111111",
	2088 => "11111111",
	2089 => "11111111",
	2090 => "11111111",
	2091 => "11111111",
	2092 => "11111111",
	2093 => "11111111",
	2094 => "11111111",
	2095 => "11111111",
	2096 => "11111111",
	2097 => "11111111",
	2098 => "11111111",
	2099 => "11111111",
	2100 => "11111111",
	2101 => "11111111",
	2102 => "11111111",
	2103 => "11111111",
	2104 => "11111111",
	2105 => "11111111",
	2106 => "11111111",
	2107 => "11111111",
	2112 => "11111111",
	2113 => "11111111",
	2114 => "11111111",
	2115 => "11111111",
	2116 => "11111111",
	2117 => "11111111",
	2118 => "11111111",
	2119 => "11111111",
	2120 => "11111111",
	2121 => "11111111",
	2122 => "11111111",
	2123 => "11111111",
	2124 => "11111111",
	2125 => "11111111",
	2126 => "11111111",
	2127 => "11111111",
	2128 => "11111111",
	2129 => "11111111",
	2130 => "11111111",
	2131 => "11111111",
	2132 => "11111111",
	2133 => "11111111",
	2134 => "11111111",
	2135 => "11111111",
	2136 => "11111111",
	2137 => "11111111",
	2138 => "11111111",
	2139 => "11111111",
	2140 => "11111111",
	2141 => "11111111",
	2142 => "11111111",
	2143 => "11111111",
	2144 => "11111111",
	2145 => "11111111",
	2146 => "11111111",
	2147 => "11111111",
	2148 => "11111111",
	2149 => "11111111",
	2150 => "11111111",
	2151 => "11111111",
	2152 => "11111111",
	2153 => "11111111",
	2154 => "11111111",
	2155 => "11111111",
	2156 => "11111111",
	2157 => "11111111",
	2158 => "11111111",
	2159 => "11111111",
	2160 => "11111111",
	2161 => "11111111",
	2162 => "11111111",
	2163 => "11111111",
	2164 => "11111111",
	2165 => "11111111",
	2166 => "11111111",
	2167 => "11111111",
	2168 => "11111111",
	2169 => "11111111",
	2170 => "11111111",
	2171 => "11111111",
	2176 => "11111111",
	2177 => "11111111",
	2178 => "11111111",
	2179 => "11111111",
	2180 => "11111111",
	2181 => "11111111",
	2182 => "11111111",
	2183 => "11111111",
	2184 => "11111111",
	2185 => "11111111",
	2186 => "11111111",
	2187 => "11111111",
	2188 => "11111111",
	2189 => "11111111",
	2190 => "11111111",
	2191 => "11111111",
	2192 => "11111111",
	2193 => "11111111",
	2194 => "11111111",
	2195 => "11111111",
	2196 => "11111111",
	2197 => "11111111",
	2198 => "11111111",
	2199 => "11111111",
	2200 => "11111111",
	2201 => "11111111",
	2202 => "11111111",
	2203 => "11111111",
	2204 => "11111111",
	2205 => "11111111",
	2206 => "11111111",
	2207 => "11111111",
	2208 => "11111111",
	2209 => "11111111",
	2210 => "11111111",
	2211 => "11111111",
	2212 => "11111111",
	2213 => "11111111",
	2214 => "11111111",
	2215 => "11111111",
	2216 => "11111111",
	2217 => "11111111",
	2218 => "11111111",
	2219 => "11111111",
	2220 => "11111111",
	2221 => "11111111",
	2222 => "11111111",
	2223 => "11111111",
	2224 => "11111111",
	2225 => "11111111",
	2226 => "11111111",
	2227 => "11111111",
	2228 => "11111111",
	2229 => "11111111",
	2230 => "11111111",
	2231 => "11111111",
	2232 => "11111111",
	2233 => "11111111",
	2234 => "11111111",
	2235 => "11111111",
	2240 => "11111111",
	2241 => "11111111",
	2242 => "11111111",
	2243 => "11111111",
	2244 => "11111111",
	2245 => "11111111",
	2246 => "11111111",
	2247 => "11111111",
	2248 => "11111111",
	2249 => "11111111",
	2250 => "11111111",
	2251 => "11111111",
	2252 => "11111111",
	2253 => "11111111",
	2254 => "11111111",
	2255 => "11111111",
	2256 => "11111111",
	2257 => "11111111",
	2258 => "11111111",
	2259 => "11111111",
	2260 => "11111111",
	2261 => "11111111",
	2262 => "11111111",
	2263 => "11111111",
	2264 => "11111111",
	2265 => "11111111",
	2266 => "11111111",
	2267 => "11111111",
	2268 => "11111111",
	2269 => "11111111",
	2270 => "11111111",
	2271 => "11111111",
	2272 => "11111111",
	2273 => "11111111",
	2274 => "11111111",
	2275 => "11111111",
	2276 => "11111111",
	2277 => "11111111",
	2278 => "11111111",
	2279 => "11111111",
	2280 => "11111111",
	2281 => "11111111",
	2282 => "11111111",
	2283 => "11111111",
	2284 => "11111111",
	2285 => "11111111",
	2286 => "11111111",
	2287 => "11111111",
	2288 => "11111111",
	2289 => "11111111",
	2290 => "11111111",
	2291 => "11111111",
	2292 => "11111111",
	2293 => "11111111",
	2294 => "11111111",
	2295 => "11111111",
	2296 => "11111111",
	2297 => "11111111",
	2298 => "11111111",
	2299 => "11111111",
	2304 => "11111111",
	2305 => "11111111",
	2306 => "11111111",
	2307 => "11111111",
	2308 => "11111111",
	2309 => "11111111",
	2310 => "11111111",
	2311 => "11111111",
	2312 => "11111111",
	2313 => "11111111",
	2314 => "11111111",
	2315 => "11111111",
	2316 => "11111111",
	2317 => "11111111",
	2318 => "11111111",
	2319 => "11111111",
	2320 => "11111111",
	2321 => "11111111",
	2322 => "11111111",
	2323 => "11111111",
	2324 => "11111111",
	2325 => "11111111",
	2326 => "11111111",
	2327 => "11111111",
	2328 => "11111111",
	2329 => "11111111",
	2330 => "11111111",
	2331 => "11111111",
	2332 => "11111111",
	2333 => "11111111",
	2334 => "11111111",
	2335 => "11111111",
	2336 => "11111111",
	2337 => "11111111",
	2338 => "11111111",
	2339 => "11111111",
	2340 => "11111111",
	2341 => "11111111",
	2342 => "11111111",
	2343 => "11111111",
	2344 => "11111111",
	2345 => "11111111",
	2346 => "11111111",
	2347 => "11111111",
	2348 => "11111111",
	2349 => "11111111",
	2350 => "11111111",
	2351 => "11111111",
	2352 => "11111111",
	2353 => "11111111",
	2354 => "11111111",
	2355 => "11111111",
	2356 => "11111111",
	2357 => "11111111",
	2358 => "11111111",
	2359 => "11111111",
	2360 => "11111111",
	2361 => "11111111",
	2362 => "11111111",
	2363 => "11111111",
	2368 => "11111111",
	2369 => "11111111",
	2370 => "11111111",
	2371 => "11111111",
	2372 => "11111111",
	2373 => "11111111",
	2374 => "11111111",
	2375 => "11111111",
	2376 => "11111111",
	2377 => "11111111",
	2378 => "11111111",
	2379 => "11111111",
	2380 => "11111111",
	2381 => "11111111",
	2382 => "11111111",
	2383 => "11111111",
	2384 => "11111111",
	2385 => "11111111",
	2386 => "11111111",
	2387 => "11111111",
	2388 => "11111111",
	2389 => "11111111",
	2390 => "11111111",
	2391 => "11111111",
	2392 => "11111111",
	2393 => "11111111",
	2394 => "11111111",
	2395 => "11111111",
	2396 => "11111111",
	2397 => "11111111",
	2398 => "11111111",
	2399 => "11111111",
	2400 => "11111111",
	2401 => "11111111",
	2402 => "11111111",
	2403 => "11111111",
	2404 => "11111111",
	2405 => "11111111",
	2406 => "11111111",
	2407 => "11111111",
	2408 => "11111111",
	2409 => "11111111",
	2410 => "11111111",
	2411 => "11111111",
	2412 => "11111111",
	2413 => "11111111",
	2414 => "11111111",
	2415 => "11111111",
	2416 => "11111111",
	2417 => "11111111",
	2418 => "11111111",
	2419 => "11111111",
	2420 => "11111111",
	2421 => "11111111",
	2422 => "11111111",
	2423 => "11111111",
	2424 => "11111111",
	2425 => "11111111",
	2426 => "11111111",
	2427 => "11111111",
	2432 => "11111111",
	2433 => "11111111",
	2434 => "11111111",
	2435 => "11111111",
	2436 => "11111111",
	2437 => "11111111",
	2438 => "11111111",
	2439 => "11111111",
	2440 => "11111111",
	2441 => "11111111",
	2442 => "11111111",
	2443 => "11111111",
	2444 => "11111111",
	2445 => "11111111",
	2446 => "11111111",
	2447 => "11111111",
	2448 => "11111111",
	2449 => "11111111",
	2450 => "11111111",
	2451 => "11111111",
	2452 => "11111111",
	2453 => "11111111",
	2454 => "11111111",
	2455 => "11111111",
	2456 => "11111111",
	2457 => "11111111",
	2458 => "11111111",
	2459 => "11111111",
	2460 => "11111111",
	2461 => "11111111",
	2462 => "11111111",
	2463 => "11111111",
	2464 => "11111111",
	2465 => "11111111",
	2466 => "11111111",
	2467 => "11111111",
	2468 => "11111111",
	2469 => "11111111",
	2470 => "11111111",
	2471 => "11111111",
	2472 => "11111111",
	2473 => "11111111",
	2474 => "11111111",
	2475 => "11111111",
	2476 => "11111111",
	2477 => "11111111",
	2478 => "11111111",
	2479 => "11111111",
	2480 => "11111111",
	2481 => "11111111",
	2482 => "11111111",
	2483 => "11111111",
	2484 => "11111111",
	2485 => "11111111",
	2486 => "11111111",
	2487 => "11111111",
	2488 => "11111111",
	2489 => "11111111",
	2490 => "11111111",
	2491 => "11111111",
	2496 => "11111111",
	2497 => "11111111",
	2498 => "11111111",
	2499 => "11111111",
	2500 => "11111111",
	2501 => "11111111",
	2502 => "11111111",
	2503 => "11111111",
	2504 => "11111111",
	2505 => "11111111",
	2506 => "11111111",
	2507 => "11111111",
	2508 => "11111111",
	2509 => "11111111",
	2510 => "11111111",
	2511 => "11111111",
	2512 => "11111111",
	2513 => "11111111",
	2514 => "11111111",
	2515 => "11111111",
	2516 => "11111111",
	2517 => "11111111",
	2518 => "11111111",
	2519 => "11111111",
	2520 => "11111111",
	2521 => "11111111",
	2522 => "11111111",
	2523 => "11111111",
	2524 => "11111111",
	2525 => "11111111",
	2526 => "11111111",
	2527 => "11111111",
	2528 => "11111111",
	2529 => "11111111",
	2530 => "11111111",
	2531 => "11111111",
	2532 => "11111111",
	2533 => "11111111",
	2534 => "11111111",
	2535 => "11111111",
	2536 => "11111111",
	2537 => "11111111",
	2538 => "11111111",
	2539 => "11111111",
	2540 => "11111111",
	2541 => "11111111",
	2542 => "11111111",
	2543 => "11111111",
	2544 => "11111111",
	2545 => "11111111",
	2546 => "11111111",
	2547 => "11111111",
	2548 => "11111111",
	2549 => "11111111",
	2550 => "11111111",
	2551 => "11111111",
	2552 => "11111111",
	2553 => "11111111",
	2554 => "11111111",
	2555 => "11111111",
	2560 => "11111111",
	2561 => "11111111",
	2562 => "11111111",
	2563 => "11111111",
	2564 => "11111111",
	2565 => "11111111",
	2566 => "11111111",
	2567 => "11111111",
	2568 => "11111111",
	2569 => "11111111",
	2570 => "11111111",
	2571 => "11111111",
	2572 => "11111111",
	2573 => "11111111",
	2574 => "11111111",
	2575 => "11111111",
	2576 => "11111111",
	2577 => "11111111",
	2578 => "11111111",
	2579 => "11111111",
	2580 => "11111111",
	2581 => "11111111",
	2582 => "11111111",
	2583 => "11111111",
	2584 => "11111111",
	2585 => "11111111",
	2586 => "11111111",
	2587 => "11111111",
	2588 => "11111111",
	2589 => "11111111",
	2590 => "11111111",
	2591 => "11111111",
	2592 => "11111111",
	2593 => "11111111",
	2594 => "11111111",
	2595 => "11111111",
	2596 => "11111111",
	2597 => "11111111",
	2598 => "11111111",
	2599 => "11111111",
	2600 => "11111111",
	2601 => "11111111",
	2602 => "11111111",
	2603 => "11111111",
	2604 => "11111111",
	2605 => "11111111",
	2606 => "11111111",
	2607 => "11111111",
	2608 => "11111111",
	2609 => "11111111",
	2610 => "11111111",
	2611 => "11111111",
	2612 => "11111111",
	2613 => "11111111",
	2614 => "11111111",
	2615 => "11111111",
	2616 => "11111111",
	2617 => "11111111",
	2618 => "11111111",
	2619 => "11111111",
	2624 => "11111111",
	2625 => "11111111",
	2626 => "11111111",
	2627 => "11111111",
	2628 => "11111111",
	2629 => "11111111",
	2630 => "11111111",
	2631 => "11111111",
	2632 => "11111111",
	2633 => "11111111",
	2634 => "11111111",
	2635 => "11111111",
	2636 => "11111111",
	2637 => "11111111",
	2638 => "11111111",
	2639 => "11111111",
	2640 => "11111111",
	2641 => "11111111",
	2642 => "11111111",
	2643 => "11111111",
	2644 => "11111111",
	2645 => "11111111",
	2646 => "11111111",
	2647 => "11111111",
	2648 => "11111111",
	2649 => "11111111",
	2650 => "11111111",
	2651 => "11111111",
	2652 => "11111111",
	2653 => "11111111",
	2654 => "11111111",
	2655 => "11111111",
	2656 => "11111111",
	2657 => "11111111",
	2658 => "11111111",
	2659 => "11111111",
	2660 => "11111111",
	2661 => "11111111",
	2662 => "11111111",
	2663 => "11111111",
	2664 => "11111111",
	2665 => "11111111",
	2666 => "11111111",
	2667 => "11111111",
	2668 => "11111111",
	2669 => "11111111",
	2670 => "11111111",
	2671 => "11111111",
	2672 => "11111111",
	2673 => "11111111",
	2674 => "11111111",
	2675 => "11111111",
	2676 => "11111111",
	2677 => "11111111",
	2678 => "11111111",
	2679 => "11111111",
	2680 => "11111111",
	2681 => "11111111",
	2682 => "11111111",
	2683 => "11111111",
	2688 => "11111111",
	2689 => "11111111",
	2690 => "11111111",
	2691 => "11111111",
	2692 => "11111111",
	2693 => "11111111",
	2694 => "11111111",
	2695 => "11111111",
	2696 => "11111111",
	2697 => "11111111",
	2698 => "11111111",
	2699 => "11111111",
	2700 => "11111111",
	2701 => "11111111",
	2702 => "11111111",
	2703 => "11111111",
	2704 => "11111111",
	2705 => "11111111",
	2706 => "11111111",
	2707 => "11111111",
	2708 => "11111111",
	2709 => "11111111",
	2710 => "11111111",
	2711 => "11111111",
	2712 => "11111111",
	2713 => "11111111",
	2714 => "11111111",
	2715 => "11111111",
	2716 => "11111111",
	2717 => "11111111",
	2718 => "11111111",
	2719 => "11111111",
	2720 => "11111111",
	2721 => "11111111",
	2722 => "11111111",
	2723 => "11111111",
	2724 => "11111111",
	2725 => "11111111",
	2726 => "11111111",
	2727 => "11111111",
	2728 => "11111111",
	2729 => "11111111",
	2730 => "11111111",
	2731 => "11111111",
	2732 => "11111111",
	2733 => "11111111",
	2734 => "11111111",
	2735 => "11111111",
	2736 => "11111111",
	2737 => "11111111",
	2738 => "11111111",
	2739 => "11111111",
	2740 => "11111111",
	2741 => "11111111",
	2742 => "11111111",
	2743 => "11111111",
	2744 => "11111111",
	2745 => "11111111",
	2746 => "11111111",
	2747 => "11111111",
	2752 => "11111111",
	2753 => "11111111",
	2754 => "11111111",
	2755 => "11111111",
	2756 => "11111111",
	2757 => "11111111",
	2758 => "11111111",
	2759 => "11111111",
	2760 => "11111111",
	2761 => "11111111",
	2762 => "11111111",
	2763 => "11111111",
	2764 => "11111111",
	2765 => "11111111",
	2766 => "11111111",
	2767 => "11111111",
	2768 => "11111111",
	2769 => "11111111",
	2770 => "11111111",
	2771 => "11111111",
	2772 => "11111111",
	2773 => "11111111",
	2774 => "11111111",
	2775 => "11111111",
	2776 => "11111111",
	2777 => "11111111",
	2778 => "11111111",
	2779 => "11111111",
	2780 => "11111111",
	2781 => "11111111",
	2782 => "11111111",
	2783 => "11111111",
	2784 => "11111111",
	2785 => "11111111",
	2786 => "11111111",
	2787 => "11111111",
	2788 => "11111111",
	2789 => "11111111",
	2790 => "11111111",
	2791 => "11111111",
	2792 => "11111111",
	2793 => "11111111",
	2794 => "11111111",
	2795 => "11111111",
	2796 => "11111111",
	2797 => "11111111",
	2798 => "11111111",
	2799 => "11111111",
	2800 => "11111111",
	2801 => "11111111",
	2802 => "11111111",
	2803 => "11111111",
	2804 => "11111111",
	2805 => "11111111",
	2806 => "11111111",
	2807 => "11111111",
	2808 => "11111111",
	2809 => "11111111",
	2810 => "11111111",
	2811 => "11111111",
	2816 => "11111111",
	2817 => "11111111",
	2818 => "11111111",
	2819 => "11111111",
	2820 => "11111111",
	2821 => "11111111",
	2822 => "11111111",
	2823 => "11111111",
	2824 => "11111111",
	2825 => "11111111",
	2826 => "11111111",
	2827 => "11111111",
	2828 => "11111111",
	2829 => "11111111",
	2830 => "11111111",
	2831 => "11111111",
	2832 => "11111111",
	2833 => "11111111",
	2834 => "11111111",
	2835 => "11111111",
	2836 => "11111111",
	2837 => "11111111",
	2838 => "11111111",
	2839 => "11111111",
	2840 => "11111111",
	2841 => "11111111",
	2842 => "11111111",
	2843 => "11111111",
	2844 => "11111111",
	2845 => "11111111",
	2846 => "11111111",
	2847 => "11111111",
	2848 => "11111111",
	2849 => "11111111",
	2850 => "11111111",
	2851 => "11111111",
	2852 => "11111111",
	2853 => "11111111",
	2854 => "11111111",
	2855 => "11111111",
	2856 => "11111111",
	2857 => "11111111",
	2858 => "11111111",
	2859 => "11111111",
	2860 => "11111111",
	2861 => "11111111",
	2862 => "11111111",
	2863 => "11111111",
	2864 => "11111111",
	2865 => "11111111",
	2866 => "11111111",
	2867 => "11111111",
	2868 => "11111111",
	2869 => "11111111",
	2870 => "11111111",
	2871 => "11111111",
	2872 => "11111111",
	2873 => "11111111",
	2874 => "11111111",
	2875 => "11111111",
	2880 => "11111111",
	2881 => "11111111",
	2882 => "11111111",
	2883 => "11111111",
	2884 => "11111111",
	2885 => "11111111",
	2886 => "11111111",
	2887 => "11111111",
	2888 => "11111111",
	2889 => "11111111",
	2890 => "11111111",
	2891 => "11111111",
	2892 => "11111111",
	2893 => "11111111",
	2894 => "11111111",
	2895 => "11111111",
	2896 => "11111111",
	2897 => "11111111",
	2898 => "11111111",
	2899 => "11111111",
	2900 => "11111111",
	2901 => "11111111",
	2902 => "11111111",
	2903 => "11111111",
	2904 => "11111111",
	2905 => "11111111",
	2906 => "11111111",
	2907 => "11111111",
	2908 => "11111111",
	2909 => "11111111",
	2910 => "11111111",
	2911 => "11111111",
	2912 => "11111111",
	2913 => "11111111",
	2914 => "11111111",
	2915 => "11111111",
	2916 => "11111111",
	2917 => "11111111",
	2918 => "11111111",
	2919 => "11111111",
	2920 => "11111111",
	2921 => "11111111",
	2922 => "11111111",
	2923 => "11111111",
	2924 => "11111111",
	2925 => "11111111",
	2926 => "11111111",
	2927 => "11111111",
	2928 => "11111111",
	2929 => "11111111",
	2930 => "11111111",
	2931 => "11111111",
	2932 => "11111111",
	2933 => "11111111",
	2934 => "11111111",
	2935 => "11111111",
	2936 => "11111111",
	2937 => "11111111",
	2938 => "11111111",
	2939 => "11111111",
	2944 => "11111111",
	2945 => "11111111",
	2946 => "11111111",
	2947 => "11111111",
	2948 => "11111111",
	2949 => "11111111",
	2950 => "11111111",
	2951 => "11111111",
	2952 => "11111111",
	2953 => "11111111",
	2954 => "11111111",
	2955 => "11111111",
	2956 => "11111111",
	2957 => "11111111",
	2958 => "11111111",
	2959 => "11111111",
	2960 => "11111111",
	2961 => "11111111",
	2962 => "11111111",
	2963 => "11111111",
	2964 => "11111111",
	2965 => "11111111",
	2966 => "11111111",
	2967 => "11111111",
	2968 => "11111111",
	2969 => "11111111",
	2970 => "11111111",
	2971 => "11111111",
	2972 => "11111111",
	2973 => "11111111",
	2974 => "11111111",
	2975 => "11111111",
	2976 => "11111111",
	2977 => "11111111",
	2978 => "11111111",
	2979 => "11111111",
	2980 => "11111111",
	2981 => "11111111",
	2982 => "11111111",
	2983 => "11111111",
	2984 => "11111111",
	2985 => "11111111",
	2986 => "11111111",
	2987 => "11111111",
	2988 => "11111111",
	2989 => "11111111",
	2990 => "11111111",
	2991 => "11111111",
	2992 => "11111111",
	2993 => "11111111",
	2994 => "11111111",
	2995 => "11111111",
	2996 => "11111111",
	2997 => "11111111",
	2998 => "11111111",
	2999 => "11111111",
	3000 => "11111111",
	3001 => "11111111",
	3002 => "11111111",
	3003 => "11111111",
	3008 => "11111111",
	3009 => "11111111",
	3010 => "11111111",
	3011 => "11111111",
	3012 => "11111111",
	3013 => "11111111",
	3014 => "11111111",
	3015 => "11111111",
	3016 => "11111111",
	3017 => "11111111",
	3018 => "11111111",
	3019 => "11111111",
	3020 => "11111111",
	3021 => "11111111",
	3022 => "11111111",
	3023 => "11111111",
	3024 => "11111111",
	3025 => "11111111",
	3026 => "11111111",
	3027 => "11111111",
	3028 => "11111111",
	3029 => "11111111",
	3030 => "11111111",
	3031 => "11111111",
	3032 => "11111111",
	3033 => "11111111",
	3034 => "11111111",
	3035 => "11111111",
	3036 => "11111111",
	3037 => "11111111",
	3038 => "11111111",
	3039 => "11111111",
	3040 => "11111111",
	3041 => "11111111",
	3042 => "11111111",
	3043 => "11111111",
	3044 => "11111111",
	3045 => "11111111",
	3046 => "11111111",
	3047 => "11111111",
	3048 => "11111111",
	3049 => "11111111",
	3050 => "11111111",
	3051 => "11111111",
	3052 => "11111111",
	3053 => "11111111",
	3054 => "11111111",
	3055 => "11111111",
	3056 => "11111111",
	3057 => "11111111",
	3058 => "11111111",
	3059 => "11111111",
	3060 => "11111111",
	3061 => "11111111",
	3062 => "11111111",
	3063 => "11111111",
	3064 => "11111111",
	3065 => "11111111",
	3066 => "11111111",
	3067 => "11111111",
	3072 => "11111111",
	3073 => "11111111",
	3074 => "11111111",
	3075 => "11111111",
	3076 => "11111111",
	3077 => "11111111",
	3078 => "11111111",
	3079 => "11111111",
	3080 => "11111111",
	3081 => "11111111",
	3082 => "11111111",
	3083 => "11111111",
	3084 => "11111111",
	3085 => "11111111",
	3086 => "11111111",
	3087 => "11111111",
	3088 => "11111111",
	3089 => "11111111",
	3090 => "11111111",
	3091 => "11111111",
	3092 => "11111111",
	3093 => "11111111",
	3094 => "11111111",
	3095 => "11111111",
	3096 => "11111111",
	3097 => "11111111",
	3098 => "11111111",
	3099 => "11111111",
	3100 => "11111111",
	3101 => "11111111",
	3102 => "11111111",
	3103 => "11111111",
	3104 => "11111111",
	3105 => "11111111",
	3106 => "11111111",
	3107 => "11111111",
	3108 => "11111111",
	3109 => "11111111",
	3110 => "11111111",
	3111 => "11111111",
	3112 => "11111111",
	3113 => "11111111",
	3114 => "11111111",
	3115 => "11111111",
	3116 => "11111111",
	3117 => "11111111",
	3118 => "11111111",
	3119 => "11111111",
	3120 => "11111111",
	3121 => "11111111",
	3122 => "11111111",
	3123 => "11111111",
	3124 => "11111111",
	3125 => "11111111",
	3126 => "11111111",
	3127 => "11111111",
	3128 => "11111111",
	3129 => "11111111",
	3130 => "11111111",
	3131 => "11111111",
	3136 => "11111111",
	3137 => "11111111",
	3138 => "11111111",
	3139 => "11111111",
	3140 => "11111111",
	3141 => "11111111",
	3142 => "11111111",
	3143 => "11111111",
	3144 => "11111111",
	3145 => "11111111",
	3146 => "11111111",
	3147 => "11111111",
	3148 => "11111111",
	3149 => "11111111",
	3150 => "11111111",
	3151 => "11111111",
	3152 => "11111111",
	3153 => "11111111",
	3154 => "11111111",
	3155 => "11111111",
	3156 => "11111111",
	3157 => "11111111",
	3158 => "11111111",
	3159 => "11111111",
	3160 => "11111111",
	3161 => "11111111",
	3162 => "11111111",
	3163 => "11111111",
	3164 => "11111111",
	3165 => "11111111",
	3166 => "11111111",
	3167 => "11111111",
	3168 => "11111111",
	3169 => "11111111",
	3170 => "11111111",
	3171 => "11111111",
	3172 => "11111111",
	3173 => "11111111",
	3174 => "11111111",
	3175 => "11111111",
	3176 => "11111111",
	3177 => "11111111",
	3178 => "11111111",
	3179 => "11111111",
	3180 => "11111111",
	3181 => "11111111",
	3182 => "11111111",
	3183 => "11111111",
	3184 => "11111111",
	3185 => "11111111",
	3186 => "11111111",
	3187 => "11111111",
	3188 => "11111111",
	3189 => "11111111",
	3190 => "11111111",
	3191 => "11111111",
	3192 => "11111111",
	3193 => "11111111",
	3194 => "11111111",
	3195 => "11111111",
	3200 => "11111111",
	3201 => "11111111",
	3202 => "11111111",
	3203 => "11111111",
	3204 => "11111111",
	3205 => "11111111",
	3206 => "11111111",
	3207 => "11111111",
	3208 => "11111111",
	3209 => "11111111",
	3210 => "11111111",
	3211 => "11111111",
	3212 => "11111111",
	3213 => "11111111",
	3214 => "11111111",
	3215 => "11111111",
	3216 => "11111111",
	3217 => "11111111",
	3218 => "11111111",
	3219 => "11111111",
	3220 => "11111111",
	3221 => "11111111",
	3222 => "11111111",
	3223 => "11111111",
	3224 => "11111111",
	3225 => "11111111",
	3226 => "11111111",
	3227 => "11111111",
	3228 => "11111111",
	3229 => "11111111",
	3230 => "11111111",
	3231 => "11111111",
	3232 => "11111111",
	3233 => "11111111",
	3234 => "11111111",
	3235 => "11111111",
	3236 => "11111111",
	3237 => "11111111",
	3238 => "11111111",
	3239 => "11111111",
	3240 => "11111111",
	3241 => "11111111",
	3242 => "11111111",
	3243 => "11111111",
	3244 => "11111111",
	3245 => "11111111",
	3246 => "11111111",
	3247 => "11111111",
	3248 => "11111111",
	3249 => "11111111",
	3250 => "11111111",
	3251 => "11111111",
	3252 => "11111111",
	3253 => "11111111",
	3254 => "11111111",
	3255 => "11111111",
	3256 => "11111111",
	3257 => "11111111",
	3258 => "11111111",
	3259 => "11111111",
	3264 => "11111111",
	3265 => "11111111",
	3266 => "11111111",
	3267 => "11111111",
	3268 => "11111111",
	3269 => "11111111",
	3270 => "11111111",
	3271 => "11111111",
	3272 => "11111111",
	3273 => "11111111",
	3274 => "11111111",
	3275 => "11111111",
	3276 => "11111111",
	3277 => "11111111",
	3278 => "11111111",
	3279 => "11111111",
	3280 => "11111111",
	3281 => "11111111",
	3282 => "11111111",
	3283 => "11111111",
	3284 => "11111111",
	3285 => "11111111",
	3286 => "11111111",
	3287 => "11111111",
	3288 => "11111111",
	3289 => "11111111",
	3290 => "11111111",
	3291 => "11111111",
	3292 => "11111111",
	3293 => "11111111",
	3294 => "11111111",
	3295 => "11111111",
	3296 => "11111111",
	3297 => "11111111",
	3298 => "11111111",
	3299 => "11111111",
	3300 => "11111111",
	3301 => "11111111",
	3302 => "11111111",
	3303 => "11111111",
	3304 => "11111111",
	3305 => "11111111",
	3306 => "11111111",
	3307 => "11111111",
	3308 => "11111111",
	3309 => "11111111",
	3310 => "11111111",
	3311 => "11111111",
	3312 => "11111111",
	3313 => "11111111",
	3314 => "11111111",
	3315 => "11111111",
	3316 => "11111111",
	3317 => "11111111",
	3318 => "11111111",
	3319 => "11111111",
	3320 => "11111111",
	3321 => "11111111",
	3322 => "11111111",
	3323 => "11111111",
	3328 => "11111111",
	3329 => "11111111",
	3330 => "11111111",
	3331 => "11111111",
	3332 => "11111111",
	3333 => "11111111",
	3334 => "11111111",
	3335 => "11111111",
	3336 => "11111111",
	3337 => "11111111",
	3338 => "11111111",
	3339 => "11111111",
	3340 => "11111111",
	3341 => "11111111",
	3342 => "11111111",
	3343 => "11111111",
	3344 => "11111111",
	3345 => "11111111",
	3346 => "11111111",
	3347 => "11111111",
	3348 => "11111111",
	3349 => "11111111",
	3350 => "11111111",
	3351 => "11111111",
	3352 => "11111111",
	3353 => "11111111",
	3354 => "11111111",
	3355 => "11111111",
	3356 => "11111111",
	3357 => "11111111",
	3358 => "11111111",
	3359 => "11111111",
	3360 => "11111111",
	3361 => "11111111",
	3362 => "11111111",
	3363 => "11111111",
	3364 => "11111111",
	3365 => "11111111",
	3366 => "11111111",
	3367 => "11111111",
	3368 => "11111111",
	3369 => "11111111",
	3370 => "11111111",
	3371 => "11111111",
	3372 => "11111111",
	3373 => "11111111",
	3374 => "11111111",
	3375 => "11111111",
	3376 => "11111111",
	3377 => "11111111",
	3378 => "11111111",
	3379 => "11111111",
	3380 => "11111111",
	3381 => "11111111",
	3382 => "11111111",
	3383 => "11111111",
	3384 => "11111111",
	3385 => "11111111",
	3386 => "11111111",
	3387 => "11111111",
	3392 => "11111111",
	3393 => "11111111",
	3394 => "11111111",
	3395 => "11111111",
	3396 => "11111111",
	3397 => "11111111",
	3398 => "11111111",
	3399 => "11111111",
	3400 => "11111111",
	3401 => "11111111",
	3402 => "11111111",
	3403 => "11111111",
	3404 => "11111111",
	3405 => "11111111",
	3406 => "11111111",
	3407 => "11111111",
	3408 => "11111111",
	3409 => "11111111",
	3410 => "11111111",
	3411 => "11111111",
	3412 => "11111111",
	3413 => "11111111",
	3414 => "11111111",
	3415 => "11111111",
	3416 => "11111111",
	3417 => "11111111",
	3418 => "11111111",
	3419 => "11111111",
	3420 => "11111111",
	3421 => "11111111",
	3422 => "11111111",
	3423 => "11111111",
	3424 => "11111111",
	3425 => "11111111",
	3426 => "11111111",
	3427 => "11111111",
	3428 => "11111111",
	3429 => "11111111",
	3430 => "11111111",
	3431 => "11111111",
	3432 => "11111111",
	3433 => "11111111",
	3434 => "11111111",
	3435 => "11111111",
	3436 => "11111111",
	3437 => "11111111",
	3438 => "11111111",
	3439 => "11111111",
	3440 => "11111111",
	3441 => "11111111",
	3442 => "11111111",
	3443 => "11111111",
	3444 => "11111111",
	3445 => "11111111",
	3446 => "11111111",
	3447 => "11111111",
	3448 => "11111111",
	3449 => "11111111",
	3450 => "11111111",
	3451 => "11111111",
	3456 => "11111111",
	3457 => "11111111",
	3458 => "11111111",
	3459 => "11111111",
	3460 => "11111111",
	3461 => "11111111",
	3462 => "11111111",
	3463 => "11111111",
	3464 => "11111111",
	3465 => "11111111",
	3466 => "11111111",
	3467 => "11111111",
	3468 => "11111111",
	3469 => "11111111",
	3470 => "11111111",
	3471 => "11111111",
	3472 => "11111111",
	3473 => "11111111",
	3474 => "11111111",
	3475 => "11111111",
	3476 => "11111111",
	3477 => "11111111",
	3478 => "11111111",
	3479 => "11111111",
	3480 => "11111111",
	3481 => "11111111",
	3482 => "11111111",
	3483 => "11111111",
	3484 => "11111111",
	3485 => "11111111",
	3486 => "11111111",
	3487 => "11111111",
	3488 => "11111111",
	3489 => "11111111",
	3490 => "11111111",
	3491 => "11111111",
	3492 => "11111111",
	3493 => "11111111",
	3494 => "11111111",
	3495 => "11111111",
	3496 => "11111111",
	3497 => "11111111",
	3498 => "11111111",
	3499 => "11111111",
	3500 => "11111111",
	3501 => "11111111",
	3502 => "11111111",
	3503 => "11111111",
	3504 => "11111111",
	3505 => "11111111",
	3506 => "11111111",
	3507 => "11111111",
	3508 => "11111111",
	3509 => "11111111",
	3510 => "11111111",
	3511 => "11111111",
	3512 => "11111111",
	3513 => "11111111",
	3514 => "11111111",
	3515 => "11111111",
	3520 => "11111111",
	3521 => "11111111",
	3522 => "11111111",
	3523 => "11111111",
	3524 => "11111111",
	3525 => "11111111",
	3526 => "11111111",
	3527 => "11111111",
	3528 => "11111111",
	3529 => "11111111",
	3530 => "11111111",
	3531 => "11111111",
	3532 => "11111111",
	3533 => "11111111",
	3534 => "11111111",
	3535 => "11111111",
	3536 => "11111111",
	3537 => "11111111",
	3538 => "11111111",
	3539 => "11111111",
	3540 => "11111111",
	3541 => "11111111",
	3542 => "11111111",
	3543 => "11111111",
	3544 => "11111111",
	3545 => "11111111",
	3546 => "11111111",
	3547 => "11111111",
	3548 => "11111111",
	3549 => "11111111",
	3550 => "11111111",
	3551 => "11111111",
	3552 => "11111111",
	3553 => "11111111",
	3554 => "11111111",
	3555 => "11111111",
	3556 => "11111111",
	3557 => "11111111",
	3558 => "11111111",
	3559 => "11111111",
	3560 => "11111111",
	3561 => "11111111",
	3562 => "11111111",
	3563 => "11111111",
	3564 => "11111111",
	3565 => "11111111",
	3566 => "11111111",
	3567 => "11111111",
	3568 => "11111111",
	3569 => "11111111",
	3570 => "11111111",
	3571 => "11111111",
	3572 => "11111111",
	3573 => "11111111",
	3574 => "11111111",
	3575 => "11111111",
	3576 => "11111111",
	3577 => "11111111",
	3578 => "11111111",
	3579 => "11111111",
	3584 => "11111111",
	3585 => "11111111",
	3586 => "11111111",
	3587 => "11111111",
	3588 => "11111111",
	3589 => "11111111",
	3590 => "11111111",
	3591 => "11111111",
	3592 => "11111111",
	3593 => "11111111",
	3594 => "11111111",
	3595 => "11111111",
	3596 => "11111111",
	3597 => "11111111",
	3598 => "11111111",
	3599 => "11111111",
	3600 => "11111111",
	3601 => "11111111",
	3602 => "11111111",
	3603 => "11111111",
	3604 => "11111111",
	3605 => "11111111",
	3606 => "11111111",
	3607 => "11111111",
	3608 => "11111111",
	3609 => "11111111",
	3610 => "11111111",
	3611 => "11111111",
	3612 => "11111111",
	3613 => "11111111",
	3614 => "11111111",
	3615 => "11111111",
	3616 => "11111111",
	3617 => "11111111",
	3618 => "11111111",
	3619 => "11111111",
	3620 => "11111111",
	3621 => "11111111",
	3622 => "11111111",
	3623 => "11111111",
	3624 => "11111111",
	3625 => "11111111",
	3626 => "11111111",
	3627 => "11111111",
	3628 => "11111111",
	3629 => "11111111",
	3630 => "11111111",
	3631 => "11111111",
	3632 => "11111111",
	3633 => "11111111",
	3634 => "11111111",
	3635 => "11111111",
	3636 => "11111111",
	3637 => "11111111",
	3638 => "11111111",
	3639 => "11111111",
	3640 => "11111111",
	3641 => "11111111",
	3642 => "11111111",
	3643 => "11111111",
	3648 => "11111111",
	3649 => "11111111",
	3650 => "11111111",
	3651 => "11111111",
	3652 => "11111111",
	3653 => "11111111",
	3654 => "11111111",
	3655 => "11111111",
	3656 => "11111111",
	3657 => "11111111",
	3658 => "11111111",
	3659 => "11111111",
	3660 => "11111111",
	3661 => "11111111",
	3662 => "11111111",
	3663 => "11111111",
	3664 => "11111111",
	3665 => "11111111",
	3666 => "11111111",
	3667 => "11111111",
	3668 => "11111111",
	3669 => "11111111",
	3670 => "11111111",
	3671 => "11111111",
	3672 => "11111111",
	3673 => "11111111",
	3674 => "11111111",
	3675 => "11111111",
	3676 => "11111111",
	3677 => "11111111",
	3678 => "11111111",
	3679 => "11111111",
	3680 => "11111111",
	3681 => "11111111",
	3682 => "11111111",
	3683 => "11111111",
	3684 => "11111111",
	3685 => "11111111",
	3686 => "11111111",
	3687 => "11111111",
	3688 => "11111111",
	3689 => "11111111",
	3690 => "11111111",
	3691 => "11111111",
	3692 => "11111111",
	3693 => "11111111",
	3694 => "11111111",
	3695 => "11111111",
	3696 => "11111111",
	3697 => "11111111",
	3698 => "11111111",
	3699 => "11111111",
	3700 => "11111111",
	3701 => "11111111",
	3702 => "11111111",
	3703 => "11111111",
	3704 => "11111111",
	3705 => "11111111",
	3706 => "11111111",
	3707 => "11111111",
	3712 => "11111111",
	3713 => "11111111",
	3714 => "11111111",
	3715 => "11111111",
	3716 => "11111111",
	3717 => "11111111",
	3718 => "11111111",
	3719 => "11111111",
	3720 => "11111111",
	3721 => "11111111",
	3722 => "11111111",
	3723 => "11111111",
	3724 => "11111111",
	3725 => "11111111",
	3726 => "11111111",
	3727 => "11111111",
	3728 => "11111111",
	3729 => "11111111",
	3730 => "11111111",
	3731 => "11111111",
	3732 => "11111111",
	3733 => "11111111",
	3734 => "11111111",
	3735 => "11111111",
	3736 => "11111111",
	3737 => "11111111",
	3738 => "11111111",
	3739 => "11111111",
	3740 => "11111111",
	3741 => "11111111",
	3742 => "11111111",
	3743 => "11111111",
	3744 => "11111111",
	3745 => "11111111",
	3746 => "11111111",
	3747 => "11111111",
	3748 => "11111111",
	3749 => "11111111",
	3750 => "11111111",
	3751 => "11111111",
	3752 => "11111111",
	3753 => "11111111",
	3754 => "11111111",
	3755 => "11111111",
	3756 => "11111111",
	3757 => "11111111",
	3758 => "11111111",
	3759 => "11111111",
	3760 => "11111111",
	3761 => "11111111",
	3762 => "11111111",
	3763 => "11111111",
	3764 => "11111111",
	3765 => "11111111",
	3766 => "11111111",
	3767 => "11111111",
	3768 => "11111111",
	3769 => "11111111",
	3770 => "11111111",
	3771 => "11111111",
	3776 => "11111111",
	3777 => "11111111",
	3778 => "11111111",
	3779 => "11111111",
	3780 => "11111111",
	3781 => "11111111",
	3782 => "11111111",
	3783 => "11111111",
	3784 => "11111111",
	3785 => "11111111",
	3786 => "11111111",
	3787 => "11111111",
	3788 => "11111111",
	3789 => "11111111",
	3790 => "11111111",
	3791 => "11111111",
	3792 => "11111111",
	3793 => "11111111",
	3794 => "11111111",
	3795 => "11111111",
	3796 => "11111111",
	3797 => "11111111",
	3798 => "11111111",
	3799 => "11111111",
	3800 => "11111111",
	3801 => "11111111",
	3802 => "11111111",
	3803 => "11111111",
	3804 => "11111111",
	3805 => "11111111",
	3806 => "11111111",
	3807 => "11111111",
	3808 => "11111111",
	3809 => "11111111",
	3810 => "11111111",
	3811 => "11111111",
	3812 => "11111111",
	3813 => "11111111",
	3814 => "11111111",
	3815 => "11111111",
	3816 => "11111111",
	3817 => "11111111",
	3818 => "11111111",
	3819 => "11111111",
	3820 => "11111111",
	3821 => "11111111",
	3822 => "11111111",
	3823 => "11111111",
	3824 => "11111111",
	3825 => "11111111",
	3826 => "11111111",
	3827 => "11111111",
	3828 => "11111111",
	3829 => "11111111",
	3830 => "11111111",
	3831 => "11111111",
	3832 => "11111111",
	3833 => "11111111",
	3834 => "11111111",
	3835 => "11111111",

	others => (others => '0')
);

begin
	
	-- process ROM
	process (CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (EN = '1') then
				DATA <= ROM(conv_integer(ADDR));
			end if;
		end if;
	end process;
	
end Behavioral;

