		4140 => x"FF",
		4141 => x"FF",
		4142 => x"FF",
		4143 => x"FF",
		4144 => x"FF",
		4145 => x"FF",
		4146 => x"FF",
		4147 => x"FF",
		4148 => x"FF",
		4149 => x"FF",
		4150 => x"FF",
		4151 => x"FF",
		4152 => x"FF",
		4153 => x"FF",
		4154 => x"FF",
		4155 => x"FF",
		4156 => x"FF",
		4157 => x"FF",
		4158 => x"FF",
		4159 => x"FF",
		4160 => x"FF",
		4161 => x"FF",
		4162 => x"FF",
		4163 => x"FF",
		4164 => x"FF",
		4165 => x"FF",
		4166 => x"FF",
		4167 => x"FF",
		4168 => x"FF",
		4169 => x"FF",
		4170 => x"FF",
		4171 => x"FF",
		4172 => x"FF",
		4173 => x"FF",
		4174 => x"FF",
		4175 => x"FF",
		4176 => x"FF",
		4177 => x"FF",
		4178 => x"FF",
		4179 => x"FF",
		4180 => x"FF",
		4181 => x"FF",
		4182 => x"FF",
		4183 => x"FF",
		4184 => x"FF",
		4185 => x"FF",
		4186 => x"FF",
		4187 => x"FF",
		4188 => x"FF",
		4189 => x"FF",
		4190 => x"FF",
		4191 => x"FF",
		4192 => x"FF",
		4193 => x"FF",
		4194 => x"FF",
		4195 => x"FF",
		4196 => x"FF",
		4197 => x"FF",
		4198 => x"FF",
		4199 => x"FF",
		4200 => x"FF",
		4201 => x"FF",
		4202 => x"FF",
		4203 => x"FF",
		4204 => x"FF",
		4205 => x"FF",
		4206 => x"FF",
		4207 => x"FF",
		4208 => x"FF",
		4209 => x"FF",
		4210 => x"FF",
		4211 => x"FF",
		4212 => x"FF",
		4213 => x"FF",
		4214 => x"FF",
		4215 => x"FF",
		4216 => x"FF",
		4217 => x"FF",
		4218 => x"FF",
		4219 => x"FF",
		4220 => x"FF",
		4221 => x"FF",
		4222 => x"FF",
		4223 => x"FF",
		4224 => x"FF",
		4225 => x"FF",
		4226 => x"FF",
		4227 => x"FF",
		4228 => x"FF",
		4229 => x"FF",
		4230 => x"FF",
		4231 => x"FF",
		4232 => x"FF",
		4233 => x"FF",
		4234 => x"FF",
		4235 => x"FF",
		4236 => x"FF",
		4237 => x"FF",
		4238 => x"FF",
		4239 => x"FF",
		4240 => x"FF",
		4241 => x"FF",
		4242 => x"FF",
		4243 => x"FF",
		4244 => x"FF",
		4245 => x"FF",
		4246 => x"FF",
		4247 => x"FF",
		4248 => x"FF",
		4249 => x"FF",
		4250 => x"FF",
		4251 => x"FF",
		4252 => x"FF",
		4253 => x"FF",
		4254 => x"FF",
		4255 => x"FF",
		4256 => x"FF",
		4257 => x"FF",
		4258 => x"FF",
		4259 => x"FF",
		4260 => x"FF",
		4261 => x"FF",
		4262 => x"FF",
		4263 => x"FF",
		4264 => x"FF",
		4265 => x"FF",
		4266 => x"FF",
		4267 => x"FF",
		4268 => x"FF",
		4269 => x"FF",
		4270 => x"FF",
		4271 => x"FF",
		4272 => x"FF",
		4273 => x"FF",
		4274 => x"FF",
		4275 => x"FF",
		4276 => x"FF",
		4277 => x"FF",
		4278 => x"FF",
		4279 => x"FF",
		4280 => x"FF",
		4281 => x"FF",
		4282 => x"FF",
		4283 => x"FF",
		4284 => x"FF",
		4285 => x"FF",
		4286 => x"FF",
		4287 => x"FF",
		4288 => x"FF",
		4289 => x"FF",
		4290 => x"FF",
		4291 => x"FF",
		4292 => x"FF",
		4293 => x"FF",
		4294 => x"FF",
		4295 => x"FF",
		4296 => x"FF",
		4297 => x"FF",
		4298 => x"FF",
		4299 => x"FF",
		4300 => x"FF",
		4301 => x"FF",
		4302 => x"FF",
		4303 => x"FF",
		4304 => x"FF",
		4305 => x"FF",
		4306 => x"FF",
		4307 => x"FF",
		4308 => x"FF",
		4309 => x"FF",
		4310 => x"FF",
		4311 => x"FF",
		4312 => x"FF",
		4313 => x"FF",
		4314 => x"FF",
		4315 => x"FF",
		4316 => x"FF",
		4317 => x"FF",
		4318 => x"FF",
		4319 => x"FF",
		4320 => x"FF",
		4321 => x"FF",
		4322 => x"FF",
		4323 => x"FF",
		4324 => x"FF",
		4325 => x"FF",
		4326 => x"FF",
		4327 => x"FF",
		4328 => x"FF",
		4329 => x"FF",
		4330 => x"FF",
		4331 => x"FF",
		4332 => x"FF",
		4333 => x"FF",
		4334 => x"FF",
		4335 => x"FF",
		4336 => x"FF",
		4337 => x"FF",
		4338 => x"FF",
		4339 => x"FF",
		4340 => x"FF",
		4341 => x"FF",
		4342 => x"FF",
		4343 => x"FF",
		4344 => x"FF",
		4345 => x"FF",
		4346 => x"FF",
		4347 => x"FF",
		4348 => x"FF",
		4349 => x"FF",
		4350 => x"FF",
		4351 => x"FF",
		4352 => x"FF",
		4353 => x"FF",
		4354 => x"FF",
		4355 => x"FF",
		4356 => x"FF",
		4357 => x"FF",
		4358 => x"FF",
		4359 => x"FF",
		4360 => x"FF",
		4361 => x"FF",
		4362 => x"FF",
		4363 => x"FF",
		4364 => x"FF",
		4365 => x"FF",
		4366 => x"FF",
		4367 => x"FF",
		4368 => x"FF",
		4369 => x"FF",
		5164 => x"FF",
		5165 => x"FF",
		5166 => x"FF",
		5167 => x"FF",
		5168 => x"FF",
		5169 => x"FF",
		5170 => x"FF",
		5171 => x"FF",
		5172 => x"FF",
		5173 => x"FF",
		5174 => x"FF",
		5175 => x"FF",
		5176 => x"FF",
		5177 => x"FF",
		5178 => x"FF",
		5179 => x"FF",
		5180 => x"FF",
		5181 => x"FF",
		5182 => x"FF",
		5183 => x"FF",
		5184 => x"FF",
		5185 => x"FF",
		5186 => x"FF",
		5187 => x"FF",
		5188 => x"FF",
		5189 => x"FF",
		5190 => x"FF",
		5191 => x"FF",
		5192 => x"FF",
		5193 => x"FF",
		5194 => x"FF",
		5195 => x"FF",
		5196 => x"FF",
		5197 => x"FF",
		5198 => x"FF",
		5199 => x"FF",
		5200 => x"FF",
		5201 => x"FF",
		5202 => x"FF",
		5203 => x"FF",
		5204 => x"FF",
		5205 => x"FF",
		5206 => x"FF",
		5207 => x"FF",
		5208 => x"FF",
		5209 => x"FF",
		5210 => x"FF",
		5211 => x"FF",
		5212 => x"FF",
		5213 => x"FF",
		5214 => x"FF",
		5215 => x"FF",
		5216 => x"FF",
		5217 => x"FF",
		5218 => x"FF",
		5219 => x"FF",
		5220 => x"FF",
		5221 => x"FF",
		5222 => x"FF",
		5223 => x"FF",
		5224 => x"FF",
		5225 => x"FF",
		5226 => x"FF",
		5227 => x"FF",
		5228 => x"FF",
		5229 => x"FF",
		5230 => x"FF",
		5231 => x"FF",
		5232 => x"FF",
		5233 => x"FF",
		5234 => x"FF",
		5235 => x"FF",
		5236 => x"FF",
		5237 => x"FF",
		5238 => x"FF",
		5239 => x"FF",
		5240 => x"FF",
		5241 => x"FF",
		5242 => x"FF",
		5243 => x"FF",
		5244 => x"FF",
		5245 => x"FF",
		5246 => x"FF",
		5247 => x"FF",
		5248 => x"FF",
		5249 => x"FF",
		5250 => x"FF",
		5251 => x"FF",
		5252 => x"FF",
		5253 => x"FF",
		5254 => x"FF",
		5255 => x"FF",
		5256 => x"FF",
		5257 => x"FF",
		5258 => x"FF",
		5259 => x"FF",
		5260 => x"FF",
		5261 => x"FF",
		5262 => x"FF",
		5263 => x"FF",
		5264 => x"FF",
		5265 => x"FF",
		5266 => x"FF",
		5267 => x"FF",
		5268 => x"FF",
		5269 => x"FF",
		5270 => x"FF",
		5271 => x"FF",
		5272 => x"FF",
		5273 => x"FF",
		5274 => x"FF",
		5275 => x"FF",
		5276 => x"FF",
		5277 => x"FF",
		5278 => x"FF",
		5279 => x"FF",
		5280 => x"FF",
		5281 => x"FF",
		5282 => x"FF",
		5283 => x"FF",
		5284 => x"FF",
		5285 => x"FF",
		5286 => x"FF",
		5287 => x"FF",
		5288 => x"FF",
		5289 => x"FF",
		5290 => x"FF",
		5291 => x"FF",
		5292 => x"FF",
		5293 => x"FF",
		5294 => x"FF",
		5295 => x"FF",
		5296 => x"FF",
		5297 => x"FF",
		5298 => x"FF",
		5299 => x"FF",
		5300 => x"FF",
		5301 => x"FF",
		5302 => x"FF",
		5303 => x"FF",
		5304 => x"FF",
		5305 => x"FF",
		5306 => x"FF",
		5307 => x"FF",
		5308 => x"FF",
		5309 => x"FF",
		5310 => x"FF",
		5311 => x"FF",
		5312 => x"FF",
		5313 => x"FF",
		5314 => x"FF",
		5315 => x"FF",
		5316 => x"FF",
		5317 => x"FF",
		5318 => x"FF",
		5319 => x"FF",
		5320 => x"FF",
		5321 => x"FF",
		5322 => x"FF",
		5323 => x"FF",
		5324 => x"FF",
		5325 => x"FF",
		5326 => x"FF",
		5327 => x"FF",
		5328 => x"FF",
		5329 => x"FF",
		5330 => x"FF",
		5331 => x"FF",
		5332 => x"FF",
		5333 => x"FF",
		5334 => x"FF",
		5335 => x"FF",
		5336 => x"FF",
		5337 => x"FF",
		5338 => x"FF",
		5339 => x"FF",
		5340 => x"FF",
		5341 => x"FF",
		5342 => x"FF",
		5343 => x"FF",
		5344 => x"FF",
		5345 => x"FF",
		5346 => x"FF",
		5347 => x"FF",
		5348 => x"FF",
		5349 => x"FF",
		5350 => x"FF",
		5351 => x"FF",
		5352 => x"FF",
		5353 => x"FF",
		5354 => x"FF",
		5355 => x"FF",
		5356 => x"FF",
		5357 => x"FF",
		5358 => x"FF",
		5359 => x"FF",
		5360 => x"FF",
		5361 => x"FF",
		5362 => x"FF",
		5363 => x"FF",
		5364 => x"FF",
		5365 => x"FF",
		5366 => x"FF",
		5367 => x"FF",
		5368 => x"FF",
		5369 => x"FF",
		5370 => x"FF",
		5371 => x"FF",
		5372 => x"FF",
		5373 => x"FF",
		5374 => x"FF",
		5375 => x"FF",
		5376 => x"FF",
		5377 => x"FF",
		5378 => x"FF",
		5379 => x"FF",
		5380 => x"FF",
		5381 => x"FF",
		5382 => x"FF",
		5383 => x"FF",
		5384 => x"FF",
		5385 => x"FF",
		5386 => x"FF",
		5387 => x"FF",
		5388 => x"FF",
		5389 => x"FF",
		5390 => x"FF",
		5391 => x"FF",
		5392 => x"FF",
		5393 => x"FF",
		6188 => x"FF",
		6189 => x"FF",
		6190 => x"FF",
		6191 => x"FF",
		6192 => x"FF",
		6193 => x"FF",
		6194 => x"FF",
		6195 => x"FF",
		6196 => x"FF",
		6197 => x"FF",
		6198 => x"FF",
		6199 => x"FF",
		6200 => x"FF",
		6201 => x"FF",
		6202 => x"FF",
		6203 => x"FF",
		6204 => x"FF",
		6205 => x"FF",
		6206 => x"FF",
		6207 => x"FF",
		6208 => x"FF",
		6209 => x"FF",
		6210 => x"FF",
		6211 => x"FF",
		6212 => x"FF",
		6213 => x"FF",
		6214 => x"FF",
		6215 => x"FF",
		6216 => x"FF",
		6217 => x"FF",
		6218 => x"FF",
		6219 => x"FF",
		6220 => x"FF",
		6221 => x"FF",
		6222 => x"FF",
		6223 => x"FF",
		6224 => x"FF",
		6225 => x"FF",
		6226 => x"FF",
		6227 => x"FF",
		6228 => x"FF",
		6229 => x"FF",
		6230 => x"FF",
		6231 => x"FF",
		6232 => x"FF",
		6233 => x"FF",
		6234 => x"FF",
		6235 => x"FF",
		6236 => x"FF",
		6237 => x"FF",
		6238 => x"FF",
		6239 => x"FF",
		6240 => x"FF",
		6241 => x"FF",
		6242 => x"FF",
		6243 => x"FF",
		6244 => x"FF",
		6245 => x"FF",
		6246 => x"FF",
		6247 => x"FF",
		6248 => x"FF",
		6249 => x"FF",
		6250 => x"FF",
		6251 => x"FF",
		6252 => x"FF",
		6253 => x"FF",
		6254 => x"FF",
		6255 => x"FF",
		6256 => x"FF",
		6257 => x"FF",
		6258 => x"FF",
		6259 => x"FF",
		6260 => x"FF",
		6261 => x"FF",
		6262 => x"FF",
		6263 => x"FF",
		6264 => x"FF",
		6265 => x"FF",
		6266 => x"FF",
		6267 => x"FF",
		6268 => x"FF",
		6269 => x"FF",
		6270 => x"FF",
		6271 => x"FF",
		6272 => x"FF",
		6273 => x"FF",
		6274 => x"FF",
		6275 => x"FF",
		6276 => x"FF",
		6277 => x"FF",
		6278 => x"FF",
		6279 => x"FF",
		6280 => x"FF",
		6281 => x"FF",
		6282 => x"FF",
		6283 => x"FF",
		6284 => x"FF",
		6285 => x"FF",
		6286 => x"FF",
		6287 => x"FF",
		6288 => x"FF",
		6289 => x"FF",
		6290 => x"FF",
		6291 => x"FF",
		6292 => x"FF",
		6293 => x"FF",
		6294 => x"FF",
		6295 => x"FF",
		6296 => x"FF",
		6297 => x"FF",
		6298 => x"FF",
		6299 => x"FF",
		6300 => x"FF",
		6301 => x"FF",
		6302 => x"FF",
		6303 => x"FF",
		6304 => x"FF",
		6305 => x"FF",
		6306 => x"FF",
		6307 => x"FF",
		6308 => x"FF",
		6309 => x"FF",
		6310 => x"FF",
		6311 => x"FF",
		6312 => x"FF",
		6313 => x"FF",
		6314 => x"FF",
		6315 => x"FF",
		6316 => x"FF",
		6317 => x"FF",
		6318 => x"FF",
		6319 => x"FF",
		6320 => x"FF",
		6321 => x"FF",
		6322 => x"FF",
		6323 => x"FF",
		6324 => x"FF",
		6325 => x"FF",
		6326 => x"FF",
		6327 => x"FF",
		6328 => x"FF",
		6329 => x"FF",
		6330 => x"FF",
		6331 => x"FF",
		6332 => x"FF",
		6333 => x"FF",
		6334 => x"FF",
		6335 => x"FF",
		6336 => x"FF",
		6337 => x"FF",
		6338 => x"FF",
		6339 => x"FF",
		6340 => x"FF",
		6341 => x"FF",
		6342 => x"FF",
		6343 => x"FF",
		6344 => x"FF",
		6345 => x"FF",
		6346 => x"FF",
		6347 => x"FF",
		6348 => x"FF",
		6349 => x"FF",
		6350 => x"FF",
		6351 => x"FF",
		6352 => x"FF",
		6353 => x"FF",
		6354 => x"FF",
		6355 => x"FF",
		6356 => x"FF",
		6357 => x"FF",
		6358 => x"FF",
		6359 => x"FF",
		6360 => x"FF",
		6361 => x"FF",
		6362 => x"FF",
		6363 => x"FF",
		6364 => x"FF",
		6365 => x"FF",
		6366 => x"FF",
		6367 => x"FF",
		6368 => x"FF",
		6369 => x"FF",
		6370 => x"FF",
		6371 => x"FF",
		6372 => x"FF",
		6373 => x"FF",
		6374 => x"FF",
		6375 => x"FF",
		6376 => x"FF",
		6377 => x"FF",
		6378 => x"FF",
		6379 => x"FF",
		6380 => x"FF",
		6381 => x"FF",
		6382 => x"FF",
		6383 => x"FF",
		6384 => x"FF",
		6385 => x"FF",
		6386 => x"FF",
		6387 => x"FF",
		6388 => x"FF",
		6389 => x"FF",
		6390 => x"FF",
		6391 => x"FF",
		6392 => x"FF",
		6393 => x"FF",
		6394 => x"FF",
		6395 => x"FF",
		6396 => x"FF",
		6397 => x"FF",
		6398 => x"FF",
		6399 => x"FF",
		6400 => x"FF",
		6401 => x"FF",
		6402 => x"FF",
		6403 => x"FF",
		6404 => x"FF",
		6405 => x"FF",
		6406 => x"FF",
		6407 => x"FF",
		6408 => x"FF",
		6409 => x"FF",
		6410 => x"FF",
		6411 => x"FF",
		6412 => x"FF",
		6413 => x"FF",
		6414 => x"FF",
		6415 => x"FF",
		6416 => x"FF",
		6417 => x"FF",
		7212 => x"FF",
		7213 => x"FF",
		7214 => x"FF",
		7215 => x"FF",
		7216 => x"FF",
		7217 => x"FF",
		7218 => x"FF",
		7219 => x"FF",
		7220 => x"FF",
		7221 => x"FF",
		7222 => x"FF",
		7223 => x"FF",
		7224 => x"FF",
		7225 => x"FF",
		7226 => x"FF",
		7227 => x"FF",
		7228 => x"FF",
		7229 => x"FF",
		7230 => x"FF",
		7231 => x"FF",
		7232 => x"FF",
		7233 => x"FF",
		7234 => x"FF",
		7235 => x"FF",
		7236 => x"FF",
		7237 => x"FF",
		7238 => x"FF",
		7239 => x"FF",
		7240 => x"FF",
		7241 => x"FF",
		7242 => x"FF",
		7243 => x"FF",
		7244 => x"FF",
		7245 => x"FF",
		7246 => x"FF",
		7247 => x"FF",
		7248 => x"FF",
		7249 => x"FF",
		7250 => x"FF",
		7251 => x"FF",
		7252 => x"FF",
		7253 => x"FF",
		7254 => x"FF",
		7255 => x"FF",
		7256 => x"FF",
		7257 => x"FF",
		7258 => x"FF",
		7259 => x"FF",
		7260 => x"FF",
		7261 => x"FF",
		7262 => x"FF",
		7263 => x"FF",
		7264 => x"FF",
		7265 => x"FF",
		7266 => x"FF",
		7267 => x"FF",
		7268 => x"FF",
		7269 => x"FF",
		7270 => x"FF",
		7271 => x"FF",
		7272 => x"FF",
		7273 => x"FF",
		7274 => x"FF",
		7275 => x"FF",
		7276 => x"FF",
		7277 => x"FF",
		7278 => x"FF",
		7279 => x"FF",
		7280 => x"FF",
		7281 => x"FF",
		7282 => x"FF",
		7283 => x"FF",
		7284 => x"FF",
		7285 => x"FF",
		7286 => x"FF",
		7287 => x"FF",
		7288 => x"FF",
		7289 => x"FF",
		7290 => x"FF",
		7291 => x"FF",
		7292 => x"FF",
		7293 => x"FF",
		7294 => x"FF",
		7295 => x"FF",
		7296 => x"FF",
		7297 => x"FF",
		7298 => x"FF",
		7299 => x"FF",
		7300 => x"FF",
		7301 => x"FF",
		7302 => x"FF",
		7303 => x"FF",
		7304 => x"FF",
		7305 => x"FF",
		7306 => x"FF",
		7307 => x"FF",
		7308 => x"FF",
		7309 => x"FF",
		7310 => x"FF",
		7311 => x"FF",
		7312 => x"FF",
		7313 => x"FF",
		7314 => x"FF",
		7315 => x"FF",
		7316 => x"FF",
		7317 => x"FF",
		7318 => x"FF",
		7319 => x"FF",
		7320 => x"FF",
		7321 => x"FF",
		7322 => x"FF",
		7323 => x"FF",
		7324 => x"FF",
		7325 => x"FF",
		7326 => x"FF",
		7327 => x"FF",
		7328 => x"FF",
		7329 => x"FF",
		7330 => x"FF",
		7331 => x"FF",
		7332 => x"FF",
		7333 => x"FF",
		7334 => x"FF",
		7335 => x"FF",
		7336 => x"FF",
		7337 => x"FF",
		7338 => x"FF",
		7339 => x"FF",
		7340 => x"FF",
		7341 => x"FF",
		7342 => x"FF",
		7343 => x"FF",
		7344 => x"FF",
		7345 => x"FF",
		7346 => x"FF",
		7347 => x"FF",
		7348 => x"FF",
		7349 => x"FF",
		7350 => x"FF",
		7351 => x"FF",
		7352 => x"FF",
		7353 => x"FF",
		7354 => x"FF",
		7355 => x"FF",
		7356 => x"FF",
		7357 => x"FF",
		7358 => x"FF",
		7359 => x"FF",
		7360 => x"FF",
		7361 => x"FF",
		7362 => x"FF",
		7363 => x"FF",
		7364 => x"FF",
		7365 => x"FF",
		7366 => x"FF",
		7367 => x"FF",
		7368 => x"FF",
		7369 => x"FF",
		7370 => x"FF",
		7371 => x"FF",
		7372 => x"FF",
		7373 => x"FF",
		7374 => x"FF",
		7375 => x"FF",
		7376 => x"FF",
		7377 => x"FF",
		7378 => x"FF",
		7379 => x"FF",
		7380 => x"FF",
		7381 => x"FF",
		7382 => x"FF",
		7383 => x"FF",
		7384 => x"FF",
		7385 => x"FF",
		7386 => x"FF",
		7387 => x"FF",
		7388 => x"FF",
		7389 => x"FF",
		7390 => x"FF",
		7391 => x"FF",
		7392 => x"FF",
		7393 => x"FF",
		7394 => x"FF",
		7395 => x"FF",
		7396 => x"FF",
		7397 => x"FF",
		7398 => x"FF",
		7399 => x"FF",
		7400 => x"FF",
		7401 => x"FF",
		7402 => x"FF",
		7403 => x"FF",
		7404 => x"FF",
		7405 => x"FF",
		7406 => x"FF",
		7407 => x"FF",
		7408 => x"FF",
		7409 => x"FF",
		7410 => x"FF",
		7411 => x"FF",
		7412 => x"FF",
		7413 => x"FF",
		7414 => x"FF",
		7415 => x"FF",
		7416 => x"FF",
		7417 => x"FF",
		7418 => x"FF",
		7419 => x"FF",
		7420 => x"FF",
		7421 => x"FF",
		7422 => x"FF",
		7423 => x"FF",
		7424 => x"FF",
		7425 => x"FF",
		7426 => x"FF",
		7427 => x"FF",
		7428 => x"FF",
		7429 => x"FF",
		7430 => x"FF",
		7431 => x"FF",
		7432 => x"FF",
		7433 => x"FF",
		7434 => x"FF",
		7435 => x"FF",
		7436 => x"FF",
		7437 => x"FF",
		7438 => x"FF",
		7439 => x"FF",
		7440 => x"FF",
		7441 => x"FF",
		8236 => x"FF",
		8237 => x"FF",
		8238 => x"FF",
		8239 => x"FF",
		8240 => x"FF",
		8241 => x"FF",
		8242 => x"FF",
		8243 => x"FF",
		8244 => x"FF",
		8245 => x"FF",
		8246 => x"FF",
		8247 => x"FF",
		8248 => x"FF",
		8249 => x"FF",
		8250 => x"FF",
		8251 => x"FF",
		8252 => x"FF",
		8253 => x"FF",
		8254 => x"FF",
		8255 => x"FF",
		8256 => x"FF",
		8257 => x"FF",
		8258 => x"FF",
		8259 => x"FF",
		8260 => x"FF",
		8261 => x"FF",
		8262 => x"FF",
		8263 => x"FF",
		8264 => x"FF",
		8265 => x"FF",
		8266 => x"FF",
		8267 => x"FF",
		8268 => x"FF",
		8269 => x"FF",
		8270 => x"FF",
		8271 => x"FF",
		8272 => x"FF",
		8273 => x"FF",
		8274 => x"FF",
		8275 => x"FF",
		8276 => x"FF",
		8277 => x"FF",
		8278 => x"FF",
		8279 => x"FF",
		8280 => x"FF",
		8281 => x"FF",
		8282 => x"FF",
		8283 => x"FF",
		8284 => x"FF",
		8285 => x"FF",
		8286 => x"FF",
		8287 => x"FF",
		8288 => x"FF",
		8289 => x"FF",
		8290 => x"FF",
		8291 => x"FF",
		8292 => x"FF",
		8293 => x"FF",
		8294 => x"FF",
		8295 => x"FF",
		8296 => x"FF",
		8297 => x"FF",
		8298 => x"FF",
		8299 => x"FF",
		8300 => x"FF",
		8301 => x"FF",
		8302 => x"FF",
		8303 => x"FF",
		8304 => x"FF",
		8305 => x"FF",
		8306 => x"FF",
		8307 => x"FF",
		8308 => x"FF",
		8309 => x"FF",
		8310 => x"FF",
		8311 => x"FF",
		8312 => x"FF",
		8313 => x"FF",
		8314 => x"FF",
		8315 => x"FF",
		8316 => x"FF",
		8317 => x"FF",
		8318 => x"FF",
		8319 => x"FF",
		8320 => x"FF",
		8321 => x"FF",
		8322 => x"FF",
		8323 => x"FF",
		8324 => x"FF",
		8325 => x"FF",
		8326 => x"FF",
		8327 => x"FF",
		8328 => x"FF",
		8329 => x"FF",
		8330 => x"FF",
		8331 => x"FF",
		8332 => x"FF",
		8333 => x"FF",
		8334 => x"FF",
		8335 => x"FF",
		8336 => x"FF",
		8337 => x"FF",
		8338 => x"FF",
		8339 => x"FF",
		8340 => x"FF",
		8341 => x"FF",
		8342 => x"FF",
		8343 => x"FF",
		8344 => x"FF",
		8345 => x"FF",
		8346 => x"FF",
		8347 => x"FF",
		8348 => x"FF",
		8349 => x"FF",
		8350 => x"FF",
		8351 => x"FF",
		8352 => x"FF",
		8353 => x"FF",
		8354 => x"FF",
		8355 => x"FF",
		8356 => x"FF",
		8357 => x"FF",
		8358 => x"FF",
		8359 => x"FF",
		8360 => x"FF",
		8361 => x"FF",
		8362 => x"FF",
		8363 => x"FF",
		8364 => x"FF",
		8365 => x"FF",
		8366 => x"FF",
		8367 => x"FF",
		8368 => x"FF",
		8369 => x"FF",
		8370 => x"FF",
		8371 => x"FF",
		8372 => x"FF",
		8373 => x"FF",
		8374 => x"FF",
		8375 => x"FF",
		8376 => x"FF",
		8377 => x"FF",
		8378 => x"FF",
		8379 => x"FF",
		8380 => x"FF",
		8381 => x"FF",
		8382 => x"FF",
		8383 => x"FF",
		8384 => x"FF",
		8385 => x"FF",
		8386 => x"FF",
		8387 => x"FF",
		8388 => x"FF",
		8389 => x"FF",
		8390 => x"FF",
		8391 => x"FF",
		8392 => x"FF",
		8393 => x"FF",
		8394 => x"FF",
		8395 => x"FF",
		8396 => x"FF",
		8397 => x"FF",
		8398 => x"FF",
		8399 => x"FF",
		8400 => x"FF",
		8401 => x"FF",
		8402 => x"FF",
		8403 => x"FF",
		8404 => x"FF",
		8405 => x"FF",
		8406 => x"FF",
		8407 => x"FF",
		8408 => x"FF",
		8409 => x"FF",
		8410 => x"FF",
		8411 => x"FF",
		8412 => x"FF",
		8413 => x"FF",
		8414 => x"FF",
		8415 => x"FF",
		8416 => x"FF",
		8417 => x"FF",
		8418 => x"FF",
		8419 => x"FF",
		8420 => x"FF",
		8421 => x"FF",
		8422 => x"FF",
		8423 => x"FF",
		8424 => x"FF",
		8425 => x"FF",
		8426 => x"FF",
		8427 => x"FF",
		8428 => x"FF",
		8429 => x"FF",
		8430 => x"FF",
		8431 => x"FF",
		8432 => x"FF",
		8433 => x"FF",
		8434 => x"FF",
		8435 => x"FF",
		8436 => x"FF",
		8437 => x"FF",
		8438 => x"FF",
		8439 => x"FF",
		8440 => x"FF",
		8441 => x"FF",
		8442 => x"FF",
		8443 => x"FF",
		8444 => x"FF",
		8445 => x"FF",
		8446 => x"FF",
		8447 => x"FF",
		8448 => x"FF",
		8449 => x"FF",
		8450 => x"FF",
		8451 => x"FF",
		8452 => x"FF",
		8453 => x"FF",
		8454 => x"FF",
		8455 => x"FF",
		8456 => x"FF",
		8457 => x"FF",
		8458 => x"FF",
		8459 => x"FF",
		8460 => x"FF",
		8461 => x"FF",
		8462 => x"FF",
		8463 => x"FF",
		8464 => x"FF",
		8465 => x"FF",
		9260 => x"FF",
		9261 => x"FF",
		9262 => x"FF",
		9263 => x"FF",
		9264 => x"FF",
		9335 => x"FF",
		9336 => x"FF",
		9337 => x"FF",
		9338 => x"FF",
		9339 => x"FF",
		9410 => x"FF",
		9411 => x"FF",
		9412 => x"FF",
		9413 => x"FF",
		9414 => x"FF",
		9485 => x"FF",
		9486 => x"FF",
		9487 => x"FF",
		9488 => x"FF",
		9489 => x"FF",
		10284 => x"FF",
		10285 => x"FF",
		10286 => x"FF",
		10287 => x"FF",
		10288 => x"FF",
		10359 => x"FF",
		10360 => x"FF",
		10361 => x"FF",
		10362 => x"FF",
		10363 => x"FF",
		10434 => x"FF",
		10435 => x"FF",
		10436 => x"FF",
		10437 => x"FF",
		10438 => x"FF",
		10509 => x"FF",
		10510 => x"FF",
		10511 => x"FF",
		10512 => x"FF",
		10513 => x"FF",
		11308 => x"FF",
		11309 => x"FF",
		11310 => x"FF",
		11311 => x"FF",
		11312 => x"FF",
		11383 => x"FF",
		11384 => x"FF",
		11385 => x"FF",
		11386 => x"FF",
		11387 => x"FF",
		11458 => x"FF",
		11459 => x"FF",
		11460 => x"FF",
		11461 => x"FF",
		11462 => x"FF",
		11533 => x"FF",
		11534 => x"FF",
		11535 => x"FF",
		11536 => x"FF",
		11537 => x"FF",
		12332 => x"FF",
		12333 => x"FF",
		12334 => x"FF",
		12335 => x"FF",
		12336 => x"FF",
		12407 => x"FF",
		12408 => x"FF",
		12409 => x"FF",
		12410 => x"FF",
		12411 => x"FF",
		12482 => x"FF",
		12483 => x"FF",
		12484 => x"FF",
		12485 => x"FF",
		12486 => x"FF",
		12557 => x"FF",
		12558 => x"FF",
		12559 => x"FF",
		12560 => x"FF",
		12561 => x"FF",
		13356 => x"FF",
		13357 => x"FF",
		13358 => x"FF",
		13359 => x"FF",
		13360 => x"FF",
		13431 => x"FF",
		13432 => x"FF",
		13433 => x"FF",
		13434 => x"FF",
		13435 => x"FF",
		13506 => x"FF",
		13507 => x"FF",
		13508 => x"FF",
		13509 => x"FF",
		13510 => x"FF",
		13581 => x"FF",
		13582 => x"FF",
		13583 => x"FF",
		13584 => x"FF",
		13585 => x"FF",
		14380 => x"FF",
		14381 => x"FF",
		14382 => x"FF",
		14383 => x"FF",
		14384 => x"FF",
		14455 => x"FF",
		14456 => x"FF",
		14457 => x"FF",
		14458 => x"FF",
		14459 => x"FF",
		14530 => x"FF",
		14531 => x"FF",
		14532 => x"FF",
		14533 => x"FF",
		14534 => x"FF",
		14605 => x"FF",
		14606 => x"FF",
		14607 => x"FF",
		14608 => x"FF",
		14609 => x"FF",
		15404 => x"FF",
		15405 => x"FF",
		15406 => x"FF",
		15407 => x"FF",
		15408 => x"FF",
		15479 => x"FF",
		15480 => x"FF",
		15481 => x"FF",
		15482 => x"FF",
		15483 => x"FF",
		15554 => x"FF",
		15555 => x"FF",
		15556 => x"FF",
		15557 => x"FF",
		15558 => x"FF",
		15629 => x"FF",
		15630 => x"FF",
		15631 => x"FF",
		15632 => x"FF",
		15633 => x"FF",
		16428 => x"FF",
		16429 => x"FF",
		16430 => x"FF",
		16431 => x"FF",
		16432 => x"FF",
		16503 => x"FF",
		16504 => x"FF",
		16505 => x"FF",
		16506 => x"FF",
		16507 => x"FF",
		16578 => x"FF",
		16579 => x"FF",
		16580 => x"FF",
		16581 => x"FF",
		16582 => x"FF",
		16653 => x"FF",
		16654 => x"FF",
		16655 => x"FF",
		16656 => x"FF",
		16657 => x"FF",
		17452 => x"FF",
		17453 => x"FF",
		17454 => x"FF",
		17455 => x"FF",
		17456 => x"FF",
		17527 => x"FF",
		17528 => x"FF",
		17529 => x"FF",
		17530 => x"FF",
		17531 => x"FF",
		17602 => x"FF",
		17603 => x"FF",
		17604 => x"FF",
		17605 => x"FF",
		17606 => x"FF",
		17677 => x"FF",
		17678 => x"FF",
		17679 => x"FF",
		17680 => x"FF",
		17681 => x"FF",
		18476 => x"FF",
		18477 => x"FF",
		18478 => x"FF",
		18479 => x"FF",
		18480 => x"FF",
		18551 => x"FF",
		18552 => x"FF",
		18553 => x"FF",
		18554 => x"FF",
		18555 => x"FF",
		18626 => x"FF",
		18627 => x"FF",
		18628 => x"FF",
		18629 => x"FF",
		18630 => x"FF",
		18701 => x"FF",
		18702 => x"FF",
		18703 => x"FF",
		18704 => x"FF",
		18705 => x"FF",
		19500 => x"FF",
		19501 => x"FF",
		19502 => x"FF",
		19503 => x"FF",
		19504 => x"FF",
		19575 => x"FF",
		19576 => x"FF",
		19577 => x"FF",
		19578 => x"FF",
		19579 => x"FF",
		19650 => x"FF",
		19651 => x"FF",
		19652 => x"FF",
		19653 => x"FF",
		19654 => x"FF",
		19725 => x"FF",
		19726 => x"FF",
		19727 => x"FF",
		19728 => x"FF",
		19729 => x"FF",
		20524 => x"FF",
		20525 => x"FF",
		20526 => x"FF",
		20527 => x"FF",
		20528 => x"FF",
		20599 => x"FF",
		20600 => x"FF",
		20601 => x"FF",
		20602 => x"FF",
		20603 => x"FF",
		20674 => x"FF",
		20675 => x"FF",
		20676 => x"FF",
		20677 => x"FF",
		20678 => x"FF",
		20749 => x"FF",
		20750 => x"FF",
		20751 => x"FF",
		20752 => x"FF",
		20753 => x"FF",
		21548 => x"FF",
		21549 => x"FF",
		21550 => x"FF",
		21551 => x"FF",
		21552 => x"FF",
		21623 => x"FF",
		21624 => x"FF",
		21625 => x"FF",
		21626 => x"FF",
		21627 => x"FF",
		21698 => x"FF",
		21699 => x"FF",
		21700 => x"FF",
		21701 => x"FF",
		21702 => x"FF",
		21773 => x"FF",
		21774 => x"FF",
		21775 => x"FF",
		21776 => x"FF",
		21777 => x"FF",
		22572 => x"FF",
		22573 => x"FF",
		22574 => x"FF",
		22575 => x"FF",
		22576 => x"FF",
		22647 => x"FF",
		22648 => x"FF",
		22649 => x"FF",
		22650 => x"FF",
		22651 => x"FF",
		22722 => x"FF",
		22723 => x"FF",
		22724 => x"FF",
		22725 => x"FF",
		22726 => x"FF",
		22797 => x"FF",
		22798 => x"FF",
		22799 => x"FF",
		22800 => x"FF",
		22801 => x"FF",
		23596 => x"FF",
		23597 => x"FF",
		23598 => x"FF",
		23599 => x"FF",
		23600 => x"FF",
		23671 => x"FF",
		23672 => x"FF",
		23673 => x"FF",
		23674 => x"FF",
		23675 => x"FF",
		23746 => x"FF",
		23747 => x"FF",
		23748 => x"FF",
		23749 => x"FF",
		23750 => x"FF",
		23821 => x"FF",
		23822 => x"FF",
		23823 => x"FF",
		23824 => x"FF",
		23825 => x"FF",
		24620 => x"FF",
		24621 => x"FF",
		24622 => x"FF",
		24623 => x"FF",
		24624 => x"FF",
		24695 => x"FF",
		24696 => x"FF",
		24697 => x"FF",
		24698 => x"FF",
		24699 => x"FF",
		24770 => x"FF",
		24771 => x"FF",
		24772 => x"FF",
		24773 => x"FF",
		24774 => x"FF",
		24845 => x"FF",
		24846 => x"FF",
		24847 => x"FF",
		24848 => x"FF",
		24849 => x"FF",
		25644 => x"FF",
		25645 => x"FF",
		25646 => x"FF",
		25647 => x"FF",
		25648 => x"FF",
		25719 => x"FF",
		25720 => x"FF",
		25721 => x"FF",
		25722 => x"FF",
		25723 => x"FF",
		25794 => x"FF",
		25795 => x"FF",
		25796 => x"FF",
		25797 => x"FF",
		25798 => x"FF",
		25869 => x"FF",
		25870 => x"FF",
		25871 => x"FF",
		25872 => x"FF",
		25873 => x"FF",
		26668 => x"FF",
		26669 => x"FF",
		26670 => x"FF",
		26671 => x"FF",
		26672 => x"FF",
		26743 => x"FF",
		26744 => x"FF",
		26745 => x"FF",
		26746 => x"FF",
		26747 => x"FF",
		26818 => x"FF",
		26819 => x"FF",
		26820 => x"FF",
		26821 => x"FF",
		26822 => x"FF",
		26893 => x"FF",
		26894 => x"FF",
		26895 => x"FF",
		26896 => x"FF",
		26897 => x"FF",
		27692 => x"FF",
		27693 => x"FF",
		27694 => x"FF",
		27695 => x"FF",
		27696 => x"FF",
		27767 => x"FF",
		27768 => x"FF",
		27769 => x"FF",
		27770 => x"FF",
		27771 => x"FF",
		27842 => x"FF",
		27843 => x"FF",
		27844 => x"FF",
		27845 => x"FF",
		27846 => x"FF",
		27917 => x"FF",
		27918 => x"FF",
		27919 => x"FF",
		27920 => x"FF",
		27921 => x"FF",
		28716 => x"FF",
		28717 => x"FF",
		28718 => x"FF",
		28719 => x"FF",
		28720 => x"FF",
		28791 => x"FF",
		28792 => x"FF",
		28793 => x"FF",
		28794 => x"FF",
		28795 => x"FF",
		28866 => x"FF",
		28867 => x"FF",
		28868 => x"FF",
		28869 => x"FF",
		28870 => x"FF",
		28941 => x"FF",
		28942 => x"FF",
		28943 => x"FF",
		28944 => x"FF",
		28945 => x"FF",
		29740 => x"FF",
		29741 => x"FF",
		29742 => x"FF",
		29743 => x"FF",
		29744 => x"FF",
		29815 => x"FF",
		29816 => x"FF",
		29817 => x"FF",
		29818 => x"FF",
		29819 => x"FF",
		29890 => x"FF",
		29891 => x"FF",
		29892 => x"FF",
		29893 => x"FF",
		29894 => x"FF",
		29965 => x"FF",
		29966 => x"FF",
		29967 => x"FF",
		29968 => x"FF",
		29969 => x"FF",
		30764 => x"FF",
		30765 => x"FF",
		30766 => x"FF",
		30767 => x"FF",
		30768 => x"FF",
		30839 => x"FF",
		30840 => x"FF",
		30841 => x"FF",
		30842 => x"FF",
		30843 => x"FF",
		30914 => x"FF",
		30915 => x"FF",
		30916 => x"FF",
		30917 => x"FF",
		30918 => x"FF",
		30989 => x"FF",
		30990 => x"FF",
		30991 => x"FF",
		30992 => x"FF",
		30993 => x"FF",
		31788 => x"FF",
		31789 => x"FF",
		31790 => x"FF",
		31791 => x"FF",
		31792 => x"FF",
		31863 => x"FF",
		31864 => x"FF",
		31865 => x"FF",
		31866 => x"FF",
		31867 => x"FF",
		31938 => x"FF",
		31939 => x"FF",
		31940 => x"FF",
		31941 => x"FF",
		31942 => x"FF",
		32013 => x"FF",
		32014 => x"FF",
		32015 => x"FF",
		32016 => x"FF",
		32017 => x"FF",
		32812 => x"FF",
		32813 => x"FF",
		32814 => x"FF",
		32815 => x"FF",
		32816 => x"FF",
		32887 => x"FF",
		32888 => x"FF",
		32889 => x"FF",
		32890 => x"FF",
		32891 => x"FF",
		32962 => x"FF",
		32963 => x"FF",
		32964 => x"FF",
		32965 => x"FF",
		32966 => x"FF",
		33037 => x"FF",
		33038 => x"FF",
		33039 => x"FF",
		33040 => x"FF",
		33041 => x"FF",
		33836 => x"FF",
		33837 => x"FF",
		33838 => x"FF",
		33839 => x"FF",
		33840 => x"FF",
		33911 => x"FF",
		33912 => x"FF",
		33913 => x"FF",
		33914 => x"FF",
		33915 => x"FF",
		33986 => x"FF",
		33987 => x"FF",
		33988 => x"FF",
		33989 => x"FF",
		33990 => x"FF",
		34061 => x"FF",
		34062 => x"FF",
		34063 => x"FF",
		34064 => x"FF",
		34065 => x"FF",
		34860 => x"FF",
		34861 => x"FF",
		34862 => x"FF",
		34863 => x"FF",
		34864 => x"FF",
		34935 => x"FF",
		34936 => x"FF",
		34937 => x"FF",
		34938 => x"FF",
		34939 => x"FF",
		35010 => x"FF",
		35011 => x"FF",
		35012 => x"FF",
		35013 => x"FF",
		35014 => x"FF",
		35085 => x"FF",
		35086 => x"FF",
		35087 => x"FF",
		35088 => x"FF",
		35089 => x"FF",
		35884 => x"FF",
		35885 => x"FF",
		35886 => x"FF",
		35887 => x"FF",
		35888 => x"FF",
		35959 => x"FF",
		35960 => x"FF",
		35961 => x"FF",
		35962 => x"FF",
		35963 => x"FF",
		36034 => x"FF",
		36035 => x"FF",
		36036 => x"FF",
		36037 => x"FF",
		36038 => x"FF",
		36109 => x"FF",
		36110 => x"FF",
		36111 => x"FF",
		36112 => x"FF",
		36113 => x"FF",
		36908 => x"FF",
		36909 => x"FF",
		36910 => x"FF",
		36911 => x"FF",
		36912 => x"FF",
		36983 => x"FF",
		36984 => x"FF",
		36985 => x"FF",
		36986 => x"FF",
		36987 => x"FF",
		37058 => x"FF",
		37059 => x"FF",
		37060 => x"FF",
		37061 => x"FF",
		37062 => x"FF",
		37133 => x"FF",
		37134 => x"FF",
		37135 => x"FF",
		37136 => x"FF",
		37137 => x"FF",
		37932 => x"FF",
		37933 => x"FF",
		37934 => x"FF",
		37935 => x"FF",
		37936 => x"FF",
		38007 => x"FF",
		38008 => x"FF",
		38009 => x"FF",
		38010 => x"FF",
		38011 => x"FF",
		38082 => x"FF",
		38083 => x"FF",
		38084 => x"FF",
		38085 => x"FF",
		38086 => x"FF",
		38157 => x"FF",
		38158 => x"FF",
		38159 => x"FF",
		38160 => x"FF",
		38161 => x"FF",
		38956 => x"FF",
		38957 => x"FF",
		38958 => x"FF",
		38959 => x"FF",
		38960 => x"FF",
		39031 => x"FF",
		39032 => x"FF",
		39033 => x"FF",
		39034 => x"FF",
		39035 => x"FF",
		39106 => x"FF",
		39107 => x"FF",
		39108 => x"FF",
		39109 => x"FF",
		39110 => x"FF",
		39181 => x"FF",
		39182 => x"FF",
		39183 => x"FF",
		39184 => x"FF",
		39185 => x"FF",
		39980 => x"FF",
		39981 => x"FF",
		39982 => x"FF",
		39983 => x"FF",
		39984 => x"FF",
		40055 => x"FF",
		40056 => x"FF",
		40057 => x"FF",
		40058 => x"FF",
		40059 => x"FF",
		40130 => x"FF",
		40131 => x"FF",
		40132 => x"FF",
		40133 => x"FF",
		40134 => x"FF",
		40205 => x"FF",
		40206 => x"FF",
		40207 => x"FF",
		40208 => x"FF",
		40209 => x"FF",
		41004 => x"FF",
		41005 => x"FF",
		41006 => x"FF",
		41007 => x"FF",
		41008 => x"FF",
		41079 => x"FF",
		41080 => x"FF",
		41081 => x"FF",
		41082 => x"FF",
		41083 => x"FF",
		41154 => x"FF",
		41155 => x"FF",
		41156 => x"FF",
		41157 => x"FF",
		41158 => x"FF",
		41229 => x"FF",
		41230 => x"FF",
		41231 => x"FF",
		41232 => x"FF",
		41233 => x"FF",
		42028 => x"FF",
		42029 => x"FF",
		42030 => x"FF",
		42031 => x"FF",
		42032 => x"FF",
		42103 => x"FF",
		42104 => x"FF",
		42105 => x"FF",
		42106 => x"FF",
		42107 => x"FF",
		42178 => x"FF",
		42179 => x"FF",
		42180 => x"FF",
		42181 => x"FF",
		42182 => x"FF",
		42253 => x"FF",
		42254 => x"FF",
		42255 => x"FF",
		42256 => x"FF",
		42257 => x"FF",
		43052 => x"FF",
		43053 => x"FF",
		43054 => x"FF",
		43055 => x"FF",
		43056 => x"FF",
		43127 => x"FF",
		43128 => x"FF",
		43129 => x"FF",
		43130 => x"FF",
		43131 => x"FF",
		43202 => x"FF",
		43203 => x"FF",
		43204 => x"FF",
		43205 => x"FF",
		43206 => x"FF",
		43277 => x"FF",
		43278 => x"FF",
		43279 => x"FF",
		43280 => x"FF",
		43281 => x"FF",
		44076 => x"FF",
		44077 => x"FF",
		44078 => x"FF",
		44079 => x"FF",
		44080 => x"FF",
		44151 => x"FF",
		44152 => x"FF",
		44153 => x"FF",
		44154 => x"FF",
		44155 => x"FF",
		44226 => x"FF",
		44227 => x"FF",
		44228 => x"FF",
		44229 => x"FF",
		44230 => x"FF",
		44301 => x"FF",
		44302 => x"FF",
		44303 => x"FF",
		44304 => x"FF",
		44305 => x"FF",
		45100 => x"FF",
		45101 => x"FF",
		45102 => x"FF",
		45103 => x"FF",
		45104 => x"FF",
		45175 => x"FF",
		45176 => x"FF",
		45177 => x"FF",
		45178 => x"FF",
		45179 => x"FF",
		45250 => x"FF",
		45251 => x"FF",
		45252 => x"FF",
		45253 => x"FF",
		45254 => x"FF",
		45325 => x"FF",
		45326 => x"FF",
		45327 => x"FF",
		45328 => x"FF",
		45329 => x"FF",
		46124 => x"FF",
		46125 => x"FF",
		46126 => x"FF",
		46127 => x"FF",
		46128 => x"FF",
		46199 => x"FF",
		46200 => x"FF",
		46201 => x"FF",
		46202 => x"FF",
		46203 => x"FF",
		46274 => x"FF",
		46275 => x"FF",
		46276 => x"FF",
		46277 => x"FF",
		46278 => x"FF",
		46349 => x"FF",
		46350 => x"FF",
		46351 => x"FF",
		46352 => x"FF",
		46353 => x"FF",
		47148 => x"FF",
		47149 => x"FF",
		47150 => x"FF",
		47151 => x"FF",
		47152 => x"FF",
		47223 => x"FF",
		47224 => x"FF",
		47225 => x"FF",
		47226 => x"FF",
		47227 => x"FF",
		47298 => x"FF",
		47299 => x"FF",
		47300 => x"FF",
		47301 => x"FF",
		47302 => x"FF",
		47373 => x"FF",
		47374 => x"FF",
		47375 => x"FF",
		47376 => x"FF",
		47377 => x"FF",
		48172 => x"FF",
		48173 => x"FF",
		48174 => x"FF",
		48175 => x"FF",
		48176 => x"FF",
		48247 => x"FF",
		48248 => x"FF",
		48249 => x"FF",
		48250 => x"FF",
		48251 => x"FF",
		48322 => x"FF",
		48323 => x"FF",
		48324 => x"FF",
		48325 => x"FF",
		48326 => x"FF",
		48397 => x"FF",
		48398 => x"FF",
		48399 => x"FF",
		48400 => x"FF",
		48401 => x"FF",
		49196 => x"FF",
		49197 => x"FF",
		49198 => x"FF",
		49199 => x"FF",
		49200 => x"FF",
		49271 => x"FF",
		49272 => x"FF",
		49273 => x"FF",
		49274 => x"FF",
		49275 => x"FF",
		49346 => x"FF",
		49347 => x"FF",
		49348 => x"FF",
		49349 => x"FF",
		49350 => x"FF",
		49421 => x"FF",
		49422 => x"FF",
		49423 => x"FF",
		49424 => x"FF",
		49425 => x"FF",
		50220 => x"FF",
		50221 => x"FF",
		50222 => x"FF",
		50223 => x"FF",
		50224 => x"FF",
		50295 => x"FF",
		50296 => x"FF",
		50297 => x"FF",
		50298 => x"FF",
		50299 => x"FF",
		50370 => x"FF",
		50371 => x"FF",
		50372 => x"FF",
		50373 => x"FF",
		50374 => x"FF",
		50445 => x"FF",
		50446 => x"FF",
		50447 => x"FF",
		50448 => x"FF",
		50449 => x"FF",
		51244 => x"FF",
		51245 => x"FF",
		51246 => x"FF",
		51247 => x"FF",
		51248 => x"FF",
		51319 => x"FF",
		51320 => x"FF",
		51321 => x"FF",
		51322 => x"FF",
		51323 => x"FF",
		51394 => x"FF",
		51395 => x"FF",
		51396 => x"FF",
		51397 => x"FF",
		51398 => x"FF",
		51469 => x"FF",
		51470 => x"FF",
		51471 => x"FF",
		51472 => x"FF",
		51473 => x"FF",
		52268 => x"FF",
		52269 => x"FF",
		52270 => x"FF",
		52271 => x"FF",
		52272 => x"FF",
		52343 => x"FF",
		52344 => x"FF",
		52345 => x"FF",
		52346 => x"FF",
		52347 => x"FF",
		52418 => x"FF",
		52419 => x"FF",
		52420 => x"FF",
		52421 => x"FF",
		52422 => x"FF",
		52493 => x"FF",
		52494 => x"FF",
		52495 => x"FF",
		52496 => x"FF",
		52497 => x"FF",
		53292 => x"FF",
		53293 => x"FF",
		53294 => x"FF",
		53295 => x"FF",
		53296 => x"FF",
		53367 => x"FF",
		53368 => x"FF",
		53369 => x"FF",
		53370 => x"FF",
		53371 => x"FF",
		53442 => x"FF",
		53443 => x"FF",
		53444 => x"FF",
		53445 => x"FF",
		53446 => x"FF",
		53517 => x"FF",
		53518 => x"FF",
		53519 => x"FF",
		53520 => x"FF",
		53521 => x"FF",
		54316 => x"FF",
		54317 => x"FF",
		54318 => x"FF",
		54319 => x"FF",
		54320 => x"FF",
		54391 => x"FF",
		54392 => x"FF",
		54393 => x"FF",
		54394 => x"FF",
		54395 => x"FF",
		54466 => x"FF",
		54467 => x"FF",
		54468 => x"FF",
		54469 => x"FF",
		54470 => x"FF",
		54541 => x"FF",
		54542 => x"FF",
		54543 => x"FF",
		54544 => x"FF",
		54545 => x"FF",
		55340 => x"FF",
		55341 => x"FF",
		55342 => x"FF",
		55343 => x"FF",
		55344 => x"FF",
		55415 => x"FF",
		55416 => x"FF",
		55417 => x"FF",
		55418 => x"FF",
		55419 => x"FF",
		55490 => x"FF",
		55491 => x"FF",
		55492 => x"FF",
		55493 => x"FF",
		55494 => x"FF",
		55565 => x"FF",
		55566 => x"FF",
		55567 => x"FF",
		55568 => x"FF",
		55569 => x"FF",
		56364 => x"FF",
		56365 => x"FF",
		56366 => x"FF",
		56367 => x"FF",
		56368 => x"FF",
		56439 => x"FF",
		56440 => x"FF",
		56441 => x"FF",
		56442 => x"FF",
		56443 => x"FF",
		56514 => x"FF",
		56515 => x"FF",
		56516 => x"FF",
		56517 => x"FF",
		56518 => x"FF",
		56589 => x"FF",
		56590 => x"FF",
		56591 => x"FF",
		56592 => x"FF",
		56593 => x"FF",
		57388 => x"FF",
		57389 => x"FF",
		57390 => x"FF",
		57391 => x"FF",
		57392 => x"FF",
		57463 => x"FF",
		57464 => x"FF",
		57465 => x"FF",
		57466 => x"FF",
		57467 => x"FF",
		57538 => x"FF",
		57539 => x"FF",
		57540 => x"FF",
		57541 => x"FF",
		57542 => x"FF",
		57613 => x"FF",
		57614 => x"FF",
		57615 => x"FF",
		57616 => x"FF",
		57617 => x"FF",
		58412 => x"FF",
		58413 => x"FF",
		58414 => x"FF",
		58415 => x"FF",
		58416 => x"FF",
		58487 => x"FF",
		58488 => x"FF",
		58489 => x"FF",
		58490 => x"FF",
		58491 => x"FF",
		58562 => x"FF",
		58563 => x"FF",
		58564 => x"FF",
		58565 => x"FF",
		58566 => x"FF",
		58637 => x"FF",
		58638 => x"FF",
		58639 => x"FF",
		58640 => x"FF",
		58641 => x"FF",
		59436 => x"FF",
		59437 => x"FF",
		59438 => x"FF",
		59439 => x"FF",
		59440 => x"FF",
		59511 => x"FF",
		59512 => x"FF",
		59513 => x"FF",
		59514 => x"FF",
		59515 => x"FF",
		59586 => x"FF",
		59587 => x"FF",
		59588 => x"FF",
		59589 => x"FF",
		59590 => x"FF",
		59661 => x"FF",
		59662 => x"FF",
		59663 => x"FF",
		59664 => x"FF",
		59665 => x"FF",
		60460 => x"FF",
		60461 => x"FF",
		60462 => x"FF",
		60463 => x"FF",
		60464 => x"FF",
		60535 => x"FF",
		60536 => x"FF",
		60537 => x"FF",
		60538 => x"FF",
		60539 => x"FF",
		60610 => x"FF",
		60611 => x"FF",
		60612 => x"FF",
		60613 => x"FF",
		60614 => x"FF",
		60685 => x"FF",
		60686 => x"FF",
		60687 => x"FF",
		60688 => x"FF",
		60689 => x"FF",
		61484 => x"FF",
		61485 => x"FF",
		61486 => x"FF",
		61487 => x"FF",
		61488 => x"FF",
		61559 => x"FF",
		61560 => x"FF",
		61561 => x"FF",
		61562 => x"FF",
		61563 => x"FF",
		61634 => x"FF",
		61635 => x"FF",
		61636 => x"FF",
		61637 => x"FF",
		61638 => x"FF",
		61709 => x"FF",
		61710 => x"FF",
		61711 => x"FF",
		61712 => x"FF",
		61713 => x"FF",
		62508 => x"FF",
		62509 => x"FF",
		62510 => x"FF",
		62511 => x"FF",
		62512 => x"FF",
		62583 => x"FF",
		62584 => x"FF",
		62585 => x"FF",
		62586 => x"FF",
		62587 => x"FF",
		62658 => x"FF",
		62659 => x"FF",
		62660 => x"FF",
		62661 => x"FF",
		62662 => x"FF",
		62733 => x"FF",
		62734 => x"FF",
		62735 => x"FF",
		62736 => x"FF",
		62737 => x"FF",
		63532 => x"FF",
		63533 => x"FF",
		63534 => x"FF",
		63535 => x"FF",
		63536 => x"FF",
		63607 => x"FF",
		63608 => x"FF",
		63609 => x"FF",
		63610 => x"FF",
		63611 => x"FF",
		63682 => x"FF",
		63683 => x"FF",
		63684 => x"FF",
		63685 => x"FF",
		63686 => x"FF",
		63757 => x"FF",
		63758 => x"FF",
		63759 => x"FF",
		63760 => x"FF",
		63761 => x"FF",
		64556 => x"FF",
		64557 => x"FF",
		64558 => x"FF",
		64559 => x"FF",
		64560 => x"FF",
		64631 => x"FF",
		64632 => x"FF",
		64633 => x"FF",
		64634 => x"FF",
		64635 => x"FF",
		64706 => x"FF",
		64707 => x"FF",
		64708 => x"FF",
		64709 => x"FF",
		64710 => x"FF",
		64781 => x"FF",
		64782 => x"FF",
		64783 => x"FF",
		64784 => x"FF",
		64785 => x"FF",
		65580 => x"FF",
		65581 => x"FF",
		65582 => x"FF",
		65583 => x"FF",
		65584 => x"FF",
		65655 => x"FF",
		65656 => x"FF",
		65657 => x"FF",
		65658 => x"FF",
		65659 => x"FF",
		65730 => x"FF",
		65731 => x"FF",
		65732 => x"FF",
		65733 => x"FF",
		65734 => x"FF",
		65805 => x"FF",
		65806 => x"FF",
		65807 => x"FF",
		65808 => x"FF",
		65809 => x"FF",
		66604 => x"FF",
		66605 => x"FF",
		66606 => x"FF",
		66607 => x"FF",
		66608 => x"FF",
		66679 => x"FF",
		66680 => x"FF",
		66681 => x"FF",
		66682 => x"FF",
		66683 => x"FF",
		66754 => x"FF",
		66755 => x"FF",
		66756 => x"FF",
		66757 => x"FF",
		66758 => x"FF",
		66829 => x"FF",
		66830 => x"FF",
		66831 => x"FF",
		66832 => x"FF",
		66833 => x"FF",
		67628 => x"FF",
		67629 => x"FF",
		67630 => x"FF",
		67631 => x"FF",
		67632 => x"FF",
		67703 => x"FF",
		67704 => x"FF",
		67705 => x"FF",
		67706 => x"FF",
		67707 => x"FF",
		67778 => x"FF",
		67779 => x"FF",
		67780 => x"FF",
		67781 => x"FF",
		67782 => x"FF",
		67853 => x"FF",
		67854 => x"FF",
		67855 => x"FF",
		67856 => x"FF",
		67857 => x"FF",
		68652 => x"FF",
		68653 => x"FF",
		68654 => x"FF",
		68655 => x"FF",
		68656 => x"FF",
		68727 => x"FF",
		68728 => x"FF",
		68729 => x"FF",
		68730 => x"FF",
		68731 => x"FF",
		68802 => x"FF",
		68803 => x"FF",
		68804 => x"FF",
		68805 => x"FF",
		68806 => x"FF",
		68877 => x"FF",
		68878 => x"FF",
		68879 => x"FF",
		68880 => x"FF",
		68881 => x"FF",
		69676 => x"FF",
		69677 => x"FF",
		69678 => x"FF",
		69679 => x"FF",
		69680 => x"FF",
		69751 => x"FF",
		69752 => x"FF",
		69753 => x"FF",
		69754 => x"FF",
		69755 => x"FF",
		69826 => x"FF",
		69827 => x"FF",
		69828 => x"FF",
		69829 => x"FF",
		69830 => x"FF",
		69901 => x"FF",
		69902 => x"FF",
		69903 => x"FF",
		69904 => x"FF",
		69905 => x"FF",
		70700 => x"FF",
		70701 => x"FF",
		70702 => x"FF",
		70703 => x"FF",
		70704 => x"FF",
		70775 => x"FF",
		70776 => x"FF",
		70777 => x"FF",
		70778 => x"FF",
		70779 => x"FF",
		70850 => x"FF",
		70851 => x"FF",
		70852 => x"FF",
		70853 => x"FF",
		70854 => x"FF",
		70925 => x"FF",
		70926 => x"FF",
		70927 => x"FF",
		70928 => x"FF",
		70929 => x"FF",
		71724 => x"FF",
		71725 => x"FF",
		71726 => x"FF",
		71727 => x"FF",
		71728 => x"FF",
		71799 => x"FF",
		71800 => x"FF",
		71801 => x"FF",
		71802 => x"FF",
		71803 => x"FF",
		71874 => x"FF",
		71875 => x"FF",
		71876 => x"FF",
		71877 => x"FF",
		71878 => x"FF",
		71949 => x"FF",
		71950 => x"FF",
		71951 => x"FF",
		71952 => x"FF",
		71953 => x"FF",
		72748 => x"FF",
		72749 => x"FF",
		72750 => x"FF",
		72751 => x"FF",
		72752 => x"FF",
		72823 => x"FF",
		72824 => x"FF",
		72825 => x"FF",
		72826 => x"FF",
		72827 => x"FF",
		72898 => x"FF",
		72899 => x"FF",
		72900 => x"FF",
		72901 => x"FF",
		72902 => x"FF",
		72973 => x"FF",
		72974 => x"FF",
		72975 => x"FF",
		72976 => x"FF",
		72977 => x"FF",
		73772 => x"FF",
		73773 => x"FF",
		73774 => x"FF",
		73775 => x"FF",
		73776 => x"FF",
		73847 => x"FF",
		73848 => x"FF",
		73849 => x"FF",
		73850 => x"FF",
		73851 => x"FF",
		73922 => x"FF",
		73923 => x"FF",
		73924 => x"FF",
		73925 => x"FF",
		73926 => x"FF",
		73997 => x"FF",
		73998 => x"FF",
		73999 => x"FF",
		74000 => x"FF",
		74001 => x"FF",
		74796 => x"FF",
		74797 => x"FF",
		74798 => x"FF",
		74799 => x"FF",
		74800 => x"FF",
		74871 => x"FF",
		74872 => x"FF",
		74873 => x"FF",
		74874 => x"FF",
		74875 => x"FF",
		74946 => x"FF",
		74947 => x"FF",
		74948 => x"FF",
		74949 => x"FF",
		74950 => x"FF",
		75021 => x"FF",
		75022 => x"FF",
		75023 => x"FF",
		75024 => x"FF",
		75025 => x"FF",
		75820 => x"FF",
		75821 => x"FF",
		75822 => x"FF",
		75823 => x"FF",
		75824 => x"FF",
		75895 => x"FF",
		75896 => x"FF",
		75897 => x"FF",
		75898 => x"FF",
		75899 => x"FF",
		75970 => x"FF",
		75971 => x"FF",
		75972 => x"FF",
		75973 => x"FF",
		75974 => x"FF",
		76045 => x"FF",
		76046 => x"FF",
		76047 => x"FF",
		76048 => x"FF",
		76049 => x"FF",
		76844 => x"FF",
		76845 => x"FF",
		76846 => x"FF",
		76847 => x"FF",
		76848 => x"FF",
		76919 => x"FF",
		76920 => x"FF",
		76921 => x"FF",
		76922 => x"FF",
		76923 => x"FF",
		76994 => x"FF",
		76995 => x"FF",
		76996 => x"FF",
		76997 => x"FF",
		76998 => x"FF",
		77069 => x"FF",
		77070 => x"FF",
		77071 => x"FF",
		77072 => x"FF",
		77073 => x"FF",
		77868 => x"FF",
		77869 => x"FF",
		77870 => x"FF",
		77871 => x"FF",
		77872 => x"FF",
		77943 => x"FF",
		77944 => x"FF",
		77945 => x"FF",
		77946 => x"FF",
		77947 => x"FF",
		78018 => x"FF",
		78019 => x"FF",
		78020 => x"FF",
		78021 => x"FF",
		78022 => x"FF",
		78093 => x"FF",
		78094 => x"FF",
		78095 => x"FF",
		78096 => x"FF",
		78097 => x"FF",
		78892 => x"FF",
		78893 => x"FF",
		78894 => x"FF",
		78895 => x"FF",
		78896 => x"FF",
		78967 => x"FF",
		78968 => x"FF",
		78969 => x"FF",
		78970 => x"FF",
		78971 => x"FF",
		79042 => x"FF",
		79043 => x"FF",
		79044 => x"FF",
		79045 => x"FF",
		79046 => x"FF",
		79117 => x"FF",
		79118 => x"FF",
		79119 => x"FF",
		79120 => x"FF",
		79121 => x"FF",
		79916 => x"FF",
		79917 => x"FF",
		79918 => x"FF",
		79919 => x"FF",
		79920 => x"FF",
		79991 => x"FF",
		79992 => x"FF",
		79993 => x"FF",
		79994 => x"FF",
		79995 => x"FF",
		80066 => x"FF",
		80067 => x"FF",
		80068 => x"FF",
		80069 => x"FF",
		80070 => x"FF",
		80141 => x"FF",
		80142 => x"FF",
		80143 => x"FF",
		80144 => x"FF",
		80145 => x"FF",
		80940 => x"FF",
		80941 => x"FF",
		80942 => x"FF",
		80943 => x"FF",
		80944 => x"FF",
		80945 => x"FF",
		80946 => x"FF",
		80947 => x"FF",
		80948 => x"FF",
		80949 => x"FF",
		80950 => x"FF",
		80951 => x"FF",
		80952 => x"FF",
		80953 => x"FF",
		80954 => x"FF",
		80955 => x"FF",
		80956 => x"FF",
		80957 => x"FF",
		80958 => x"FF",
		80959 => x"FF",
		80960 => x"FF",
		80961 => x"FF",
		80962 => x"FF",
		80963 => x"FF",
		80964 => x"FF",
		80965 => x"FF",
		80966 => x"FF",
		80967 => x"FF",
		80968 => x"FF",
		80969 => x"FF",
		80970 => x"FF",
		80971 => x"FF",
		80972 => x"FF",
		80973 => x"FF",
		80974 => x"FF",
		80975 => x"FF",
		80976 => x"FF",
		80977 => x"FF",
		80978 => x"FF",
		80979 => x"FF",
		80980 => x"FF",
		80981 => x"FF",
		80982 => x"FF",
		80983 => x"FF",
		80984 => x"FF",
		80985 => x"FF",
		80986 => x"FF",
		80987 => x"FF",
		80988 => x"FF",
		80989 => x"FF",
		80990 => x"FF",
		80991 => x"FF",
		80992 => x"FF",
		80993 => x"FF",
		80994 => x"FF",
		80995 => x"FF",
		80996 => x"FF",
		80997 => x"FF",
		80998 => x"FF",
		80999 => x"FF",
		81000 => x"FF",
		81001 => x"FF",
		81002 => x"FF",
		81003 => x"FF",
		81004 => x"FF",
		81005 => x"FF",
		81006 => x"FF",
		81007 => x"FF",
		81008 => x"FF",
		81009 => x"FF",
		81010 => x"FF",
		81011 => x"FF",
		81012 => x"FF",
		81013 => x"FF",
		81014 => x"FF",
		81015 => x"FF",
		81016 => x"FF",
		81017 => x"FF",
		81018 => x"FF",
		81019 => x"FF",
		81020 => x"FF",
		81021 => x"FF",
		81022 => x"FF",
		81023 => x"FF",
		81024 => x"FF",
		81025 => x"FF",
		81026 => x"FF",
		81027 => x"FF",
		81028 => x"FF",
		81029 => x"FF",
		81030 => x"FF",
		81031 => x"FF",
		81032 => x"FF",
		81033 => x"FF",
		81034 => x"FF",
		81035 => x"FF",
		81036 => x"FF",
		81037 => x"FF",
		81038 => x"FF",
		81039 => x"FF",
		81040 => x"FF",
		81041 => x"FF",
		81042 => x"FF",
		81043 => x"FF",
		81044 => x"FF",
		81045 => x"FF",
		81046 => x"FF",
		81047 => x"FF",
		81048 => x"FF",
		81049 => x"FF",
		81050 => x"FF",
		81051 => x"FF",
		81052 => x"FF",
		81053 => x"FF",
		81054 => x"FF",
		81055 => x"FF",
		81056 => x"FF",
		81057 => x"FF",
		81058 => x"FF",
		81059 => x"FF",
		81060 => x"FF",
		81061 => x"FF",
		81062 => x"FF",
		81063 => x"FF",
		81064 => x"FF",
		81065 => x"FF",
		81066 => x"FF",
		81067 => x"FF",
		81068 => x"FF",
		81069 => x"FF",
		81070 => x"FF",
		81071 => x"FF",
		81072 => x"FF",
		81073 => x"FF",
		81074 => x"FF",
		81075 => x"FF",
		81076 => x"FF",
		81077 => x"FF",
		81078 => x"FF",
		81079 => x"FF",
		81080 => x"FF",
		81081 => x"FF",
		81082 => x"FF",
		81083 => x"FF",
		81084 => x"FF",
		81085 => x"FF",
		81086 => x"FF",
		81087 => x"FF",
		81088 => x"FF",
		81089 => x"FF",
		81090 => x"FF",
		81091 => x"FF",
		81092 => x"FF",
		81093 => x"FF",
		81094 => x"FF",
		81095 => x"FF",
		81096 => x"FF",
		81097 => x"FF",
		81098 => x"FF",
		81099 => x"FF",
		81100 => x"FF",
		81101 => x"FF",
		81102 => x"FF",
		81103 => x"FF",
		81104 => x"FF",
		81105 => x"FF",
		81106 => x"FF",
		81107 => x"FF",
		81108 => x"FF",
		81109 => x"FF",
		81110 => x"FF",
		81111 => x"FF",
		81112 => x"FF",
		81113 => x"FF",
		81114 => x"FF",
		81115 => x"FF",
		81116 => x"FF",
		81117 => x"FF",
		81118 => x"FF",
		81119 => x"FF",
		81120 => x"FF",
		81121 => x"FF",
		81122 => x"FF",
		81123 => x"FF",
		81124 => x"FF",
		81125 => x"FF",
		81126 => x"FF",
		81127 => x"FF",
		81128 => x"FF",
		81129 => x"FF",
		81130 => x"FF",
		81131 => x"FF",
		81132 => x"FF",
		81133 => x"FF",
		81134 => x"FF",
		81135 => x"FF",
		81136 => x"FF",
		81137 => x"FF",
		81138 => x"FF",
		81139 => x"FF",
		81140 => x"FF",
		81141 => x"FF",
		81142 => x"FF",
		81143 => x"FF",
		81144 => x"FF",
		81145 => x"FF",
		81146 => x"FF",
		81147 => x"FF",
		81148 => x"FF",
		81149 => x"FF",
		81150 => x"FF",
		81151 => x"FF",
		81152 => x"FF",
		81153 => x"FF",
		81154 => x"FF",
		81155 => x"FF",
		81156 => x"FF",
		81157 => x"FF",
		81158 => x"FF",
		81159 => x"FF",
		81160 => x"FF",
		81161 => x"FF",
		81162 => x"FF",
		81163 => x"FF",
		81164 => x"FF",
		81165 => x"FF",
		81166 => x"FF",
		81167 => x"FF",
		81168 => x"FF",
		81169 => x"FF",
		81964 => x"FF",
		81965 => x"FF",
		81966 => x"FF",
		81967 => x"FF",
		81968 => x"FF",
		81969 => x"FF",
		81970 => x"FF",
		81971 => x"FF",
		81972 => x"FF",
		81973 => x"FF",
		81974 => x"FF",
		81975 => x"FF",
		81976 => x"FF",
		81977 => x"FF",
		81978 => x"FF",
		81979 => x"FF",
		81980 => x"FF",
		81981 => x"FF",
		81982 => x"FF",
		81983 => x"FF",
		81984 => x"FF",
		81985 => x"FF",
		81986 => x"FF",
		81987 => x"FF",
		81988 => x"FF",
		81989 => x"FF",
		81990 => x"FF",
		81991 => x"FF",
		81992 => x"FF",
		81993 => x"FF",
		81994 => x"FF",
		81995 => x"FF",
		81996 => x"FF",
		81997 => x"FF",
		81998 => x"FF",
		81999 => x"FF",
		82000 => x"FF",
		82001 => x"FF",
		82002 => x"FF",
		82003 => x"FF",
		82004 => x"FF",
		82005 => x"FF",
		82006 => x"FF",
		82007 => x"FF",
		82008 => x"FF",
		82009 => x"FF",
		82010 => x"FF",
		82011 => x"FF",
		82012 => x"FF",
		82013 => x"FF",
		82014 => x"FF",
		82015 => x"FF",
		82016 => x"FF",
		82017 => x"FF",
		82018 => x"FF",
		82019 => x"FF",
		82020 => x"FF",
		82021 => x"FF",
		82022 => x"FF",
		82023 => x"FF",
		82024 => x"FF",
		82025 => x"FF",
		82026 => x"FF",
		82027 => x"FF",
		82028 => x"FF",
		82029 => x"FF",
		82030 => x"FF",
		82031 => x"FF",
		82032 => x"FF",
		82033 => x"FF",
		82034 => x"FF",
		82035 => x"FF",
		82036 => x"FF",
		82037 => x"FF",
		82038 => x"FF",
		82039 => x"FF",
		82040 => x"FF",
		82041 => x"FF",
		82042 => x"FF",
		82043 => x"FF",
		82044 => x"FF",
		82045 => x"FF",
		82046 => x"FF",
		82047 => x"FF",
		82048 => x"FF",
		82049 => x"FF",
		82050 => x"FF",
		82051 => x"FF",
		82052 => x"FF",
		82053 => x"FF",
		82054 => x"FF",
		82055 => x"FF",
		82056 => x"FF",
		82057 => x"FF",
		82058 => x"FF",
		82059 => x"FF",
		82060 => x"FF",
		82061 => x"FF",
		82062 => x"FF",
		82063 => x"FF",
		82064 => x"FF",
		82065 => x"FF",
		82066 => x"FF",
		82067 => x"FF",
		82068 => x"FF",
		82069 => x"FF",
		82070 => x"FF",
		82071 => x"FF",
		82072 => x"FF",
		82073 => x"FF",
		82074 => x"FF",
		82075 => x"FF",
		82076 => x"FF",
		82077 => x"FF",
		82078 => x"FF",
		82079 => x"FF",
		82080 => x"FF",
		82081 => x"FF",
		82082 => x"FF",
		82083 => x"FF",
		82084 => x"FF",
		82085 => x"FF",
		82086 => x"FF",
		82087 => x"FF",
		82088 => x"FF",
		82089 => x"FF",
		82090 => x"FF",
		82091 => x"FF",
		82092 => x"FF",
		82093 => x"FF",
		82094 => x"FF",
		82095 => x"FF",
		82096 => x"FF",
		82097 => x"FF",
		82098 => x"FF",
		82099 => x"FF",
		82100 => x"FF",
		82101 => x"FF",
		82102 => x"FF",
		82103 => x"FF",
		82104 => x"FF",
		82105 => x"FF",
		82106 => x"FF",
		82107 => x"FF",
		82108 => x"FF",
		82109 => x"FF",
		82110 => x"FF",
		82111 => x"FF",
		82112 => x"FF",
		82113 => x"FF",
		82114 => x"FF",
		82115 => x"FF",
		82116 => x"FF",
		82117 => x"FF",
		82118 => x"FF",
		82119 => x"FF",
		82120 => x"FF",
		82121 => x"FF",
		82122 => x"FF",
		82123 => x"FF",
		82124 => x"FF",
		82125 => x"FF",
		82126 => x"FF",
		82127 => x"FF",
		82128 => x"FF",
		82129 => x"FF",
		82130 => x"FF",
		82131 => x"FF",
		82132 => x"FF",
		82133 => x"FF",
		82134 => x"FF",
		82135 => x"FF",
		82136 => x"FF",
		82137 => x"FF",
		82138 => x"FF",
		82139 => x"FF",
		82140 => x"FF",
		82141 => x"FF",
		82142 => x"FF",
		82143 => x"FF",
		82144 => x"FF",
		82145 => x"FF",
		82146 => x"FF",
		82147 => x"FF",
		82148 => x"FF",
		82149 => x"FF",
		82150 => x"FF",
		82151 => x"FF",
		82152 => x"FF",
		82153 => x"FF",
		82154 => x"FF",
		82155 => x"FF",
		82156 => x"FF",
		82157 => x"FF",
		82158 => x"FF",
		82159 => x"FF",
		82160 => x"FF",
		82161 => x"FF",
		82162 => x"FF",
		82163 => x"FF",
		82164 => x"FF",
		82165 => x"FF",
		82166 => x"FF",
		82167 => x"FF",
		82168 => x"FF",
		82169 => x"FF",
		82170 => x"FF",
		82171 => x"FF",
		82172 => x"FF",
		82173 => x"FF",
		82174 => x"FF",
		82175 => x"FF",
		82176 => x"FF",
		82177 => x"FF",
		82178 => x"FF",
		82179 => x"FF",
		82180 => x"FF",
		82181 => x"FF",
		82182 => x"FF",
		82183 => x"FF",
		82184 => x"FF",
		82185 => x"FF",
		82186 => x"FF",
		82187 => x"FF",
		82188 => x"FF",
		82189 => x"FF",
		82190 => x"FF",
		82191 => x"FF",
		82192 => x"FF",
		82193 => x"FF",
		82988 => x"FF",
		82989 => x"FF",
		82990 => x"FF",
		82991 => x"FF",
		82992 => x"FF",
		82993 => x"FF",
		82994 => x"FF",
		82995 => x"FF",
		82996 => x"FF",
		82997 => x"FF",
		82998 => x"FF",
		82999 => x"FF",
		83000 => x"FF",
		83001 => x"FF",
		83002 => x"FF",
		83003 => x"FF",
		83004 => x"FF",
		83005 => x"FF",
		83006 => x"FF",
		83007 => x"FF",
		83008 => x"FF",
		83009 => x"FF",
		83010 => x"FF",
		83011 => x"FF",
		83012 => x"FF",
		83013 => x"FF",
		83014 => x"FF",
		83015 => x"FF",
		83016 => x"FF",
		83017 => x"FF",
		83018 => x"FF",
		83019 => x"FF",
		83020 => x"FF",
		83021 => x"FF",
		83022 => x"FF",
		83023 => x"FF",
		83024 => x"FF",
		83025 => x"FF",
		83026 => x"FF",
		83027 => x"FF",
		83028 => x"FF",
		83029 => x"FF",
		83030 => x"FF",
		83031 => x"FF",
		83032 => x"FF",
		83033 => x"FF",
		83034 => x"FF",
		83035 => x"FF",
		83036 => x"FF",
		83037 => x"FF",
		83038 => x"FF",
		83039 => x"FF",
		83040 => x"FF",
		83041 => x"FF",
		83042 => x"FF",
		83043 => x"FF",
		83044 => x"FF",
		83045 => x"FF",
		83046 => x"FF",
		83047 => x"FF",
		83048 => x"FF",
		83049 => x"FF",
		83050 => x"FF",
		83051 => x"FF",
		83052 => x"FF",
		83053 => x"FF",
		83054 => x"FF",
		83055 => x"FF",
		83056 => x"FF",
		83057 => x"FF",
		83058 => x"FF",
		83059 => x"FF",
		83060 => x"FF",
		83061 => x"FF",
		83062 => x"FF",
		83063 => x"FF",
		83064 => x"FF",
		83065 => x"FF",
		83066 => x"FF",
		83067 => x"FF",
		83068 => x"FF",
		83069 => x"FF",
		83070 => x"FF",
		83071 => x"FF",
		83072 => x"FF",
		83073 => x"FF",
		83074 => x"FF",
		83075 => x"FF",
		83076 => x"FF",
		83077 => x"FF",
		83078 => x"FF",
		83079 => x"FF",
		83080 => x"FF",
		83081 => x"FF",
		83082 => x"FF",
		83083 => x"FF",
		83084 => x"FF",
		83085 => x"FF",
		83086 => x"FF",
		83087 => x"FF",
		83088 => x"FF",
		83089 => x"FF",
		83090 => x"FF",
		83091 => x"FF",
		83092 => x"FF",
		83093 => x"FF",
		83094 => x"FF",
		83095 => x"FF",
		83096 => x"FF",
		83097 => x"FF",
		83098 => x"FF",
		83099 => x"FF",
		83100 => x"FF",
		83101 => x"FF",
		83102 => x"FF",
		83103 => x"FF",
		83104 => x"FF",
		83105 => x"FF",
		83106 => x"FF",
		83107 => x"FF",
		83108 => x"FF",
		83109 => x"FF",
		83110 => x"FF",
		83111 => x"FF",
		83112 => x"FF",
		83113 => x"FF",
		83114 => x"FF",
		83115 => x"FF",
		83116 => x"FF",
		83117 => x"FF",
		83118 => x"FF",
		83119 => x"FF",
		83120 => x"FF",
		83121 => x"FF",
		83122 => x"FF",
		83123 => x"FF",
		83124 => x"FF",
		83125 => x"FF",
		83126 => x"FF",
		83127 => x"FF",
		83128 => x"FF",
		83129 => x"FF",
		83130 => x"FF",
		83131 => x"FF",
		83132 => x"FF",
		83133 => x"FF",
		83134 => x"FF",
		83135 => x"FF",
		83136 => x"FF",
		83137 => x"FF",
		83138 => x"FF",
		83139 => x"FF",
		83140 => x"FF",
		83141 => x"FF",
		83142 => x"FF",
		83143 => x"FF",
		83144 => x"FF",
		83145 => x"FF",
		83146 => x"FF",
		83147 => x"FF",
		83148 => x"FF",
		83149 => x"FF",
		83150 => x"FF",
		83151 => x"FF",
		83152 => x"FF",
		83153 => x"FF",
		83154 => x"FF",
		83155 => x"FF",
		83156 => x"FF",
		83157 => x"FF",
		83158 => x"FF",
		83159 => x"FF",
		83160 => x"FF",
		83161 => x"FF",
		83162 => x"FF",
		83163 => x"FF",
		83164 => x"FF",
		83165 => x"FF",
		83166 => x"FF",
		83167 => x"FF",
		83168 => x"FF",
		83169 => x"FF",
		83170 => x"FF",
		83171 => x"FF",
		83172 => x"FF",
		83173 => x"FF",
		83174 => x"FF",
		83175 => x"FF",
		83176 => x"FF",
		83177 => x"FF",
		83178 => x"FF",
		83179 => x"FF",
		83180 => x"FF",
		83181 => x"FF",
		83182 => x"FF",
		83183 => x"FF",
		83184 => x"FF",
		83185 => x"FF",
		83186 => x"FF",
		83187 => x"FF",
		83188 => x"FF",
		83189 => x"FF",
		83190 => x"FF",
		83191 => x"FF",
		83192 => x"FF",
		83193 => x"FF",
		83194 => x"FF",
		83195 => x"FF",
		83196 => x"FF",
		83197 => x"FF",
		83198 => x"FF",
		83199 => x"FF",
		83200 => x"FF",
		83201 => x"FF",
		83202 => x"FF",
		83203 => x"FF",
		83204 => x"FF",
		83205 => x"FF",
		83206 => x"FF",
		83207 => x"FF",
		83208 => x"FF",
		83209 => x"FF",
		83210 => x"FF",
		83211 => x"FF",
		83212 => x"FF",
		83213 => x"FF",
		83214 => x"FF",
		83215 => x"FF",
		83216 => x"FF",
		83217 => x"FF",
		84012 => x"FF",
		84013 => x"FF",
		84014 => x"FF",
		84015 => x"FF",
		84016 => x"FF",
		84017 => x"FF",
		84018 => x"FF",
		84019 => x"FF",
		84020 => x"FF",
		84021 => x"FF",
		84022 => x"FF",
		84023 => x"FF",
		84024 => x"FF",
		84025 => x"FF",
		84026 => x"FF",
		84027 => x"FF",
		84028 => x"FF",
		84029 => x"FF",
		84030 => x"FF",
		84031 => x"FF",
		84032 => x"FF",
		84033 => x"FF",
		84034 => x"FF",
		84035 => x"FF",
		84036 => x"FF",
		84037 => x"FF",
		84038 => x"FF",
		84039 => x"FF",
		84040 => x"FF",
		84041 => x"FF",
		84042 => x"FF",
		84043 => x"FF",
		84044 => x"FF",
		84045 => x"FF",
		84046 => x"FF",
		84047 => x"FF",
		84048 => x"FF",
		84049 => x"FF",
		84050 => x"FF",
		84051 => x"FF",
		84052 => x"FF",
		84053 => x"FF",
		84054 => x"FF",
		84055 => x"FF",
		84056 => x"FF",
		84057 => x"FF",
		84058 => x"FF",
		84059 => x"FF",
		84060 => x"FF",
		84061 => x"FF",
		84062 => x"FF",
		84063 => x"FF",
		84064 => x"FF",
		84065 => x"FF",
		84066 => x"FF",
		84067 => x"FF",
		84068 => x"FF",
		84069 => x"FF",
		84070 => x"FF",
		84071 => x"FF",
		84072 => x"FF",
		84073 => x"FF",
		84074 => x"FF",
		84075 => x"FF",
		84076 => x"FF",
		84077 => x"FF",
		84078 => x"FF",
		84079 => x"FF",
		84080 => x"FF",
		84081 => x"FF",
		84082 => x"FF",
		84083 => x"FF",
		84084 => x"FF",
		84085 => x"FF",
		84086 => x"FF",
		84087 => x"FF",
		84088 => x"FF",
		84089 => x"FF",
		84090 => x"FF",
		84091 => x"FF",
		84092 => x"FF",
		84093 => x"FF",
		84094 => x"FF",
		84095 => x"FF",
		84096 => x"FF",
		84097 => x"FF",
		84098 => x"FF",
		84099 => x"FF",
		84100 => x"FF",
		84101 => x"FF",
		84102 => x"FF",
		84103 => x"FF",
		84104 => x"FF",
		84105 => x"FF",
		84106 => x"FF",
		84107 => x"FF",
		84108 => x"FF",
		84109 => x"FF",
		84110 => x"FF",
		84111 => x"FF",
		84112 => x"FF",
		84113 => x"FF",
		84114 => x"FF",
		84115 => x"FF",
		84116 => x"FF",
		84117 => x"FF",
		84118 => x"FF",
		84119 => x"FF",
		84120 => x"FF",
		84121 => x"FF",
		84122 => x"FF",
		84123 => x"FF",
		84124 => x"FF",
		84125 => x"FF",
		84126 => x"FF",
		84127 => x"FF",
		84128 => x"FF",
		84129 => x"FF",
		84130 => x"FF",
		84131 => x"FF",
		84132 => x"FF",
		84133 => x"FF",
		84134 => x"FF",
		84135 => x"FF",
		84136 => x"FF",
		84137 => x"FF",
		84138 => x"FF",
		84139 => x"FF",
		84140 => x"FF",
		84141 => x"FF",
		84142 => x"FF",
		84143 => x"FF",
		84144 => x"FF",
		84145 => x"FF",
		84146 => x"FF",
		84147 => x"FF",
		84148 => x"FF",
		84149 => x"FF",
		84150 => x"FF",
		84151 => x"FF",
		84152 => x"FF",
		84153 => x"FF",
		84154 => x"FF",
		84155 => x"FF",
		84156 => x"FF",
		84157 => x"FF",
		84158 => x"FF",
		84159 => x"FF",
		84160 => x"FF",
		84161 => x"FF",
		84162 => x"FF",
		84163 => x"FF",
		84164 => x"FF",
		84165 => x"FF",
		84166 => x"FF",
		84167 => x"FF",
		84168 => x"FF",
		84169 => x"FF",
		84170 => x"FF",
		84171 => x"FF",
		84172 => x"FF",
		84173 => x"FF",
		84174 => x"FF",
		84175 => x"FF",
		84176 => x"FF",
		84177 => x"FF",
		84178 => x"FF",
		84179 => x"FF",
		84180 => x"FF",
		84181 => x"FF",
		84182 => x"FF",
		84183 => x"FF",
		84184 => x"FF",
		84185 => x"FF",
		84186 => x"FF",
		84187 => x"FF",
		84188 => x"FF",
		84189 => x"FF",
		84190 => x"FF",
		84191 => x"FF",
		84192 => x"FF",
		84193 => x"FF",
		84194 => x"FF",
		84195 => x"FF",
		84196 => x"FF",
		84197 => x"FF",
		84198 => x"FF",
		84199 => x"FF",
		84200 => x"FF",
		84201 => x"FF",
		84202 => x"FF",
		84203 => x"FF",
		84204 => x"FF",
		84205 => x"FF",
		84206 => x"FF",
		84207 => x"FF",
		84208 => x"FF",
		84209 => x"FF",
		84210 => x"FF",
		84211 => x"FF",
		84212 => x"FF",
		84213 => x"FF",
		84214 => x"FF",
		84215 => x"FF",
		84216 => x"FF",
		84217 => x"FF",
		84218 => x"FF",
		84219 => x"FF",
		84220 => x"FF",
		84221 => x"FF",
		84222 => x"FF",
		84223 => x"FF",
		84224 => x"FF",
		84225 => x"FF",
		84226 => x"FF",
		84227 => x"FF",
		84228 => x"FF",
		84229 => x"FF",
		84230 => x"FF",
		84231 => x"FF",
		84232 => x"FF",
		84233 => x"FF",
		84234 => x"FF",
		84235 => x"FF",
		84236 => x"FF",
		84237 => x"FF",
		84238 => x"FF",
		84239 => x"FF",
		84240 => x"FF",
		84241 => x"FF",
		85036 => x"FF",
		85037 => x"FF",
		85038 => x"FF",
		85039 => x"FF",
		85040 => x"FF",
		85041 => x"FF",
		85042 => x"FF",
		85043 => x"FF",
		85044 => x"FF",
		85045 => x"FF",
		85046 => x"FF",
		85047 => x"FF",
		85048 => x"FF",
		85049 => x"FF",
		85050 => x"FF",
		85051 => x"FF",
		85052 => x"FF",
		85053 => x"FF",
		85054 => x"FF",
		85055 => x"FF",
		85056 => x"FF",
		85057 => x"FF",
		85058 => x"FF",
		85059 => x"FF",
		85060 => x"FF",
		85061 => x"FF",
		85062 => x"FF",
		85063 => x"FF",
		85064 => x"FF",
		85065 => x"FF",
		85066 => x"FF",
		85067 => x"FF",
		85068 => x"FF",
		85069 => x"FF",
		85070 => x"FF",
		85071 => x"FF",
		85072 => x"FF",
		85073 => x"FF",
		85074 => x"FF",
		85075 => x"FF",
		85076 => x"FF",
		85077 => x"FF",
		85078 => x"FF",
		85079 => x"FF",
		85080 => x"FF",
		85081 => x"FF",
		85082 => x"FF",
		85083 => x"FF",
		85084 => x"FF",
		85085 => x"FF",
		85086 => x"FF",
		85087 => x"FF",
		85088 => x"FF",
		85089 => x"FF",
		85090 => x"FF",
		85091 => x"FF",
		85092 => x"FF",
		85093 => x"FF",
		85094 => x"FF",
		85095 => x"FF",
		85096 => x"FF",
		85097 => x"FF",
		85098 => x"FF",
		85099 => x"FF",
		85100 => x"FF",
		85101 => x"FF",
		85102 => x"FF",
		85103 => x"FF",
		85104 => x"FF",
		85105 => x"FF",
		85106 => x"FF",
		85107 => x"FF",
		85108 => x"FF",
		85109 => x"FF",
		85110 => x"FF",
		85111 => x"FF",
		85112 => x"FF",
		85113 => x"FF",
		85114 => x"FF",
		85115 => x"FF",
		85116 => x"FF",
		85117 => x"FF",
		85118 => x"FF",
		85119 => x"FF",
		85120 => x"FF",
		85121 => x"FF",
		85122 => x"FF",
		85123 => x"FF",
		85124 => x"FF",
		85125 => x"FF",
		85126 => x"FF",
		85127 => x"FF",
		85128 => x"FF",
		85129 => x"FF",
		85130 => x"FF",
		85131 => x"FF",
		85132 => x"FF",
		85133 => x"FF",
		85134 => x"FF",
		85135 => x"FF",
		85136 => x"FF",
		85137 => x"FF",
		85138 => x"FF",
		85139 => x"FF",
		85140 => x"FF",
		85141 => x"FF",
		85142 => x"FF",
		85143 => x"FF",
		85144 => x"FF",
		85145 => x"FF",
		85146 => x"FF",
		85147 => x"FF",
		85148 => x"FF",
		85149 => x"FF",
		85150 => x"FF",
		85151 => x"FF",
		85152 => x"FF",
		85153 => x"FF",
		85154 => x"FF",
		85155 => x"FF",
		85156 => x"FF",
		85157 => x"FF",
		85158 => x"FF",
		85159 => x"FF",
		85160 => x"FF",
		85161 => x"FF",
		85162 => x"FF",
		85163 => x"FF",
		85164 => x"FF",
		85165 => x"FF",
		85166 => x"FF",
		85167 => x"FF",
		85168 => x"FF",
		85169 => x"FF",
		85170 => x"FF",
		85171 => x"FF",
		85172 => x"FF",
		85173 => x"FF",
		85174 => x"FF",
		85175 => x"FF",
		85176 => x"FF",
		85177 => x"FF",
		85178 => x"FF",
		85179 => x"FF",
		85180 => x"FF",
		85181 => x"FF",
		85182 => x"FF",
		85183 => x"FF",
		85184 => x"FF",
		85185 => x"FF",
		85186 => x"FF",
		85187 => x"FF",
		85188 => x"FF",
		85189 => x"FF",
		85190 => x"FF",
		85191 => x"FF",
		85192 => x"FF",
		85193 => x"FF",
		85194 => x"FF",
		85195 => x"FF",
		85196 => x"FF",
		85197 => x"FF",
		85198 => x"FF",
		85199 => x"FF",
		85200 => x"FF",
		85201 => x"FF",
		85202 => x"FF",
		85203 => x"FF",
		85204 => x"FF",
		85205 => x"FF",
		85206 => x"FF",
		85207 => x"FF",
		85208 => x"FF",
		85209 => x"FF",
		85210 => x"FF",
		85211 => x"FF",
		85212 => x"FF",
		85213 => x"FF",
		85214 => x"FF",
		85215 => x"FF",
		85216 => x"FF",
		85217 => x"FF",
		85218 => x"FF",
		85219 => x"FF",
		85220 => x"FF",
		85221 => x"FF",
		85222 => x"FF",
		85223 => x"FF",
		85224 => x"FF",
		85225 => x"FF",
		85226 => x"FF",
		85227 => x"FF",
		85228 => x"FF",
		85229 => x"FF",
		85230 => x"FF",
		85231 => x"FF",
		85232 => x"FF",
		85233 => x"FF",
		85234 => x"FF",
		85235 => x"FF",
		85236 => x"FF",
		85237 => x"FF",
		85238 => x"FF",
		85239 => x"FF",
		85240 => x"FF",
		85241 => x"FF",
		85242 => x"FF",
		85243 => x"FF",
		85244 => x"FF",
		85245 => x"FF",
		85246 => x"FF",
		85247 => x"FF",
		85248 => x"FF",
		85249 => x"FF",
		85250 => x"FF",
		85251 => x"FF",
		85252 => x"FF",
		85253 => x"FF",
		85254 => x"FF",
		85255 => x"FF",
		85256 => x"FF",
		85257 => x"FF",
		85258 => x"FF",
		85259 => x"FF",
		85260 => x"FF",
		85261 => x"FF",
		85262 => x"FF",
		85263 => x"FF",
		85264 => x"FF",
		85265 => x"FF",
		86060 => x"FF",
		86061 => x"FF",
		86062 => x"FF",
		86063 => x"FF",
		86064 => x"FF",
		86135 => x"FF",
		86136 => x"FF",
		86137 => x"FF",
		86138 => x"FF",
		86139 => x"FF",
		86210 => x"FF",
		86211 => x"FF",
		86212 => x"FF",
		86213 => x"FF",
		86214 => x"FF",
		86285 => x"FF",
		86286 => x"FF",
		86287 => x"FF",
		86288 => x"FF",
		86289 => x"FF",
		87084 => x"FF",
		87085 => x"FF",
		87086 => x"FF",
		87087 => x"FF",
		87088 => x"FF",
		87159 => x"FF",
		87160 => x"FF",
		87161 => x"FF",
		87162 => x"FF",
		87163 => x"FF",
		87234 => x"FF",
		87235 => x"FF",
		87236 => x"FF",
		87237 => x"FF",
		87238 => x"FF",
		87309 => x"FF",
		87310 => x"FF",
		87311 => x"FF",
		87312 => x"FF",
		87313 => x"FF",
		88108 => x"FF",
		88109 => x"FF",
		88110 => x"FF",
		88111 => x"FF",
		88112 => x"FF",
		88183 => x"FF",
		88184 => x"FF",
		88185 => x"FF",
		88186 => x"FF",
		88187 => x"FF",
		88258 => x"FF",
		88259 => x"FF",
		88260 => x"FF",
		88261 => x"FF",
		88262 => x"FF",
		88333 => x"FF",
		88334 => x"FF",
		88335 => x"FF",
		88336 => x"FF",
		88337 => x"FF",
		89132 => x"FF",
		89133 => x"FF",
		89134 => x"FF",
		89135 => x"FF",
		89136 => x"FF",
		89207 => x"FF",
		89208 => x"FF",
		89209 => x"FF",
		89210 => x"FF",
		89211 => x"FF",
		89282 => x"FF",
		89283 => x"FF",
		89284 => x"FF",
		89285 => x"FF",
		89286 => x"FF",
		89357 => x"FF",
		89358 => x"FF",
		89359 => x"FF",
		89360 => x"FF",
		89361 => x"FF",
		90156 => x"FF",
		90157 => x"FF",
		90158 => x"FF",
		90159 => x"FF",
		90160 => x"FF",
		90231 => x"FF",
		90232 => x"FF",
		90233 => x"FF",
		90234 => x"FF",
		90235 => x"FF",
		90306 => x"FF",
		90307 => x"FF",
		90308 => x"FF",
		90309 => x"FF",
		90310 => x"FF",
		90381 => x"FF",
		90382 => x"FF",
		90383 => x"FF",
		90384 => x"FF",
		90385 => x"FF",
		91180 => x"FF",
		91181 => x"FF",
		91182 => x"FF",
		91183 => x"FF",
		91184 => x"FF",
		91255 => x"FF",
		91256 => x"FF",
		91257 => x"FF",
		91258 => x"FF",
		91259 => x"FF",
		91330 => x"FF",
		91331 => x"FF",
		91332 => x"FF",
		91333 => x"FF",
		91334 => x"FF",
		91405 => x"FF",
		91406 => x"FF",
		91407 => x"FF",
		91408 => x"FF",
		91409 => x"FF",
		92204 => x"FF",
		92205 => x"FF",
		92206 => x"FF",
		92207 => x"FF",
		92208 => x"FF",
		92279 => x"FF",
		92280 => x"FF",
		92281 => x"FF",
		92282 => x"FF",
		92283 => x"FF",
		92354 => x"FF",
		92355 => x"FF",
		92356 => x"FF",
		92357 => x"FF",
		92358 => x"FF",
		92429 => x"FF",
		92430 => x"FF",
		92431 => x"FF",
		92432 => x"FF",
		92433 => x"FF",
		93228 => x"FF",
		93229 => x"FF",
		93230 => x"FF",
		93231 => x"FF",
		93232 => x"FF",
		93303 => x"FF",
		93304 => x"FF",
		93305 => x"FF",
		93306 => x"FF",
		93307 => x"FF",
		93378 => x"FF",
		93379 => x"FF",
		93380 => x"FF",
		93381 => x"FF",
		93382 => x"FF",
		93453 => x"FF",
		93454 => x"FF",
		93455 => x"FF",
		93456 => x"FF",
		93457 => x"FF",
		94252 => x"FF",
		94253 => x"FF",
		94254 => x"FF",
		94255 => x"FF",
		94256 => x"FF",
		94327 => x"FF",
		94328 => x"FF",
		94329 => x"FF",
		94330 => x"FF",
		94331 => x"FF",
		94402 => x"FF",
		94403 => x"FF",
		94404 => x"FF",
		94405 => x"FF",
		94406 => x"FF",
		94477 => x"FF",
		94478 => x"FF",
		94479 => x"FF",
		94480 => x"FF",
		94481 => x"FF",
		95276 => x"FF",
		95277 => x"FF",
		95278 => x"FF",
		95279 => x"FF",
		95280 => x"FF",
		95351 => x"FF",
		95352 => x"FF",
		95353 => x"FF",
		95354 => x"FF",
		95355 => x"FF",
		95426 => x"FF",
		95427 => x"FF",
		95428 => x"FF",
		95429 => x"FF",
		95430 => x"FF",
		95501 => x"FF",
		95502 => x"FF",
		95503 => x"FF",
		95504 => x"FF",
		95505 => x"FF",
		96300 => x"FF",
		96301 => x"FF",
		96302 => x"FF",
		96303 => x"FF",
		96304 => x"FF",
		96375 => x"FF",
		96376 => x"FF",
		96377 => x"FF",
		96378 => x"FF",
		96379 => x"FF",
		96450 => x"FF",
		96451 => x"FF",
		96452 => x"FF",
		96453 => x"FF",
		96454 => x"FF",
		96525 => x"FF",
		96526 => x"FF",
		96527 => x"FF",
		96528 => x"FF",
		96529 => x"FF",
		97324 => x"FF",
		97325 => x"FF",
		97326 => x"FF",
		97327 => x"FF",
		97328 => x"FF",
		97399 => x"FF",
		97400 => x"FF",
		97401 => x"FF",
		97402 => x"FF",
		97403 => x"FF",
		97474 => x"FF",
		97475 => x"FF",
		97476 => x"FF",
		97477 => x"FF",
		97478 => x"FF",
		97549 => x"FF",
		97550 => x"FF",
		97551 => x"FF",
		97552 => x"FF",
		97553 => x"FF",
		98348 => x"FF",
		98349 => x"FF",
		98350 => x"FF",
		98351 => x"FF",
		98352 => x"FF",
		98423 => x"FF",
		98424 => x"FF",
		98425 => x"FF",
		98426 => x"FF",
		98427 => x"FF",
		98498 => x"FF",
		98499 => x"FF",
		98500 => x"FF",
		98501 => x"FF",
		98502 => x"FF",
		98573 => x"FF",
		98574 => x"FF",
		98575 => x"FF",
		98576 => x"FF",
		98577 => x"FF",
		99372 => x"FF",
		99373 => x"FF",
		99374 => x"FF",
		99375 => x"FF",
		99376 => x"FF",
		99447 => x"FF",
		99448 => x"FF",
		99449 => x"FF",
		99450 => x"FF",
		99451 => x"FF",
		99522 => x"FF",
		99523 => x"FF",
		99524 => x"FF",
		99525 => x"FF",
		99526 => x"FF",
		99597 => x"FF",
		99598 => x"FF",
		99599 => x"FF",
		99600 => x"FF",
		99601 => x"FF",
		100396 => x"FF",
		100397 => x"FF",
		100398 => x"FF",
		100399 => x"FF",
		100400 => x"FF",
		100471 => x"FF",
		100472 => x"FF",
		100473 => x"FF",
		100474 => x"FF",
		100475 => x"FF",
		100546 => x"FF",
		100547 => x"FF",
		100548 => x"FF",
		100549 => x"FF",
		100550 => x"FF",
		100621 => x"FF",
		100622 => x"FF",
		100623 => x"FF",
		100624 => x"FF",
		100625 => x"FF",
		101420 => x"FF",
		101421 => x"FF",
		101422 => x"FF",
		101423 => x"FF",
		101424 => x"FF",
		101495 => x"FF",
		101496 => x"FF",
		101497 => x"FF",
		101498 => x"FF",
		101499 => x"FF",
		101570 => x"FF",
		101571 => x"FF",
		101572 => x"FF",
		101573 => x"FF",
		101574 => x"FF",
		101645 => x"FF",
		101646 => x"FF",
		101647 => x"FF",
		101648 => x"FF",
		101649 => x"FF",
		102444 => x"FF",
		102445 => x"FF",
		102446 => x"FF",
		102447 => x"FF",
		102448 => x"FF",
		102519 => x"FF",
		102520 => x"FF",
		102521 => x"FF",
		102522 => x"FF",
		102523 => x"FF",
		102594 => x"FF",
		102595 => x"FF",
		102596 => x"FF",
		102597 => x"FF",
		102598 => x"FF",
		102669 => x"FF",
		102670 => x"FF",
		102671 => x"FF",
		102672 => x"FF",
		102673 => x"FF",
		103468 => x"FF",
		103469 => x"FF",
		103470 => x"FF",
		103471 => x"FF",
		103472 => x"FF",
		103543 => x"FF",
		103544 => x"FF",
		103545 => x"FF",
		103546 => x"FF",
		103547 => x"FF",
		103618 => x"FF",
		103619 => x"FF",
		103620 => x"FF",
		103621 => x"FF",
		103622 => x"FF",
		103693 => x"FF",
		103694 => x"FF",
		103695 => x"FF",
		103696 => x"FF",
		103697 => x"FF",
		104492 => x"FF",
		104493 => x"FF",
		104494 => x"FF",
		104495 => x"FF",
		104496 => x"FF",
		104567 => x"FF",
		104568 => x"FF",
		104569 => x"FF",
		104570 => x"FF",
		104571 => x"FF",
		104642 => x"FF",
		104643 => x"FF",
		104644 => x"FF",
		104645 => x"FF",
		104646 => x"FF",
		104717 => x"FF",
		104718 => x"FF",
		104719 => x"FF",
		104720 => x"FF",
		104721 => x"FF",
		105516 => x"FF",
		105517 => x"FF",
		105518 => x"FF",
		105519 => x"FF",
		105520 => x"FF",
		105591 => x"FF",
		105592 => x"FF",
		105593 => x"FF",
		105594 => x"FF",
		105595 => x"FF",
		105666 => x"FF",
		105667 => x"FF",
		105668 => x"FF",
		105669 => x"FF",
		105670 => x"FF",
		105741 => x"FF",
		105742 => x"FF",
		105743 => x"FF",
		105744 => x"FF",
		105745 => x"FF",
		106540 => x"FF",
		106541 => x"FF",
		106542 => x"FF",
		106543 => x"FF",
		106544 => x"FF",
		106615 => x"FF",
		106616 => x"FF",
		106617 => x"FF",
		106618 => x"FF",
		106619 => x"FF",
		106690 => x"FF",
		106691 => x"FF",
		106692 => x"FF",
		106693 => x"FF",
		106694 => x"FF",
		106765 => x"FF",
		106766 => x"FF",
		106767 => x"FF",
		106768 => x"FF",
		106769 => x"FF",
		107564 => x"FF",
		107565 => x"FF",
		107566 => x"FF",
		107567 => x"FF",
		107568 => x"FF",
		107639 => x"FF",
		107640 => x"FF",
		107641 => x"FF",
		107642 => x"FF",
		107643 => x"FF",
		107714 => x"FF",
		107715 => x"FF",
		107716 => x"FF",
		107717 => x"FF",
		107718 => x"FF",
		107789 => x"FF",
		107790 => x"FF",
		107791 => x"FF",
		107792 => x"FF",
		107793 => x"FF",
		108588 => x"FF",
		108589 => x"FF",
		108590 => x"FF",
		108591 => x"FF",
		108592 => x"FF",
		108663 => x"FF",
		108664 => x"FF",
		108665 => x"FF",
		108666 => x"FF",
		108667 => x"FF",
		108738 => x"FF",
		108739 => x"FF",
		108740 => x"FF",
		108741 => x"FF",
		108742 => x"FF",
		108813 => x"FF",
		108814 => x"FF",
		108815 => x"FF",
		108816 => x"FF",
		108817 => x"FF",
		109612 => x"FF",
		109613 => x"FF",
		109614 => x"FF",
		109615 => x"FF",
		109616 => x"FF",
		109687 => x"FF",
		109688 => x"FF",
		109689 => x"FF",
		109690 => x"FF",
		109691 => x"FF",
		109762 => x"FF",
		109763 => x"FF",
		109764 => x"FF",
		109765 => x"FF",
		109766 => x"FF",
		109837 => x"FF",
		109838 => x"FF",
		109839 => x"FF",
		109840 => x"FF",
		109841 => x"FF",
		110636 => x"FF",
		110637 => x"FF",
		110638 => x"FF",
		110639 => x"FF",
		110640 => x"FF",
		110711 => x"FF",
		110712 => x"FF",
		110713 => x"FF",
		110714 => x"FF",
		110715 => x"FF",
		110786 => x"FF",
		110787 => x"FF",
		110788 => x"FF",
		110789 => x"FF",
		110790 => x"FF",
		110861 => x"FF",
		110862 => x"FF",
		110863 => x"FF",
		110864 => x"FF",
		110865 => x"FF",
		111660 => x"FF",
		111661 => x"FF",
		111662 => x"FF",
		111663 => x"FF",
		111664 => x"FF",
		111735 => x"FF",
		111736 => x"FF",
		111737 => x"FF",
		111738 => x"FF",
		111739 => x"FF",
		111810 => x"FF",
		111811 => x"FF",
		111812 => x"FF",
		111813 => x"FF",
		111814 => x"FF",
		111885 => x"FF",
		111886 => x"FF",
		111887 => x"FF",
		111888 => x"FF",
		111889 => x"FF",
		112684 => x"FF",
		112685 => x"FF",
		112686 => x"FF",
		112687 => x"FF",
		112688 => x"FF",
		112759 => x"FF",
		112760 => x"FF",
		112761 => x"FF",
		112762 => x"FF",
		112763 => x"FF",
		112834 => x"FF",
		112835 => x"FF",
		112836 => x"FF",
		112837 => x"FF",
		112838 => x"FF",
		112909 => x"FF",
		112910 => x"FF",
		112911 => x"FF",
		112912 => x"FF",
		112913 => x"FF",
		113708 => x"FF",
		113709 => x"FF",
		113710 => x"FF",
		113711 => x"FF",
		113712 => x"FF",
		113783 => x"FF",
		113784 => x"FF",
		113785 => x"FF",
		113786 => x"FF",
		113787 => x"FF",
		113858 => x"FF",
		113859 => x"FF",
		113860 => x"FF",
		113861 => x"FF",
		113862 => x"FF",
		113933 => x"FF",
		113934 => x"FF",
		113935 => x"FF",
		113936 => x"FF",
		113937 => x"FF",
		114732 => x"FF",
		114733 => x"FF",
		114734 => x"FF",
		114735 => x"FF",
		114736 => x"FF",
		114807 => x"FF",
		114808 => x"FF",
		114809 => x"FF",
		114810 => x"FF",
		114811 => x"FF",
		114882 => x"FF",
		114883 => x"FF",
		114884 => x"FF",
		114885 => x"FF",
		114886 => x"FF",
		114957 => x"FF",
		114958 => x"FF",
		114959 => x"FF",
		114960 => x"FF",
		114961 => x"FF",
		115756 => x"FF",
		115757 => x"FF",
		115758 => x"FF",
		115759 => x"FF",
		115760 => x"FF",
		115831 => x"FF",
		115832 => x"FF",
		115833 => x"FF",
		115834 => x"FF",
		115835 => x"FF",
		115906 => x"FF",
		115907 => x"FF",
		115908 => x"FF",
		115909 => x"FF",
		115910 => x"FF",
		115981 => x"FF",
		115982 => x"FF",
		115983 => x"FF",
		115984 => x"FF",
		115985 => x"FF",
		116780 => x"FF",
		116781 => x"FF",
		116782 => x"FF",
		116783 => x"FF",
		116784 => x"FF",
		116855 => x"FF",
		116856 => x"FF",
		116857 => x"FF",
		116858 => x"FF",
		116859 => x"FF",
		116930 => x"FF",
		116931 => x"FF",
		116932 => x"FF",
		116933 => x"FF",
		116934 => x"FF",
		117005 => x"FF",
		117006 => x"FF",
		117007 => x"FF",
		117008 => x"FF",
		117009 => x"FF",
		117804 => x"FF",
		117805 => x"FF",
		117806 => x"FF",
		117807 => x"FF",
		117808 => x"FF",
		117879 => x"FF",
		117880 => x"FF",
		117881 => x"FF",
		117882 => x"FF",
		117883 => x"FF",
		117954 => x"FF",
		117955 => x"FF",
		117956 => x"FF",
		117957 => x"FF",
		117958 => x"FF",
		118029 => x"FF",
		118030 => x"FF",
		118031 => x"FF",
		118032 => x"FF",
		118033 => x"FF",
		118828 => x"FF",
		118829 => x"FF",
		118830 => x"FF",
		118831 => x"FF",
		118832 => x"FF",
		118903 => x"FF",
		118904 => x"FF",
		118905 => x"FF",
		118906 => x"FF",
		118907 => x"FF",
		118978 => x"FF",
		118979 => x"FF",
		118980 => x"FF",
		118981 => x"FF",
		118982 => x"FF",
		119053 => x"FF",
		119054 => x"FF",
		119055 => x"FF",
		119056 => x"FF",
		119057 => x"FF",
		119852 => x"FF",
		119853 => x"FF",
		119854 => x"FF",
		119855 => x"FF",
		119856 => x"FF",
		119927 => x"FF",
		119928 => x"FF",
		119929 => x"FF",
		119930 => x"FF",
		119931 => x"FF",
		120002 => x"FF",
		120003 => x"FF",
		120004 => x"FF",
		120005 => x"FF",
		120006 => x"FF",
		120077 => x"FF",
		120078 => x"FF",
		120079 => x"FF",
		120080 => x"FF",
		120081 => x"FF",
		120876 => x"FF",
		120877 => x"FF",
		120878 => x"FF",
		120879 => x"FF",
		120880 => x"FF",
		120951 => x"FF",
		120952 => x"FF",
		120953 => x"FF",
		120954 => x"FF",
		120955 => x"FF",
		121026 => x"FF",
		121027 => x"FF",
		121028 => x"FF",
		121029 => x"FF",
		121030 => x"FF",
		121101 => x"FF",
		121102 => x"FF",
		121103 => x"FF",
		121104 => x"FF",
		121105 => x"FF",
		121900 => x"FF",
		121901 => x"FF",
		121902 => x"FF",
		121903 => x"FF",
		121904 => x"FF",
		121975 => x"FF",
		121976 => x"FF",
		121977 => x"FF",
		121978 => x"FF",
		121979 => x"FF",
		122050 => x"FF",
		122051 => x"FF",
		122052 => x"FF",
		122053 => x"FF",
		122054 => x"FF",
		122125 => x"FF",
		122126 => x"FF",
		122127 => x"FF",
		122128 => x"FF",
		122129 => x"FF",
		122924 => x"FF",
		122925 => x"FF",
		122926 => x"FF",
		122927 => x"FF",
		122928 => x"FF",
		122999 => x"FF",
		123000 => x"FF",
		123001 => x"FF",
		123002 => x"FF",
		123003 => x"FF",
		123074 => x"FF",
		123075 => x"FF",
		123076 => x"FF",
		123077 => x"FF",
		123078 => x"FF",
		123149 => x"FF",
		123150 => x"FF",
		123151 => x"FF",
		123152 => x"FF",
		123153 => x"FF",
		123948 => x"FF",
		123949 => x"FF",
		123950 => x"FF",
		123951 => x"FF",
		123952 => x"FF",
		124023 => x"FF",
		124024 => x"FF",
		124025 => x"FF",
		124026 => x"FF",
		124027 => x"FF",
		124098 => x"FF",
		124099 => x"FF",
		124100 => x"FF",
		124101 => x"FF",
		124102 => x"FF",
		124173 => x"FF",
		124174 => x"FF",
		124175 => x"FF",
		124176 => x"FF",
		124177 => x"FF",
		124972 => x"FF",
		124973 => x"FF",
		124974 => x"FF",
		124975 => x"FF",
		124976 => x"FF",
		125047 => x"FF",
		125048 => x"FF",
		125049 => x"FF",
		125050 => x"FF",
		125051 => x"FF",
		125122 => x"FF",
		125123 => x"FF",
		125124 => x"FF",
		125125 => x"FF",
		125126 => x"FF",
		125197 => x"FF",
		125198 => x"FF",
		125199 => x"FF",
		125200 => x"FF",
		125201 => x"FF",
		125996 => x"FF",
		125997 => x"FF",
		125998 => x"FF",
		125999 => x"FF",
		126000 => x"FF",
		126071 => x"FF",
		126072 => x"FF",
		126073 => x"FF",
		126074 => x"FF",
		126075 => x"FF",
		126146 => x"FF",
		126147 => x"FF",
		126148 => x"FF",
		126149 => x"FF",
		126150 => x"FF",
		126221 => x"FF",
		126222 => x"FF",
		126223 => x"FF",
		126224 => x"FF",
		126225 => x"FF",
		127020 => x"FF",
		127021 => x"FF",
		127022 => x"FF",
		127023 => x"FF",
		127024 => x"FF",
		127095 => x"FF",
		127096 => x"FF",
		127097 => x"FF",
		127098 => x"FF",
		127099 => x"FF",
		127170 => x"FF",
		127171 => x"FF",
		127172 => x"FF",
		127173 => x"FF",
		127174 => x"FF",
		127245 => x"FF",
		127246 => x"FF",
		127247 => x"FF",
		127248 => x"FF",
		127249 => x"FF",
		128044 => x"FF",
		128045 => x"FF",
		128046 => x"FF",
		128047 => x"FF",
		128048 => x"FF",
		128119 => x"FF",
		128120 => x"FF",
		128121 => x"FF",
		128122 => x"FF",
		128123 => x"FF",
		128194 => x"FF",
		128195 => x"FF",
		128196 => x"FF",
		128197 => x"FF",
		128198 => x"FF",
		128269 => x"FF",
		128270 => x"FF",
		128271 => x"FF",
		128272 => x"FF",
		128273 => x"FF",
		129068 => x"FF",
		129069 => x"FF",
		129070 => x"FF",
		129071 => x"FF",
		129072 => x"FF",
		129143 => x"FF",
		129144 => x"FF",
		129145 => x"FF",
		129146 => x"FF",
		129147 => x"FF",
		129218 => x"FF",
		129219 => x"FF",
		129220 => x"FF",
		129221 => x"FF",
		129222 => x"FF",
		129293 => x"FF",
		129294 => x"FF",
		129295 => x"FF",
		129296 => x"FF",
		129297 => x"FF",
		130092 => x"FF",
		130093 => x"FF",
		130094 => x"FF",
		130095 => x"FF",
		130096 => x"FF",
		130167 => x"FF",
		130168 => x"FF",
		130169 => x"FF",
		130170 => x"FF",
		130171 => x"FF",
		130242 => x"FF",
		130243 => x"FF",
		130244 => x"FF",
		130245 => x"FF",
		130246 => x"FF",
		130317 => x"FF",
		130318 => x"FF",
		130319 => x"FF",
		130320 => x"FF",
		130321 => x"FF",
		131116 => x"FF",
		131117 => x"FF",
		131118 => x"FF",
		131119 => x"FF",
		131120 => x"FF",
		131191 => x"FF",
		131192 => x"FF",
		131193 => x"FF",
		131194 => x"FF",
		131195 => x"FF",
		131266 => x"FF",
		131267 => x"FF",
		131268 => x"FF",
		131269 => x"FF",
		131270 => x"FF",
		131341 => x"FF",
		131342 => x"FF",
		131343 => x"FF",
		131344 => x"FF",
		131345 => x"FF",
		132140 => x"FF",
		132141 => x"FF",
		132142 => x"FF",
		132143 => x"FF",
		132144 => x"FF",
		132215 => x"FF",
		132216 => x"FF",
		132217 => x"FF",
		132218 => x"FF",
		132219 => x"FF",
		132290 => x"FF",
		132291 => x"FF",
		132292 => x"FF",
		132293 => x"FF",
		132294 => x"FF",
		132365 => x"FF",
		132366 => x"FF",
		132367 => x"FF",
		132368 => x"FF",
		132369 => x"FF",
		133164 => x"FF",
		133165 => x"FF",
		133166 => x"FF",
		133167 => x"FF",
		133168 => x"FF",
		133239 => x"FF",
		133240 => x"FF",
		133241 => x"FF",
		133242 => x"FF",
		133243 => x"FF",
		133314 => x"FF",
		133315 => x"FF",
		133316 => x"FF",
		133317 => x"FF",
		133318 => x"FF",
		133389 => x"FF",
		133390 => x"FF",
		133391 => x"FF",
		133392 => x"FF",
		133393 => x"FF",
		134188 => x"FF",
		134189 => x"FF",
		134190 => x"FF",
		134191 => x"FF",
		134192 => x"FF",
		134263 => x"FF",
		134264 => x"FF",
		134265 => x"FF",
		134266 => x"FF",
		134267 => x"FF",
		134338 => x"FF",
		134339 => x"FF",
		134340 => x"FF",
		134341 => x"FF",
		134342 => x"FF",
		134413 => x"FF",
		134414 => x"FF",
		134415 => x"FF",
		134416 => x"FF",
		134417 => x"FF",
		135212 => x"FF",
		135213 => x"FF",
		135214 => x"FF",
		135215 => x"FF",
		135216 => x"FF",
		135287 => x"FF",
		135288 => x"FF",
		135289 => x"FF",
		135290 => x"FF",
		135291 => x"FF",
		135362 => x"FF",
		135363 => x"FF",
		135364 => x"FF",
		135365 => x"FF",
		135366 => x"FF",
		135437 => x"FF",
		135438 => x"FF",
		135439 => x"FF",
		135440 => x"FF",
		135441 => x"FF",
		136236 => x"FF",
		136237 => x"FF",
		136238 => x"FF",
		136239 => x"FF",
		136240 => x"FF",
		136311 => x"FF",
		136312 => x"FF",
		136313 => x"FF",
		136314 => x"FF",
		136315 => x"FF",
		136386 => x"FF",
		136387 => x"FF",
		136388 => x"FF",
		136389 => x"FF",
		136390 => x"FF",
		136461 => x"FF",
		136462 => x"FF",
		136463 => x"FF",
		136464 => x"FF",
		136465 => x"FF",
		137260 => x"FF",
		137261 => x"FF",
		137262 => x"FF",
		137263 => x"FF",
		137264 => x"FF",
		137335 => x"FF",
		137336 => x"FF",
		137337 => x"FF",
		137338 => x"FF",
		137339 => x"FF",
		137410 => x"FF",
		137411 => x"FF",
		137412 => x"FF",
		137413 => x"FF",
		137414 => x"FF",
		137485 => x"FF",
		137486 => x"FF",
		137487 => x"FF",
		137488 => x"FF",
		137489 => x"FF",
		138284 => x"FF",
		138285 => x"FF",
		138286 => x"FF",
		138287 => x"FF",
		138288 => x"FF",
		138359 => x"FF",
		138360 => x"FF",
		138361 => x"FF",
		138362 => x"FF",
		138363 => x"FF",
		138434 => x"FF",
		138435 => x"FF",
		138436 => x"FF",
		138437 => x"FF",
		138438 => x"FF",
		138509 => x"FF",
		138510 => x"FF",
		138511 => x"FF",
		138512 => x"FF",
		138513 => x"FF",
		139308 => x"FF",
		139309 => x"FF",
		139310 => x"FF",
		139311 => x"FF",
		139312 => x"FF",
		139383 => x"FF",
		139384 => x"FF",
		139385 => x"FF",
		139386 => x"FF",
		139387 => x"FF",
		139458 => x"FF",
		139459 => x"FF",
		139460 => x"FF",
		139461 => x"FF",
		139462 => x"FF",
		139533 => x"FF",
		139534 => x"FF",
		139535 => x"FF",
		139536 => x"FF",
		139537 => x"FF",
		140332 => x"FF",
		140333 => x"FF",
		140334 => x"FF",
		140335 => x"FF",
		140336 => x"FF",
		140407 => x"FF",
		140408 => x"FF",
		140409 => x"FF",
		140410 => x"FF",
		140411 => x"FF",
		140482 => x"FF",
		140483 => x"FF",
		140484 => x"FF",
		140485 => x"FF",
		140486 => x"FF",
		140557 => x"FF",
		140558 => x"FF",
		140559 => x"FF",
		140560 => x"FF",
		140561 => x"FF",
		141356 => x"FF",
		141357 => x"FF",
		141358 => x"FF",
		141359 => x"FF",
		141360 => x"FF",
		141431 => x"FF",
		141432 => x"FF",
		141433 => x"FF",
		141434 => x"FF",
		141435 => x"FF",
		141506 => x"FF",
		141507 => x"FF",
		141508 => x"FF",
		141509 => x"FF",
		141510 => x"FF",
		141581 => x"FF",
		141582 => x"FF",
		141583 => x"FF",
		141584 => x"FF",
		141585 => x"FF",
		142380 => x"FF",
		142381 => x"FF",
		142382 => x"FF",
		142383 => x"FF",
		142384 => x"FF",
		142455 => x"FF",
		142456 => x"FF",
		142457 => x"FF",
		142458 => x"FF",
		142459 => x"FF",
		142530 => x"FF",
		142531 => x"FF",
		142532 => x"FF",
		142533 => x"FF",
		142534 => x"FF",
		142605 => x"FF",
		142606 => x"FF",
		142607 => x"FF",
		142608 => x"FF",
		142609 => x"FF",
		143404 => x"FF",
		143405 => x"FF",
		143406 => x"FF",
		143407 => x"FF",
		143408 => x"FF",
		143479 => x"FF",
		143480 => x"FF",
		143481 => x"FF",
		143482 => x"FF",
		143483 => x"FF",
		143554 => x"FF",
		143555 => x"FF",
		143556 => x"FF",
		143557 => x"FF",
		143558 => x"FF",
		143629 => x"FF",
		143630 => x"FF",
		143631 => x"FF",
		143632 => x"FF",
		143633 => x"FF",
		144428 => x"FF",
		144429 => x"FF",
		144430 => x"FF",
		144431 => x"FF",
		144432 => x"FF",
		144503 => x"FF",
		144504 => x"FF",
		144505 => x"FF",
		144506 => x"FF",
		144507 => x"FF",
		144578 => x"FF",
		144579 => x"FF",
		144580 => x"FF",
		144581 => x"FF",
		144582 => x"FF",
		144653 => x"FF",
		144654 => x"FF",
		144655 => x"FF",
		144656 => x"FF",
		144657 => x"FF",
		145452 => x"FF",
		145453 => x"FF",
		145454 => x"FF",
		145455 => x"FF",
		145456 => x"FF",
		145527 => x"FF",
		145528 => x"FF",
		145529 => x"FF",
		145530 => x"FF",
		145531 => x"FF",
		145602 => x"FF",
		145603 => x"FF",
		145604 => x"FF",
		145605 => x"FF",
		145606 => x"FF",
		145677 => x"FF",
		145678 => x"FF",
		145679 => x"FF",
		145680 => x"FF",
		145681 => x"FF",
		146476 => x"FF",
		146477 => x"FF",
		146478 => x"FF",
		146479 => x"FF",
		146480 => x"FF",
		146551 => x"FF",
		146552 => x"FF",
		146553 => x"FF",
		146554 => x"FF",
		146555 => x"FF",
		146626 => x"FF",
		146627 => x"FF",
		146628 => x"FF",
		146629 => x"FF",
		146630 => x"FF",
		146701 => x"FF",
		146702 => x"FF",
		146703 => x"FF",
		146704 => x"FF",
		146705 => x"FF",
		147500 => x"FF",
		147501 => x"FF",
		147502 => x"FF",
		147503 => x"FF",
		147504 => x"FF",
		147575 => x"FF",
		147576 => x"FF",
		147577 => x"FF",
		147578 => x"FF",
		147579 => x"FF",
		147650 => x"FF",
		147651 => x"FF",
		147652 => x"FF",
		147653 => x"FF",
		147654 => x"FF",
		147725 => x"FF",
		147726 => x"FF",
		147727 => x"FF",
		147728 => x"FF",
		147729 => x"FF",
		148524 => x"FF",
		148525 => x"FF",
		148526 => x"FF",
		148527 => x"FF",
		148528 => x"FF",
		148599 => x"FF",
		148600 => x"FF",
		148601 => x"FF",
		148602 => x"FF",
		148603 => x"FF",
		148674 => x"FF",
		148675 => x"FF",
		148676 => x"FF",
		148677 => x"FF",
		148678 => x"FF",
		148749 => x"FF",
		148750 => x"FF",
		148751 => x"FF",
		148752 => x"FF",
		148753 => x"FF",
		149548 => x"FF",
		149549 => x"FF",
		149550 => x"FF",
		149551 => x"FF",
		149552 => x"FF",
		149623 => x"FF",
		149624 => x"FF",
		149625 => x"FF",
		149626 => x"FF",
		149627 => x"FF",
		149698 => x"FF",
		149699 => x"FF",
		149700 => x"FF",
		149701 => x"FF",
		149702 => x"FF",
		149773 => x"FF",
		149774 => x"FF",
		149775 => x"FF",
		149776 => x"FF",
		149777 => x"FF",
		150572 => x"FF",
		150573 => x"FF",
		150574 => x"FF",
		150575 => x"FF",
		150576 => x"FF",
		150647 => x"FF",
		150648 => x"FF",
		150649 => x"FF",
		150650 => x"FF",
		150651 => x"FF",
		150722 => x"FF",
		150723 => x"FF",
		150724 => x"FF",
		150725 => x"FF",
		150726 => x"FF",
		150797 => x"FF",
		150798 => x"FF",
		150799 => x"FF",
		150800 => x"FF",
		150801 => x"FF",
		151596 => x"FF",
		151597 => x"FF",
		151598 => x"FF",
		151599 => x"FF",
		151600 => x"FF",
		151671 => x"FF",
		151672 => x"FF",
		151673 => x"FF",
		151674 => x"FF",
		151675 => x"FF",
		151746 => x"FF",
		151747 => x"FF",
		151748 => x"FF",
		151749 => x"FF",
		151750 => x"FF",
		151821 => x"FF",
		151822 => x"FF",
		151823 => x"FF",
		151824 => x"FF",
		151825 => x"FF",
		152620 => x"FF",
		152621 => x"FF",
		152622 => x"FF",
		152623 => x"FF",
		152624 => x"FF",
		152695 => x"FF",
		152696 => x"FF",
		152697 => x"FF",
		152698 => x"FF",
		152699 => x"FF",
		152770 => x"FF",
		152771 => x"FF",
		152772 => x"FF",
		152773 => x"FF",
		152774 => x"FF",
		152845 => x"FF",
		152846 => x"FF",
		152847 => x"FF",
		152848 => x"FF",
		152849 => x"FF",
		153644 => x"FF",
		153645 => x"FF",
		153646 => x"FF",
		153647 => x"FF",
		153648 => x"FF",
		153719 => x"FF",
		153720 => x"FF",
		153721 => x"FF",
		153722 => x"FF",
		153723 => x"FF",
		153794 => x"FF",
		153795 => x"FF",
		153796 => x"FF",
		153797 => x"FF",
		153798 => x"FF",
		153869 => x"FF",
		153870 => x"FF",
		153871 => x"FF",
		153872 => x"FF",
		153873 => x"FF",
		154668 => x"FF",
		154669 => x"FF",
		154670 => x"FF",
		154671 => x"FF",
		154672 => x"FF",
		154743 => x"FF",
		154744 => x"FF",
		154745 => x"FF",
		154746 => x"FF",
		154747 => x"FF",
		154818 => x"FF",
		154819 => x"FF",
		154820 => x"FF",
		154821 => x"FF",
		154822 => x"FF",
		154893 => x"FF",
		154894 => x"FF",
		154895 => x"FF",
		154896 => x"FF",
		154897 => x"FF",
		155692 => x"FF",
		155693 => x"FF",
		155694 => x"FF",
		155695 => x"FF",
		155696 => x"FF",
		155767 => x"FF",
		155768 => x"FF",
		155769 => x"FF",
		155770 => x"FF",
		155771 => x"FF",
		155842 => x"FF",
		155843 => x"FF",
		155844 => x"FF",
		155845 => x"FF",
		155846 => x"FF",
		155917 => x"FF",
		155918 => x"FF",
		155919 => x"FF",
		155920 => x"FF",
		155921 => x"FF",
		156716 => x"FF",
		156717 => x"FF",
		156718 => x"FF",
		156719 => x"FF",
		156720 => x"FF",
		156791 => x"FF",
		156792 => x"FF",
		156793 => x"FF",
		156794 => x"FF",
		156795 => x"FF",
		156866 => x"FF",
		156867 => x"FF",
		156868 => x"FF",
		156869 => x"FF",
		156870 => x"FF",
		156941 => x"FF",
		156942 => x"FF",
		156943 => x"FF",
		156944 => x"FF",
		156945 => x"FF",
		157740 => x"FF",
		157741 => x"FF",
		157742 => x"FF",
		157743 => x"FF",
		157744 => x"FF",
		157745 => x"FF",
		157746 => x"FF",
		157747 => x"FF",
		157748 => x"FF",
		157749 => x"FF",
		157750 => x"FF",
		157751 => x"FF",
		157752 => x"FF",
		157753 => x"FF",
		157754 => x"FF",
		157755 => x"FF",
		157756 => x"FF",
		157757 => x"FF",
		157758 => x"FF",
		157759 => x"FF",
		157760 => x"FF",
		157761 => x"FF",
		157762 => x"FF",
		157763 => x"FF",
		157764 => x"FF",
		157765 => x"FF",
		157766 => x"FF",
		157767 => x"FF",
		157768 => x"FF",
		157769 => x"FF",
		157770 => x"FF",
		157771 => x"FF",
		157772 => x"FF",
		157773 => x"FF",
		157774 => x"FF",
		157775 => x"FF",
		157776 => x"FF",
		157777 => x"FF",
		157778 => x"FF",
		157779 => x"FF",
		157780 => x"FF",
		157781 => x"FF",
		157782 => x"FF",
		157783 => x"FF",
		157784 => x"FF",
		157785 => x"FF",
		157786 => x"FF",
		157787 => x"FF",
		157788 => x"FF",
		157789 => x"FF",
		157790 => x"FF",
		157791 => x"FF",
		157792 => x"FF",
		157793 => x"FF",
		157794 => x"FF",
		157795 => x"FF",
		157796 => x"FF",
		157797 => x"FF",
		157798 => x"FF",
		157799 => x"FF",
		157800 => x"FF",
		157801 => x"FF",
		157802 => x"FF",
		157803 => x"FF",
		157804 => x"FF",
		157805 => x"FF",
		157806 => x"FF",
		157807 => x"FF",
		157808 => x"FF",
		157809 => x"FF",
		157810 => x"FF",
		157811 => x"FF",
		157812 => x"FF",
		157813 => x"FF",
		157814 => x"FF",
		157815 => x"FF",
		157816 => x"FF",
		157817 => x"FF",
		157818 => x"FF",
		157819 => x"FF",
		157820 => x"FF",
		157821 => x"FF",
		157822 => x"FF",
		157823 => x"FF",
		157824 => x"FF",
		157825 => x"FF",
		157826 => x"FF",
		157827 => x"FF",
		157828 => x"FF",
		157829 => x"FF",
		157830 => x"FF",
		157831 => x"FF",
		157832 => x"FF",
		157833 => x"FF",
		157834 => x"FF",
		157835 => x"FF",
		157836 => x"FF",
		157837 => x"FF",
		157838 => x"FF",
		157839 => x"FF",
		157840 => x"FF",
		157841 => x"FF",
		157842 => x"FF",
		157843 => x"FF",
		157844 => x"FF",
		157845 => x"FF",
		157846 => x"FF",
		157847 => x"FF",
		157848 => x"FF",
		157849 => x"FF",
		157850 => x"FF",
		157851 => x"FF",
		157852 => x"FF",
		157853 => x"FF",
		157854 => x"FF",
		157855 => x"FF",
		157856 => x"FF",
		157857 => x"FF",
		157858 => x"FF",
		157859 => x"FF",
		157860 => x"FF",
		157861 => x"FF",
		157862 => x"FF",
		157863 => x"FF",
		157864 => x"FF",
		157865 => x"FF",
		157866 => x"FF",
		157867 => x"FF",
		157868 => x"FF",
		157869 => x"FF",
		157870 => x"FF",
		157871 => x"FF",
		157872 => x"FF",
		157873 => x"FF",
		157874 => x"FF",
		157875 => x"FF",
		157876 => x"FF",
		157877 => x"FF",
		157878 => x"FF",
		157879 => x"FF",
		157880 => x"FF",
		157881 => x"FF",
		157882 => x"FF",
		157883 => x"FF",
		157884 => x"FF",
		157885 => x"FF",
		157886 => x"FF",
		157887 => x"FF",
		157888 => x"FF",
		157889 => x"FF",
		157890 => x"FF",
		157891 => x"FF",
		157892 => x"FF",
		157893 => x"FF",
		157894 => x"FF",
		157895 => x"FF",
		157896 => x"FF",
		157897 => x"FF",
		157898 => x"FF",
		157899 => x"FF",
		157900 => x"FF",
		157901 => x"FF",
		157902 => x"FF",
		157903 => x"FF",
		157904 => x"FF",
		157905 => x"FF",
		157906 => x"FF",
		157907 => x"FF",
		157908 => x"FF",
		157909 => x"FF",
		157910 => x"FF",
		157911 => x"FF",
		157912 => x"FF",
		157913 => x"FF",
		157914 => x"FF",
		157915 => x"FF",
		157916 => x"FF",
		157917 => x"FF",
		157918 => x"FF",
		157919 => x"FF",
		157920 => x"FF",
		157921 => x"FF",
		157922 => x"FF",
		157923 => x"FF",
		157924 => x"FF",
		157925 => x"FF",
		157926 => x"FF",
		157927 => x"FF",
		157928 => x"FF",
		157929 => x"FF",
		157930 => x"FF",
		157931 => x"FF",
		157932 => x"FF",
		157933 => x"FF",
		157934 => x"FF",
		157935 => x"FF",
		157936 => x"FF",
		157937 => x"FF",
		157938 => x"FF",
		157939 => x"FF",
		157940 => x"FF",
		157941 => x"FF",
		157942 => x"FF",
		157943 => x"FF",
		157944 => x"FF",
		157945 => x"FF",
		157946 => x"FF",
		157947 => x"FF",
		157948 => x"FF",
		157949 => x"FF",
		157950 => x"FF",
		157951 => x"FF",
		157952 => x"FF",
		157953 => x"FF",
		157954 => x"FF",
		157955 => x"FF",
		157956 => x"FF",
		157957 => x"FF",
		157958 => x"FF",
		157959 => x"FF",
		157960 => x"FF",
		157961 => x"FF",
		157962 => x"FF",
		157963 => x"FF",
		157964 => x"FF",
		157965 => x"FF",
		157966 => x"FF",
		157967 => x"FF",
		157968 => x"FF",
		157969 => x"FF",
		158764 => x"FF",
		158765 => x"FF",
		158766 => x"FF",
		158767 => x"FF",
		158768 => x"FF",
		158769 => x"FF",
		158770 => x"FF",
		158771 => x"FF",
		158772 => x"FF",
		158773 => x"FF",
		158774 => x"FF",
		158775 => x"FF",
		158776 => x"FF",
		158777 => x"FF",
		158778 => x"FF",
		158779 => x"FF",
		158780 => x"FF",
		158781 => x"FF",
		158782 => x"FF",
		158783 => x"FF",
		158784 => x"FF",
		158785 => x"FF",
		158786 => x"FF",
		158787 => x"FF",
		158788 => x"FF",
		158789 => x"FF",
		158790 => x"FF",
		158791 => x"FF",
		158792 => x"FF",
		158793 => x"FF",
		158794 => x"FF",
		158795 => x"FF",
		158796 => x"FF",
		158797 => x"FF",
		158798 => x"FF",
		158799 => x"FF",
		158800 => x"FF",
		158801 => x"FF",
		158802 => x"FF",
		158803 => x"FF",
		158804 => x"FF",
		158805 => x"FF",
		158806 => x"FF",
		158807 => x"FF",
		158808 => x"FF",
		158809 => x"FF",
		158810 => x"FF",
		158811 => x"FF",
		158812 => x"FF",
		158813 => x"FF",
		158814 => x"FF",
		158815 => x"FF",
		158816 => x"FF",
		158817 => x"FF",
		158818 => x"FF",
		158819 => x"FF",
		158820 => x"FF",
		158821 => x"FF",
		158822 => x"FF",
		158823 => x"FF",
		158824 => x"FF",
		158825 => x"FF",
		158826 => x"FF",
		158827 => x"FF",
		158828 => x"FF",
		158829 => x"FF",
		158830 => x"FF",
		158831 => x"FF",
		158832 => x"FF",
		158833 => x"FF",
		158834 => x"FF",
		158835 => x"FF",
		158836 => x"FF",
		158837 => x"FF",
		158838 => x"FF",
		158839 => x"FF",
		158840 => x"FF",
		158841 => x"FF",
		158842 => x"FF",
		158843 => x"FF",
		158844 => x"FF",
		158845 => x"FF",
		158846 => x"FF",
		158847 => x"FF",
		158848 => x"FF",
		158849 => x"FF",
		158850 => x"FF",
		158851 => x"FF",
		158852 => x"FF",
		158853 => x"FF",
		158854 => x"FF",
		158855 => x"FF",
		158856 => x"FF",
		158857 => x"FF",
		158858 => x"FF",
		158859 => x"FF",
		158860 => x"FF",
		158861 => x"FF",
		158862 => x"FF",
		158863 => x"FF",
		158864 => x"FF",
		158865 => x"FF",
		158866 => x"FF",
		158867 => x"FF",
		158868 => x"FF",
		158869 => x"FF",
		158870 => x"FF",
		158871 => x"FF",
		158872 => x"FF",
		158873 => x"FF",
		158874 => x"FF",
		158875 => x"FF",
		158876 => x"FF",
		158877 => x"FF",
		158878 => x"FF",
		158879 => x"FF",
		158880 => x"FF",
		158881 => x"FF",
		158882 => x"FF",
		158883 => x"FF",
		158884 => x"FF",
		158885 => x"FF",
		158886 => x"FF",
		158887 => x"FF",
		158888 => x"FF",
		158889 => x"FF",
		158890 => x"FF",
		158891 => x"FF",
		158892 => x"FF",
		158893 => x"FF",
		158894 => x"FF",
		158895 => x"FF",
		158896 => x"FF",
		158897 => x"FF",
		158898 => x"FF",
		158899 => x"FF",
		158900 => x"FF",
		158901 => x"FF",
		158902 => x"FF",
		158903 => x"FF",
		158904 => x"FF",
		158905 => x"FF",
		158906 => x"FF",
		158907 => x"FF",
		158908 => x"FF",
		158909 => x"FF",
		158910 => x"FF",
		158911 => x"FF",
		158912 => x"FF",
		158913 => x"FF",
		158914 => x"FF",
		158915 => x"FF",
		158916 => x"FF",
		158917 => x"FF",
		158918 => x"FF",
		158919 => x"FF",
		158920 => x"FF",
		158921 => x"FF",
		158922 => x"FF",
		158923 => x"FF",
		158924 => x"FF",
		158925 => x"FF",
		158926 => x"FF",
		158927 => x"FF",
		158928 => x"FF",
		158929 => x"FF",
		158930 => x"FF",
		158931 => x"FF",
		158932 => x"FF",
		158933 => x"FF",
		158934 => x"FF",
		158935 => x"FF",
		158936 => x"FF",
		158937 => x"FF",
		158938 => x"FF",
		158939 => x"FF",
		158940 => x"FF",
		158941 => x"FF",
		158942 => x"FF",
		158943 => x"FF",
		158944 => x"FF",
		158945 => x"FF",
		158946 => x"FF",
		158947 => x"FF",
		158948 => x"FF",
		158949 => x"FF",
		158950 => x"FF",
		158951 => x"FF",
		158952 => x"FF",
		158953 => x"FF",
		158954 => x"FF",
		158955 => x"FF",
		158956 => x"FF",
		158957 => x"FF",
		158958 => x"FF",
		158959 => x"FF",
		158960 => x"FF",
		158961 => x"FF",
		158962 => x"FF",
		158963 => x"FF",
		158964 => x"FF",
		158965 => x"FF",
		158966 => x"FF",
		158967 => x"FF",
		158968 => x"FF",
		158969 => x"FF",
		158970 => x"FF",
		158971 => x"FF",
		158972 => x"FF",
		158973 => x"FF",
		158974 => x"FF",
		158975 => x"FF",
		158976 => x"FF",
		158977 => x"FF",
		158978 => x"FF",
		158979 => x"FF",
		158980 => x"FF",
		158981 => x"FF",
		158982 => x"FF",
		158983 => x"FF",
		158984 => x"FF",
		158985 => x"FF",
		158986 => x"FF",
		158987 => x"FF",
		158988 => x"FF",
		158989 => x"FF",
		158990 => x"FF",
		158991 => x"FF",
		158992 => x"FF",
		158993 => x"FF",
		159788 => x"FF",
		159789 => x"FF",
		159790 => x"FF",
		159791 => x"FF",
		159792 => x"FF",
		159793 => x"FF",
		159794 => x"FF",
		159795 => x"FF",
		159796 => x"FF",
		159797 => x"FF",
		159798 => x"FF",
		159799 => x"FF",
		159800 => x"FF",
		159801 => x"FF",
		159802 => x"FF",
		159803 => x"FF",
		159804 => x"FF",
		159805 => x"FF",
		159806 => x"FF",
		159807 => x"FF",
		159808 => x"FF",
		159809 => x"FF",
		159810 => x"FF",
		159811 => x"FF",
		159812 => x"FF",
		159813 => x"FF",
		159814 => x"FF",
		159815 => x"FF",
		159816 => x"FF",
		159817 => x"FF",
		159818 => x"FF",
		159819 => x"FF",
		159820 => x"FF",
		159821 => x"FF",
		159822 => x"FF",
		159823 => x"FF",
		159824 => x"FF",
		159825 => x"FF",
		159826 => x"FF",
		159827 => x"FF",
		159828 => x"FF",
		159829 => x"FF",
		159830 => x"FF",
		159831 => x"FF",
		159832 => x"FF",
		159833 => x"FF",
		159834 => x"FF",
		159835 => x"FF",
		159836 => x"FF",
		159837 => x"FF",
		159838 => x"FF",
		159839 => x"FF",
		159840 => x"FF",
		159841 => x"FF",
		159842 => x"FF",
		159843 => x"FF",
		159844 => x"FF",
		159845 => x"FF",
		159846 => x"FF",
		159847 => x"FF",
		159848 => x"FF",
		159849 => x"FF",
		159850 => x"FF",
		159851 => x"FF",
		159852 => x"FF",
		159853 => x"FF",
		159854 => x"FF",
		159855 => x"FF",
		159856 => x"FF",
		159857 => x"FF",
		159858 => x"FF",
		159859 => x"FF",
		159860 => x"FF",
		159861 => x"FF",
		159862 => x"FF",
		159863 => x"FF",
		159864 => x"FF",
		159865 => x"FF",
		159866 => x"FF",
		159867 => x"FF",
		159868 => x"FF",
		159869 => x"FF",
		159870 => x"FF",
		159871 => x"FF",
		159872 => x"FF",
		159873 => x"FF",
		159874 => x"FF",
		159875 => x"FF",
		159876 => x"FF",
		159877 => x"FF",
		159878 => x"FF",
		159879 => x"FF",
		159880 => x"FF",
		159881 => x"FF",
		159882 => x"FF",
		159883 => x"FF",
		159884 => x"FF",
		159885 => x"FF",
		159886 => x"FF",
		159887 => x"FF",
		159888 => x"FF",
		159889 => x"FF",
		159890 => x"FF",
		159891 => x"FF",
		159892 => x"FF",
		159893 => x"FF",
		159894 => x"FF",
		159895 => x"FF",
		159896 => x"FF",
		159897 => x"FF",
		159898 => x"FF",
		159899 => x"FF",
		159900 => x"FF",
		159901 => x"FF",
		159902 => x"FF",
		159903 => x"FF",
		159904 => x"FF",
		159905 => x"FF",
		159906 => x"FF",
		159907 => x"FF",
		159908 => x"FF",
		159909 => x"FF",
		159910 => x"FF",
		159911 => x"FF",
		159912 => x"FF",
		159913 => x"FF",
		159914 => x"FF",
		159915 => x"FF",
		159916 => x"FF",
		159917 => x"FF",
		159918 => x"FF",
		159919 => x"FF",
		159920 => x"FF",
		159921 => x"FF",
		159922 => x"FF",
		159923 => x"FF",
		159924 => x"FF",
		159925 => x"FF",
		159926 => x"FF",
		159927 => x"FF",
		159928 => x"FF",
		159929 => x"FF",
		159930 => x"FF",
		159931 => x"FF",
		159932 => x"FF",
		159933 => x"FF",
		159934 => x"FF",
		159935 => x"FF",
		159936 => x"FF",
		159937 => x"FF",
		159938 => x"FF",
		159939 => x"FF",
		159940 => x"FF",
		159941 => x"FF",
		159942 => x"FF",
		159943 => x"FF",
		159944 => x"FF",
		159945 => x"FF",
		159946 => x"FF",
		159947 => x"FF",
		159948 => x"FF",
		159949 => x"FF",
		159950 => x"FF",
		159951 => x"FF",
		159952 => x"FF",
		159953 => x"FF",
		159954 => x"FF",
		159955 => x"FF",
		159956 => x"FF",
		159957 => x"FF",
		159958 => x"FF",
		159959 => x"FF",
		159960 => x"FF",
		159961 => x"FF",
		159962 => x"FF",
		159963 => x"FF",
		159964 => x"FF",
		159965 => x"FF",
		159966 => x"FF",
		159967 => x"FF",
		159968 => x"FF",
		159969 => x"FF",
		159970 => x"FF",
		159971 => x"FF",
		159972 => x"FF",
		159973 => x"FF",
		159974 => x"FF",
		159975 => x"FF",
		159976 => x"FF",
		159977 => x"FF",
		159978 => x"FF",
		159979 => x"FF",
		159980 => x"FF",
		159981 => x"FF",
		159982 => x"FF",
		159983 => x"FF",
		159984 => x"FF",
		159985 => x"FF",
		159986 => x"FF",
		159987 => x"FF",
		159988 => x"FF",
		159989 => x"FF",
		159990 => x"FF",
		159991 => x"FF",
		159992 => x"FF",
		159993 => x"FF",
		159994 => x"FF",
		159995 => x"FF",
		159996 => x"FF",
		159997 => x"FF",
		159998 => x"FF",
		159999 => x"FF",
		160000 => x"FF",
		160001 => x"FF",
		160002 => x"FF",
		160003 => x"FF",
		160004 => x"FF",
		160005 => x"FF",
		160006 => x"FF",
		160007 => x"FF",
		160008 => x"FF",
		160009 => x"FF",
		160010 => x"FF",
		160011 => x"FF",
		160012 => x"FF",
		160013 => x"FF",
		160014 => x"FF",
		160015 => x"FF",
		160016 => x"FF",
		160017 => x"FF",
		160812 => x"FF",
		160813 => x"FF",
		160814 => x"FF",
		160815 => x"FF",
		160816 => x"FF",
		160817 => x"FF",
		160818 => x"FF",
		160819 => x"FF",
		160820 => x"FF",
		160821 => x"FF",
		160822 => x"FF",
		160823 => x"FF",
		160824 => x"FF",
		160825 => x"FF",
		160826 => x"FF",
		160827 => x"FF",
		160828 => x"FF",
		160829 => x"FF",
		160830 => x"FF",
		160831 => x"FF",
		160832 => x"FF",
		160833 => x"FF",
		160834 => x"FF",
		160835 => x"FF",
		160836 => x"FF",
		160837 => x"FF",
		160838 => x"FF",
		160839 => x"FF",
		160840 => x"FF",
		160841 => x"FF",
		160842 => x"FF",
		160843 => x"FF",
		160844 => x"FF",
		160845 => x"FF",
		160846 => x"FF",
		160847 => x"FF",
		160848 => x"FF",
		160849 => x"FF",
		160850 => x"FF",
		160851 => x"FF",
		160852 => x"FF",
		160853 => x"FF",
		160854 => x"FF",
		160855 => x"FF",
		160856 => x"FF",
		160857 => x"FF",
		160858 => x"FF",
		160859 => x"FF",
		160860 => x"FF",
		160861 => x"FF",
		160862 => x"FF",
		160863 => x"FF",
		160864 => x"FF",
		160865 => x"FF",
		160866 => x"FF",
		160867 => x"FF",
		160868 => x"FF",
		160869 => x"FF",
		160870 => x"FF",
		160871 => x"FF",
		160872 => x"FF",
		160873 => x"FF",
		160874 => x"FF",
		160875 => x"FF",
		160876 => x"FF",
		160877 => x"FF",
		160878 => x"FF",
		160879 => x"FF",
		160880 => x"FF",
		160881 => x"FF",
		160882 => x"FF",
		160883 => x"FF",
		160884 => x"FF",
		160885 => x"FF",
		160886 => x"FF",
		160887 => x"FF",
		160888 => x"FF",
		160889 => x"FF",
		160890 => x"FF",
		160891 => x"FF",
		160892 => x"FF",
		160893 => x"FF",
		160894 => x"FF",
		160895 => x"FF",
		160896 => x"FF",
		160897 => x"FF",
		160898 => x"FF",
		160899 => x"FF",
		160900 => x"FF",
		160901 => x"FF",
		160902 => x"FF",
		160903 => x"FF",
		160904 => x"FF",
		160905 => x"FF",
		160906 => x"FF",
		160907 => x"FF",
		160908 => x"FF",
		160909 => x"FF",
		160910 => x"FF",
		160911 => x"FF",
		160912 => x"FF",
		160913 => x"FF",
		160914 => x"FF",
		160915 => x"FF",
		160916 => x"FF",
		160917 => x"FF",
		160918 => x"FF",
		160919 => x"FF",
		160920 => x"FF",
		160921 => x"FF",
		160922 => x"FF",
		160923 => x"FF",
		160924 => x"FF",
		160925 => x"FF",
		160926 => x"FF",
		160927 => x"FF",
		160928 => x"FF",
		160929 => x"FF",
		160930 => x"FF",
		160931 => x"FF",
		160932 => x"FF",
		160933 => x"FF",
		160934 => x"FF",
		160935 => x"FF",
		160936 => x"FF",
		160937 => x"FF",
		160938 => x"FF",
		160939 => x"FF",
		160940 => x"FF",
		160941 => x"FF",
		160942 => x"FF",
		160943 => x"FF",
		160944 => x"FF",
		160945 => x"FF",
		160946 => x"FF",
		160947 => x"FF",
		160948 => x"FF",
		160949 => x"FF",
		160950 => x"FF",
		160951 => x"FF",
		160952 => x"FF",
		160953 => x"FF",
		160954 => x"FF",
		160955 => x"FF",
		160956 => x"FF",
		160957 => x"FF",
		160958 => x"FF",
		160959 => x"FF",
		160960 => x"FF",
		160961 => x"FF",
		160962 => x"FF",
		160963 => x"FF",
		160964 => x"FF",
		160965 => x"FF",
		160966 => x"FF",
		160967 => x"FF",
		160968 => x"FF",
		160969 => x"FF",
		160970 => x"FF",
		160971 => x"FF",
		160972 => x"FF",
		160973 => x"FF",
		160974 => x"FF",
		160975 => x"FF",
		160976 => x"FF",
		160977 => x"FF",
		160978 => x"FF",
		160979 => x"FF",
		160980 => x"FF",
		160981 => x"FF",
		160982 => x"FF",
		160983 => x"FF",
		160984 => x"FF",
		160985 => x"FF",
		160986 => x"FF",
		160987 => x"FF",
		160988 => x"FF",
		160989 => x"FF",
		160990 => x"FF",
		160991 => x"FF",
		160992 => x"FF",
		160993 => x"FF",
		160994 => x"FF",
		160995 => x"FF",
		160996 => x"FF",
		160997 => x"FF",
		160998 => x"FF",
		160999 => x"FF",
		161000 => x"FF",
		161001 => x"FF",
		161002 => x"FF",
		161003 => x"FF",
		161004 => x"FF",
		161005 => x"FF",
		161006 => x"FF",
		161007 => x"FF",
		161008 => x"FF",
		161009 => x"FF",
		161010 => x"FF",
		161011 => x"FF",
		161012 => x"FF",
		161013 => x"FF",
		161014 => x"FF",
		161015 => x"FF",
		161016 => x"FF",
		161017 => x"FF",
		161018 => x"FF",
		161019 => x"FF",
		161020 => x"FF",
		161021 => x"FF",
		161022 => x"FF",
		161023 => x"FF",
		161024 => x"FF",
		161025 => x"FF",
		161026 => x"FF",
		161027 => x"FF",
		161028 => x"FF",
		161029 => x"FF",
		161030 => x"FF",
		161031 => x"FF",
		161032 => x"FF",
		161033 => x"FF",
		161034 => x"FF",
		161035 => x"FF",
		161036 => x"FF",
		161037 => x"FF",
		161038 => x"FF",
		161039 => x"FF",
		161040 => x"FF",
		161041 => x"FF",
		161836 => x"FF",
		161837 => x"FF",
		161838 => x"FF",
		161839 => x"FF",
		161840 => x"FF",
		161841 => x"FF",
		161842 => x"FF",
		161843 => x"FF",
		161844 => x"FF",
		161845 => x"FF",
		161846 => x"FF",
		161847 => x"FF",
		161848 => x"FF",
		161849 => x"FF",
		161850 => x"FF",
		161851 => x"FF",
		161852 => x"FF",
		161853 => x"FF",
		161854 => x"FF",
		161855 => x"FF",
		161856 => x"FF",
		161857 => x"FF",
		161858 => x"FF",
		161859 => x"FF",
		161860 => x"FF",
		161861 => x"FF",
		161862 => x"FF",
		161863 => x"FF",
		161864 => x"FF",
		161865 => x"FF",
		161866 => x"FF",
		161867 => x"FF",
		161868 => x"FF",
		161869 => x"FF",
		161870 => x"FF",
		161871 => x"FF",
		161872 => x"FF",
		161873 => x"FF",
		161874 => x"FF",
		161875 => x"FF",
		161876 => x"FF",
		161877 => x"FF",
		161878 => x"FF",
		161879 => x"FF",
		161880 => x"FF",
		161881 => x"FF",
		161882 => x"FF",
		161883 => x"FF",
		161884 => x"FF",
		161885 => x"FF",
		161886 => x"FF",
		161887 => x"FF",
		161888 => x"FF",
		161889 => x"FF",
		161890 => x"FF",
		161891 => x"FF",
		161892 => x"FF",
		161893 => x"FF",
		161894 => x"FF",
		161895 => x"FF",
		161896 => x"FF",
		161897 => x"FF",
		161898 => x"FF",
		161899 => x"FF",
		161900 => x"FF",
		161901 => x"FF",
		161902 => x"FF",
		161903 => x"FF",
		161904 => x"FF",
		161905 => x"FF",
		161906 => x"FF",
		161907 => x"FF",
		161908 => x"FF",
		161909 => x"FF",
		161910 => x"FF",
		161911 => x"FF",
		161912 => x"FF",
		161913 => x"FF",
		161914 => x"FF",
		161915 => x"FF",
		161916 => x"FF",
		161917 => x"FF",
		161918 => x"FF",
		161919 => x"FF",
		161920 => x"FF",
		161921 => x"FF",
		161922 => x"FF",
		161923 => x"FF",
		161924 => x"FF",
		161925 => x"FF",
		161926 => x"FF",
		161927 => x"FF",
		161928 => x"FF",
		161929 => x"FF",
		161930 => x"FF",
		161931 => x"FF",
		161932 => x"FF",
		161933 => x"FF",
		161934 => x"FF",
		161935 => x"FF",
		161936 => x"FF",
		161937 => x"FF",
		161938 => x"FF",
		161939 => x"FF",
		161940 => x"FF",
		161941 => x"FF",
		161942 => x"FF",
		161943 => x"FF",
		161944 => x"FF",
		161945 => x"FF",
		161946 => x"FF",
		161947 => x"FF",
		161948 => x"FF",
		161949 => x"FF",
		161950 => x"FF",
		161951 => x"FF",
		161952 => x"FF",
		161953 => x"FF",
		161954 => x"FF",
		161955 => x"FF",
		161956 => x"FF",
		161957 => x"FF",
		161958 => x"FF",
		161959 => x"FF",
		161960 => x"FF",
		161961 => x"FF",
		161962 => x"FF",
		161963 => x"FF",
		161964 => x"FF",
		161965 => x"FF",
		161966 => x"FF",
		161967 => x"FF",
		161968 => x"FF",
		161969 => x"FF",
		161970 => x"FF",
		161971 => x"FF",
		161972 => x"FF",
		161973 => x"FF",
		161974 => x"FF",
		161975 => x"FF",
		161976 => x"FF",
		161977 => x"FF",
		161978 => x"FF",
		161979 => x"FF",
		161980 => x"FF",
		161981 => x"FF",
		161982 => x"FF",
		161983 => x"FF",
		161984 => x"FF",
		161985 => x"FF",
		161986 => x"FF",
		161987 => x"FF",
		161988 => x"FF",
		161989 => x"FF",
		161990 => x"FF",
		161991 => x"FF",
		161992 => x"FF",
		161993 => x"FF",
		161994 => x"FF",
		161995 => x"FF",
		161996 => x"FF",
		161997 => x"FF",
		161998 => x"FF",
		161999 => x"FF",
		162000 => x"FF",
		162001 => x"FF",
		162002 => x"FF",
		162003 => x"FF",
		162004 => x"FF",
		162005 => x"FF",
		162006 => x"FF",
		162007 => x"FF",
		162008 => x"FF",
		162009 => x"FF",
		162010 => x"FF",
		162011 => x"FF",
		162012 => x"FF",
		162013 => x"FF",
		162014 => x"FF",
		162015 => x"FF",
		162016 => x"FF",
		162017 => x"FF",
		162018 => x"FF",
		162019 => x"FF",
		162020 => x"FF",
		162021 => x"FF",
		162022 => x"FF",
		162023 => x"FF",
		162024 => x"FF",
		162025 => x"FF",
		162026 => x"FF",
		162027 => x"FF",
		162028 => x"FF",
		162029 => x"FF",
		162030 => x"FF",
		162031 => x"FF",
		162032 => x"FF",
		162033 => x"FF",
		162034 => x"FF",
		162035 => x"FF",
		162036 => x"FF",
		162037 => x"FF",
		162038 => x"FF",
		162039 => x"FF",
		162040 => x"FF",
		162041 => x"FF",
		162042 => x"FF",
		162043 => x"FF",
		162044 => x"FF",
		162045 => x"FF",
		162046 => x"FF",
		162047 => x"FF",
		162048 => x"FF",
		162049 => x"FF",
		162050 => x"FF",
		162051 => x"FF",
		162052 => x"FF",
		162053 => x"FF",
		162054 => x"FF",
		162055 => x"FF",
		162056 => x"FF",
		162057 => x"FF",
		162058 => x"FF",
		162059 => x"FF",
		162060 => x"FF",
		162061 => x"FF",
		162062 => x"FF",
		162063 => x"FF",
		162064 => x"FF",
		162065 => x"FF",
		162860 => x"FF",
		162861 => x"FF",
		162862 => x"FF",
		162863 => x"FF",
		162864 => x"FF",
		162935 => x"FF",
		162936 => x"FF",
		162937 => x"FF",
		162938 => x"FF",
		162939 => x"FF",
		163010 => x"FF",
		163011 => x"FF",
		163012 => x"FF",
		163013 => x"FF",
		163014 => x"FF",
		163085 => x"FF",
		163086 => x"FF",
		163087 => x"FF",
		163088 => x"FF",
		163089 => x"FF",
		163884 => x"FF",
		163885 => x"FF",
		163886 => x"FF",
		163887 => x"FF",
		163888 => x"FF",
		163959 => x"FF",
		163960 => x"FF",
		163961 => x"FF",
		163962 => x"FF",
		163963 => x"FF",
		164034 => x"FF",
		164035 => x"FF",
		164036 => x"FF",
		164037 => x"FF",
		164038 => x"FF",
		164109 => x"FF",
		164110 => x"FF",
		164111 => x"FF",
		164112 => x"FF",
		164113 => x"FF",
		164908 => x"FF",
		164909 => x"FF",
		164910 => x"FF",
		164911 => x"FF",
		164912 => x"FF",
		164983 => x"FF",
		164984 => x"FF",
		164985 => x"FF",
		164986 => x"FF",
		164987 => x"FF",
		165058 => x"FF",
		165059 => x"FF",
		165060 => x"FF",
		165061 => x"FF",
		165062 => x"FF",
		165133 => x"FF",
		165134 => x"FF",
		165135 => x"FF",
		165136 => x"FF",
		165137 => x"FF",
		165932 => x"FF",
		165933 => x"FF",
		165934 => x"FF",
		165935 => x"FF",
		165936 => x"FF",
		166007 => x"FF",
		166008 => x"FF",
		166009 => x"FF",
		166010 => x"FF",
		166011 => x"FF",
		166082 => x"FF",
		166083 => x"FF",
		166084 => x"FF",
		166085 => x"FF",
		166086 => x"FF",
		166157 => x"FF",
		166158 => x"FF",
		166159 => x"FF",
		166160 => x"FF",
		166161 => x"FF",
		166956 => x"FF",
		166957 => x"FF",
		166958 => x"FF",
		166959 => x"FF",
		166960 => x"FF",
		167031 => x"FF",
		167032 => x"FF",
		167033 => x"FF",
		167034 => x"FF",
		167035 => x"FF",
		167106 => x"FF",
		167107 => x"FF",
		167108 => x"FF",
		167109 => x"FF",
		167110 => x"FF",
		167181 => x"FF",
		167182 => x"FF",
		167183 => x"FF",
		167184 => x"FF",
		167185 => x"FF",
		167980 => x"FF",
		167981 => x"FF",
		167982 => x"FF",
		167983 => x"FF",
		167984 => x"FF",
		168055 => x"FF",
		168056 => x"FF",
		168057 => x"FF",
		168058 => x"FF",
		168059 => x"FF",
		168130 => x"FF",
		168131 => x"FF",
		168132 => x"FF",
		168133 => x"FF",
		168134 => x"FF",
		168205 => x"FF",
		168206 => x"FF",
		168207 => x"FF",
		168208 => x"FF",
		168209 => x"FF",
		169004 => x"FF",
		169005 => x"FF",
		169006 => x"FF",
		169007 => x"FF",
		169008 => x"FF",
		169079 => x"FF",
		169080 => x"FF",
		169081 => x"FF",
		169082 => x"FF",
		169083 => x"FF",
		169154 => x"FF",
		169155 => x"FF",
		169156 => x"FF",
		169157 => x"FF",
		169158 => x"FF",
		169229 => x"FF",
		169230 => x"FF",
		169231 => x"FF",
		169232 => x"FF",
		169233 => x"FF",
		170028 => x"FF",
		170029 => x"FF",
		170030 => x"FF",
		170031 => x"FF",
		170032 => x"FF",
		170103 => x"FF",
		170104 => x"FF",
		170105 => x"FF",
		170106 => x"FF",
		170107 => x"FF",
		170178 => x"FF",
		170179 => x"FF",
		170180 => x"FF",
		170181 => x"FF",
		170182 => x"FF",
		170253 => x"FF",
		170254 => x"FF",
		170255 => x"FF",
		170256 => x"FF",
		170257 => x"FF",
		171052 => x"FF",
		171053 => x"FF",
		171054 => x"FF",
		171055 => x"FF",
		171056 => x"FF",
		171127 => x"FF",
		171128 => x"FF",
		171129 => x"FF",
		171130 => x"FF",
		171131 => x"FF",
		171202 => x"FF",
		171203 => x"FF",
		171204 => x"FF",
		171205 => x"FF",
		171206 => x"FF",
		171277 => x"FF",
		171278 => x"FF",
		171279 => x"FF",
		171280 => x"FF",
		171281 => x"FF",
		172076 => x"FF",
		172077 => x"FF",
		172078 => x"FF",
		172079 => x"FF",
		172080 => x"FF",
		172151 => x"FF",
		172152 => x"FF",
		172153 => x"FF",
		172154 => x"FF",
		172155 => x"FF",
		172226 => x"FF",
		172227 => x"FF",
		172228 => x"FF",
		172229 => x"FF",
		172230 => x"FF",
		172301 => x"FF",
		172302 => x"FF",
		172303 => x"FF",
		172304 => x"FF",
		172305 => x"FF",
		173100 => x"FF",
		173101 => x"FF",
		173102 => x"FF",
		173103 => x"FF",
		173104 => x"FF",
		173175 => x"FF",
		173176 => x"FF",
		173177 => x"FF",
		173178 => x"FF",
		173179 => x"FF",
		173250 => x"FF",
		173251 => x"FF",
		173252 => x"FF",
		173253 => x"FF",
		173254 => x"FF",
		173325 => x"FF",
		173326 => x"FF",
		173327 => x"FF",
		173328 => x"FF",
		173329 => x"FF",
		174124 => x"FF",
		174125 => x"FF",
		174126 => x"FF",
		174127 => x"FF",
		174128 => x"FF",
		174199 => x"FF",
		174200 => x"FF",
		174201 => x"FF",
		174202 => x"FF",
		174203 => x"FF",
		174274 => x"FF",
		174275 => x"FF",
		174276 => x"FF",
		174277 => x"FF",
		174278 => x"FF",
		174349 => x"FF",
		174350 => x"FF",
		174351 => x"FF",
		174352 => x"FF",
		174353 => x"FF",
		175148 => x"FF",
		175149 => x"FF",
		175150 => x"FF",
		175151 => x"FF",
		175152 => x"FF",
		175223 => x"FF",
		175224 => x"FF",
		175225 => x"FF",
		175226 => x"FF",
		175227 => x"FF",
		175298 => x"FF",
		175299 => x"FF",
		175300 => x"FF",
		175301 => x"FF",
		175302 => x"FF",
		175373 => x"FF",
		175374 => x"FF",
		175375 => x"FF",
		175376 => x"FF",
		175377 => x"FF",
		176172 => x"FF",
		176173 => x"FF",
		176174 => x"FF",
		176175 => x"FF",
		176176 => x"FF",
		176247 => x"FF",
		176248 => x"FF",
		176249 => x"FF",
		176250 => x"FF",
		176251 => x"FF",
		176322 => x"FF",
		176323 => x"FF",
		176324 => x"FF",
		176325 => x"FF",
		176326 => x"FF",
		176397 => x"FF",
		176398 => x"FF",
		176399 => x"FF",
		176400 => x"FF",
		176401 => x"FF",
		177196 => x"FF",
		177197 => x"FF",
		177198 => x"FF",
		177199 => x"FF",
		177200 => x"FF",
		177271 => x"FF",
		177272 => x"FF",
		177273 => x"FF",
		177274 => x"FF",
		177275 => x"FF",
		177346 => x"FF",
		177347 => x"FF",
		177348 => x"FF",
		177349 => x"FF",
		177350 => x"FF",
		177421 => x"FF",
		177422 => x"FF",
		177423 => x"FF",
		177424 => x"FF",
		177425 => x"FF",
		178220 => x"FF",
		178221 => x"FF",
		178222 => x"FF",
		178223 => x"FF",
		178224 => x"FF",
		178295 => x"FF",
		178296 => x"FF",
		178297 => x"FF",
		178298 => x"FF",
		178299 => x"FF",
		178370 => x"FF",
		178371 => x"FF",
		178372 => x"FF",
		178373 => x"FF",
		178374 => x"FF",
		178445 => x"FF",
		178446 => x"FF",
		178447 => x"FF",
		178448 => x"FF",
		178449 => x"FF",
		179244 => x"FF",
		179245 => x"FF",
		179246 => x"FF",
		179247 => x"FF",
		179248 => x"FF",
		179319 => x"FF",
		179320 => x"FF",
		179321 => x"FF",
		179322 => x"FF",
		179323 => x"FF",
		179394 => x"FF",
		179395 => x"FF",
		179396 => x"FF",
		179397 => x"FF",
		179398 => x"FF",
		179469 => x"FF",
		179470 => x"FF",
		179471 => x"FF",
		179472 => x"FF",
		179473 => x"FF",
		180268 => x"FF",
		180269 => x"FF",
		180270 => x"FF",
		180271 => x"FF",
		180272 => x"FF",
		180343 => x"FF",
		180344 => x"FF",
		180345 => x"FF",
		180346 => x"FF",
		180347 => x"FF",
		180418 => x"FF",
		180419 => x"FF",
		180420 => x"FF",
		180421 => x"FF",
		180422 => x"FF",
		180493 => x"FF",
		180494 => x"FF",
		180495 => x"FF",
		180496 => x"FF",
		180497 => x"FF",
		181292 => x"FF",
		181293 => x"FF",
		181294 => x"FF",
		181295 => x"FF",
		181296 => x"FF",
		181367 => x"FF",
		181368 => x"FF",
		181369 => x"FF",
		181370 => x"FF",
		181371 => x"FF",
		181442 => x"FF",
		181443 => x"FF",
		181444 => x"FF",
		181445 => x"FF",
		181446 => x"FF",
		181517 => x"FF",
		181518 => x"FF",
		181519 => x"FF",
		181520 => x"FF",
		181521 => x"FF",
		182316 => x"FF",
		182317 => x"FF",
		182318 => x"FF",
		182319 => x"FF",
		182320 => x"FF",
		182391 => x"FF",
		182392 => x"FF",
		182393 => x"FF",
		182394 => x"FF",
		182395 => x"FF",
		182466 => x"FF",
		182467 => x"FF",
		182468 => x"FF",
		182469 => x"FF",
		182470 => x"FF",
		182541 => x"FF",
		182542 => x"FF",
		182543 => x"FF",
		182544 => x"FF",
		182545 => x"FF",
		183340 => x"FF",
		183341 => x"FF",
		183342 => x"FF",
		183343 => x"FF",
		183344 => x"FF",
		183415 => x"FF",
		183416 => x"FF",
		183417 => x"FF",
		183418 => x"FF",
		183419 => x"FF",
		183490 => x"FF",
		183491 => x"FF",
		183492 => x"FF",
		183493 => x"FF",
		183494 => x"FF",
		183565 => x"FF",
		183566 => x"FF",
		183567 => x"FF",
		183568 => x"FF",
		183569 => x"FF",
		184364 => x"FF",
		184365 => x"FF",
		184366 => x"FF",
		184367 => x"FF",
		184368 => x"FF",
		184439 => x"FF",
		184440 => x"FF",
		184441 => x"FF",
		184442 => x"FF",
		184443 => x"FF",
		184514 => x"FF",
		184515 => x"FF",
		184516 => x"FF",
		184517 => x"FF",
		184518 => x"FF",
		184589 => x"FF",
		184590 => x"FF",
		184591 => x"FF",
		184592 => x"FF",
		184593 => x"FF",
		185388 => x"FF",
		185389 => x"FF",
		185390 => x"FF",
		185391 => x"FF",
		185392 => x"FF",
		185463 => x"FF",
		185464 => x"FF",
		185465 => x"FF",
		185466 => x"FF",
		185467 => x"FF",
		185538 => x"FF",
		185539 => x"FF",
		185540 => x"FF",
		185541 => x"FF",
		185542 => x"FF",
		185613 => x"FF",
		185614 => x"FF",
		185615 => x"FF",
		185616 => x"FF",
		185617 => x"FF",
		186412 => x"FF",
		186413 => x"FF",
		186414 => x"FF",
		186415 => x"FF",
		186416 => x"FF",
		186487 => x"FF",
		186488 => x"FF",
		186489 => x"FF",
		186490 => x"FF",
		186491 => x"FF",
		186562 => x"FF",
		186563 => x"FF",
		186564 => x"FF",
		186565 => x"FF",
		186566 => x"FF",
		186637 => x"FF",
		186638 => x"FF",
		186639 => x"FF",
		186640 => x"FF",
		186641 => x"FF",
		187436 => x"FF",
		187437 => x"FF",
		187438 => x"FF",
		187439 => x"FF",
		187440 => x"FF",
		187511 => x"FF",
		187512 => x"FF",
		187513 => x"FF",
		187514 => x"FF",
		187515 => x"FF",
		187586 => x"FF",
		187587 => x"FF",
		187588 => x"FF",
		187589 => x"FF",
		187590 => x"FF",
		187661 => x"FF",
		187662 => x"FF",
		187663 => x"FF",
		187664 => x"FF",
		187665 => x"FF",
		188460 => x"FF",
		188461 => x"FF",
		188462 => x"FF",
		188463 => x"FF",
		188464 => x"FF",
		188535 => x"FF",
		188536 => x"FF",
		188537 => x"FF",
		188538 => x"FF",
		188539 => x"FF",
		188610 => x"FF",
		188611 => x"FF",
		188612 => x"FF",
		188613 => x"FF",
		188614 => x"FF",
		188685 => x"FF",
		188686 => x"FF",
		188687 => x"FF",
		188688 => x"FF",
		188689 => x"FF",
		189484 => x"FF",
		189485 => x"FF",
		189486 => x"FF",
		189487 => x"FF",
		189488 => x"FF",
		189559 => x"FF",
		189560 => x"FF",
		189561 => x"FF",
		189562 => x"FF",
		189563 => x"FF",
		189634 => x"FF",
		189635 => x"FF",
		189636 => x"FF",
		189637 => x"FF",
		189638 => x"FF",
		189709 => x"FF",
		189710 => x"FF",
		189711 => x"FF",
		189712 => x"FF",
		189713 => x"FF",
		190508 => x"FF",
		190509 => x"FF",
		190510 => x"FF",
		190511 => x"FF",
		190512 => x"FF",
		190583 => x"FF",
		190584 => x"FF",
		190585 => x"FF",
		190586 => x"FF",
		190587 => x"FF",
		190658 => x"FF",
		190659 => x"FF",
		190660 => x"FF",
		190661 => x"FF",
		190662 => x"FF",
		190733 => x"FF",
		190734 => x"FF",
		190735 => x"FF",
		190736 => x"FF",
		190737 => x"FF",
		191532 => x"FF",
		191533 => x"FF",
		191534 => x"FF",
		191535 => x"FF",
		191536 => x"FF",
		191607 => x"FF",
		191608 => x"FF",
		191609 => x"FF",
		191610 => x"FF",
		191611 => x"FF",
		191682 => x"FF",
		191683 => x"FF",
		191684 => x"FF",
		191685 => x"FF",
		191686 => x"FF",
		191757 => x"FF",
		191758 => x"FF",
		191759 => x"FF",
		191760 => x"FF",
		191761 => x"FF",
		192556 => x"FF",
		192557 => x"FF",
		192558 => x"FF",
		192559 => x"FF",
		192560 => x"FF",
		192631 => x"FF",
		192632 => x"FF",
		192633 => x"FF",
		192634 => x"FF",
		192635 => x"FF",
		192706 => x"FF",
		192707 => x"FF",
		192708 => x"FF",
		192709 => x"FF",
		192710 => x"FF",
		192781 => x"FF",
		192782 => x"FF",
		192783 => x"FF",
		192784 => x"FF",
		192785 => x"FF",
		193580 => x"FF",
		193581 => x"FF",
		193582 => x"FF",
		193583 => x"FF",
		193584 => x"FF",
		193655 => x"FF",
		193656 => x"FF",
		193657 => x"FF",
		193658 => x"FF",
		193659 => x"FF",
		193730 => x"FF",
		193731 => x"FF",
		193732 => x"FF",
		193733 => x"FF",
		193734 => x"FF",
		193805 => x"FF",
		193806 => x"FF",
		193807 => x"FF",
		193808 => x"FF",
		193809 => x"FF",
		194604 => x"FF",
		194605 => x"FF",
		194606 => x"FF",
		194607 => x"FF",
		194608 => x"FF",
		194679 => x"FF",
		194680 => x"FF",
		194681 => x"FF",
		194682 => x"FF",
		194683 => x"FF",
		194754 => x"FF",
		194755 => x"FF",
		194756 => x"FF",
		194757 => x"FF",
		194758 => x"FF",
		194829 => x"FF",
		194830 => x"FF",
		194831 => x"FF",
		194832 => x"FF",
		194833 => x"FF",
		195628 => x"FF",
		195629 => x"FF",
		195630 => x"FF",
		195631 => x"FF",
		195632 => x"FF",
		195703 => x"FF",
		195704 => x"FF",
		195705 => x"FF",
		195706 => x"FF",
		195707 => x"FF",
		195778 => x"FF",
		195779 => x"FF",
		195780 => x"FF",
		195781 => x"FF",
		195782 => x"FF",
		195853 => x"FF",
		195854 => x"FF",
		195855 => x"FF",
		195856 => x"FF",
		195857 => x"FF",
		196652 => x"FF",
		196653 => x"FF",
		196654 => x"FF",
		196655 => x"FF",
		196656 => x"FF",
		196727 => x"FF",
		196728 => x"FF",
		196729 => x"FF",
		196730 => x"FF",
		196731 => x"FF",
		196802 => x"FF",
		196803 => x"FF",
		196804 => x"FF",
		196805 => x"FF",
		196806 => x"FF",
		196877 => x"FF",
		196878 => x"FF",
		196879 => x"FF",
		196880 => x"FF",
		196881 => x"FF",
		197676 => x"FF",
		197677 => x"FF",
		197678 => x"FF",
		197679 => x"FF",
		197680 => x"FF",
		197751 => x"FF",
		197752 => x"FF",
		197753 => x"FF",
		197754 => x"FF",
		197755 => x"FF",
		197826 => x"FF",
		197827 => x"FF",
		197828 => x"FF",
		197829 => x"FF",
		197830 => x"FF",
		197901 => x"FF",
		197902 => x"FF",
		197903 => x"FF",
		197904 => x"FF",
		197905 => x"FF",
		198700 => x"FF",
		198701 => x"FF",
		198702 => x"FF",
		198703 => x"FF",
		198704 => x"FF",
		198775 => x"FF",
		198776 => x"FF",
		198777 => x"FF",
		198778 => x"FF",
		198779 => x"FF",
		198850 => x"FF",
		198851 => x"FF",
		198852 => x"FF",
		198853 => x"FF",
		198854 => x"FF",
		198925 => x"FF",
		198926 => x"FF",
		198927 => x"FF",
		198928 => x"FF",
		198929 => x"FF",
		199724 => x"FF",
		199725 => x"FF",
		199726 => x"FF",
		199727 => x"FF",
		199728 => x"FF",
		199799 => x"FF",
		199800 => x"FF",
		199801 => x"FF",
		199802 => x"FF",
		199803 => x"FF",
		199874 => x"FF",
		199875 => x"FF",
		199876 => x"FF",
		199877 => x"FF",
		199878 => x"FF",
		199949 => x"FF",
		199950 => x"FF",
		199951 => x"FF",
		199952 => x"FF",
		199953 => x"FF",
		200748 => x"FF",
		200749 => x"FF",
		200750 => x"FF",
		200751 => x"FF",
		200752 => x"FF",
		200823 => x"FF",
		200824 => x"FF",
		200825 => x"FF",
		200826 => x"FF",
		200827 => x"FF",
		200898 => x"FF",
		200899 => x"FF",
		200900 => x"FF",
		200901 => x"FF",
		200902 => x"FF",
		200973 => x"FF",
		200974 => x"FF",
		200975 => x"FF",
		200976 => x"FF",
		200977 => x"FF",
		201772 => x"FF",
		201773 => x"FF",
		201774 => x"FF",
		201775 => x"FF",
		201776 => x"FF",
		201847 => x"FF",
		201848 => x"FF",
		201849 => x"FF",
		201850 => x"FF",
		201851 => x"FF",
		201922 => x"FF",
		201923 => x"FF",
		201924 => x"FF",
		201925 => x"FF",
		201926 => x"FF",
		201997 => x"FF",
		201998 => x"FF",
		201999 => x"FF",
		202000 => x"FF",
		202001 => x"FF",
		202796 => x"FF",
		202797 => x"FF",
		202798 => x"FF",
		202799 => x"FF",
		202800 => x"FF",
		202871 => x"FF",
		202872 => x"FF",
		202873 => x"FF",
		202874 => x"FF",
		202875 => x"FF",
		202946 => x"FF",
		202947 => x"FF",
		202948 => x"FF",
		202949 => x"FF",
		202950 => x"FF",
		203021 => x"FF",
		203022 => x"FF",
		203023 => x"FF",
		203024 => x"FF",
		203025 => x"FF",
		203820 => x"FF",
		203821 => x"FF",
		203822 => x"FF",
		203823 => x"FF",
		203824 => x"FF",
		203895 => x"FF",
		203896 => x"FF",
		203897 => x"FF",
		203898 => x"FF",
		203899 => x"FF",
		203970 => x"FF",
		203971 => x"FF",
		203972 => x"FF",
		203973 => x"FF",
		203974 => x"FF",
		204045 => x"FF",
		204046 => x"FF",
		204047 => x"FF",
		204048 => x"FF",
		204049 => x"FF",
		204844 => x"FF",
		204845 => x"FF",
		204846 => x"FF",
		204847 => x"FF",
		204848 => x"FF",
		204919 => x"FF",
		204920 => x"FF",
		204921 => x"FF",
		204922 => x"FF",
		204923 => x"FF",
		204994 => x"FF",
		204995 => x"FF",
		204996 => x"FF",
		204997 => x"FF",
		204998 => x"FF",
		205069 => x"FF",
		205070 => x"FF",
		205071 => x"FF",
		205072 => x"FF",
		205073 => x"FF",
		205868 => x"FF",
		205869 => x"FF",
		205870 => x"FF",
		205871 => x"FF",
		205872 => x"FF",
		205943 => x"FF",
		205944 => x"FF",
		205945 => x"FF",
		205946 => x"FF",
		205947 => x"FF",
		206018 => x"FF",
		206019 => x"FF",
		206020 => x"FF",
		206021 => x"FF",
		206022 => x"FF",
		206093 => x"FF",
		206094 => x"FF",
		206095 => x"FF",
		206096 => x"FF",
		206097 => x"FF",
		206892 => x"FF",
		206893 => x"FF",
		206894 => x"FF",
		206895 => x"FF",
		206896 => x"FF",
		206967 => x"FF",
		206968 => x"FF",
		206969 => x"FF",
		206970 => x"FF",
		206971 => x"FF",
		207042 => x"FF",
		207043 => x"FF",
		207044 => x"FF",
		207045 => x"FF",
		207046 => x"FF",
		207117 => x"FF",
		207118 => x"FF",
		207119 => x"FF",
		207120 => x"FF",
		207121 => x"FF",
		207916 => x"FF",
		207917 => x"FF",
		207918 => x"FF",
		207919 => x"FF",
		207920 => x"FF",
		207991 => x"FF",
		207992 => x"FF",
		207993 => x"FF",
		207994 => x"FF",
		207995 => x"FF",
		208066 => x"FF",
		208067 => x"FF",
		208068 => x"FF",
		208069 => x"FF",
		208070 => x"FF",
		208141 => x"FF",
		208142 => x"FF",
		208143 => x"FF",
		208144 => x"FF",
		208145 => x"FF",
		208940 => x"FF",
		208941 => x"FF",
		208942 => x"FF",
		208943 => x"FF",
		208944 => x"FF",
		209015 => x"FF",
		209016 => x"FF",
		209017 => x"FF",
		209018 => x"FF",
		209019 => x"FF",
		209090 => x"FF",
		209091 => x"FF",
		209092 => x"FF",
		209093 => x"FF",
		209094 => x"FF",
		209165 => x"FF",
		209166 => x"FF",
		209167 => x"FF",
		209168 => x"FF",
		209169 => x"FF",
		209964 => x"FF",
		209965 => x"FF",
		209966 => x"FF",
		209967 => x"FF",
		209968 => x"FF",
		210039 => x"FF",
		210040 => x"FF",
		210041 => x"FF",
		210042 => x"FF",
		210043 => x"FF",
		210114 => x"FF",
		210115 => x"FF",
		210116 => x"FF",
		210117 => x"FF",
		210118 => x"FF",
		210189 => x"FF",
		210190 => x"FF",
		210191 => x"FF",
		210192 => x"FF",
		210193 => x"FF",
		210988 => x"FF",
		210989 => x"FF",
		210990 => x"FF",
		210991 => x"FF",
		210992 => x"FF",
		211063 => x"FF",
		211064 => x"FF",
		211065 => x"FF",
		211066 => x"FF",
		211067 => x"FF",
		211138 => x"FF",
		211139 => x"FF",
		211140 => x"FF",
		211141 => x"FF",
		211142 => x"FF",
		211213 => x"FF",
		211214 => x"FF",
		211215 => x"FF",
		211216 => x"FF",
		211217 => x"FF",
		212012 => x"FF",
		212013 => x"FF",
		212014 => x"FF",
		212015 => x"FF",
		212016 => x"FF",
		212087 => x"FF",
		212088 => x"FF",
		212089 => x"FF",
		212090 => x"FF",
		212091 => x"FF",
		212162 => x"FF",
		212163 => x"FF",
		212164 => x"FF",
		212165 => x"FF",
		212166 => x"FF",
		212237 => x"FF",
		212238 => x"FF",
		212239 => x"FF",
		212240 => x"FF",
		212241 => x"FF",
		213036 => x"FF",
		213037 => x"FF",
		213038 => x"FF",
		213039 => x"FF",
		213040 => x"FF",
		213111 => x"FF",
		213112 => x"FF",
		213113 => x"FF",
		213114 => x"FF",
		213115 => x"FF",
		213186 => x"FF",
		213187 => x"FF",
		213188 => x"FF",
		213189 => x"FF",
		213190 => x"FF",
		213261 => x"FF",
		213262 => x"FF",
		213263 => x"FF",
		213264 => x"FF",
		213265 => x"FF",
		214060 => x"FF",
		214061 => x"FF",
		214062 => x"FF",
		214063 => x"FF",
		214064 => x"FF",
		214135 => x"FF",
		214136 => x"FF",
		214137 => x"FF",
		214138 => x"FF",
		214139 => x"FF",
		214210 => x"FF",
		214211 => x"FF",
		214212 => x"FF",
		214213 => x"FF",
		214214 => x"FF",
		214285 => x"FF",
		214286 => x"FF",
		214287 => x"FF",
		214288 => x"FF",
		214289 => x"FF",
		215084 => x"FF",
		215085 => x"FF",
		215086 => x"FF",
		215087 => x"FF",
		215088 => x"FF",
		215159 => x"FF",
		215160 => x"FF",
		215161 => x"FF",
		215162 => x"FF",
		215163 => x"FF",
		215234 => x"FF",
		215235 => x"FF",
		215236 => x"FF",
		215237 => x"FF",
		215238 => x"FF",
		215309 => x"FF",
		215310 => x"FF",
		215311 => x"FF",
		215312 => x"FF",
		215313 => x"FF",
		216108 => x"FF",
		216109 => x"FF",
		216110 => x"FF",
		216111 => x"FF",
		216112 => x"FF",
		216183 => x"FF",
		216184 => x"FF",
		216185 => x"FF",
		216186 => x"FF",
		216187 => x"FF",
		216258 => x"FF",
		216259 => x"FF",
		216260 => x"FF",
		216261 => x"FF",
		216262 => x"FF",
		216333 => x"FF",
		216334 => x"FF",
		216335 => x"FF",
		216336 => x"FF",
		216337 => x"FF",
		217132 => x"FF",
		217133 => x"FF",
		217134 => x"FF",
		217135 => x"FF",
		217136 => x"FF",
		217207 => x"FF",
		217208 => x"FF",
		217209 => x"FF",
		217210 => x"FF",
		217211 => x"FF",
		217282 => x"FF",
		217283 => x"FF",
		217284 => x"FF",
		217285 => x"FF",
		217286 => x"FF",
		217357 => x"FF",
		217358 => x"FF",
		217359 => x"FF",
		217360 => x"FF",
		217361 => x"FF",
		218156 => x"FF",
		218157 => x"FF",
		218158 => x"FF",
		218159 => x"FF",
		218160 => x"FF",
		218231 => x"FF",
		218232 => x"FF",
		218233 => x"FF",
		218234 => x"FF",
		218235 => x"FF",
		218306 => x"FF",
		218307 => x"FF",
		218308 => x"FF",
		218309 => x"FF",
		218310 => x"FF",
		218381 => x"FF",
		218382 => x"FF",
		218383 => x"FF",
		218384 => x"FF",
		218385 => x"FF",
		219180 => x"FF",
		219181 => x"FF",
		219182 => x"FF",
		219183 => x"FF",
		219184 => x"FF",
		219255 => x"FF",
		219256 => x"FF",
		219257 => x"FF",
		219258 => x"FF",
		219259 => x"FF",
		219330 => x"FF",
		219331 => x"FF",
		219332 => x"FF",
		219333 => x"FF",
		219334 => x"FF",
		219405 => x"FF",
		219406 => x"FF",
		219407 => x"FF",
		219408 => x"FF",
		219409 => x"FF",
		220204 => x"FF",
		220205 => x"FF",
		220206 => x"FF",
		220207 => x"FF",
		220208 => x"FF",
		220279 => x"FF",
		220280 => x"FF",
		220281 => x"FF",
		220282 => x"FF",
		220283 => x"FF",
		220354 => x"FF",
		220355 => x"FF",
		220356 => x"FF",
		220357 => x"FF",
		220358 => x"FF",
		220429 => x"FF",
		220430 => x"FF",
		220431 => x"FF",
		220432 => x"FF",
		220433 => x"FF",
		221228 => x"FF",
		221229 => x"FF",
		221230 => x"FF",
		221231 => x"FF",
		221232 => x"FF",
		221303 => x"FF",
		221304 => x"FF",
		221305 => x"FF",
		221306 => x"FF",
		221307 => x"FF",
		221378 => x"FF",
		221379 => x"FF",
		221380 => x"FF",
		221381 => x"FF",
		221382 => x"FF",
		221453 => x"FF",
		221454 => x"FF",
		221455 => x"FF",
		221456 => x"FF",
		221457 => x"FF",
		222252 => x"FF",
		222253 => x"FF",
		222254 => x"FF",
		222255 => x"FF",
		222256 => x"FF",
		222327 => x"FF",
		222328 => x"FF",
		222329 => x"FF",
		222330 => x"FF",
		222331 => x"FF",
		222402 => x"FF",
		222403 => x"FF",
		222404 => x"FF",
		222405 => x"FF",
		222406 => x"FF",
		222477 => x"FF",
		222478 => x"FF",
		222479 => x"FF",
		222480 => x"FF",
		222481 => x"FF",
		223276 => x"FF",
		223277 => x"FF",
		223278 => x"FF",
		223279 => x"FF",
		223280 => x"FF",
		223351 => x"FF",
		223352 => x"FF",
		223353 => x"FF",
		223354 => x"FF",
		223355 => x"FF",
		223426 => x"FF",
		223427 => x"FF",
		223428 => x"FF",
		223429 => x"FF",
		223430 => x"FF",
		223501 => x"FF",
		223502 => x"FF",
		223503 => x"FF",
		223504 => x"FF",
		223505 => x"FF",
		224300 => x"FF",
		224301 => x"FF",
		224302 => x"FF",
		224303 => x"FF",
		224304 => x"FF",
		224375 => x"FF",
		224376 => x"FF",
		224377 => x"FF",
		224378 => x"FF",
		224379 => x"FF",
		224450 => x"FF",
		224451 => x"FF",
		224452 => x"FF",
		224453 => x"FF",
		224454 => x"FF",
		224525 => x"FF",
		224526 => x"FF",
		224527 => x"FF",
		224528 => x"FF",
		224529 => x"FF",
		225324 => x"FF",
		225325 => x"FF",
		225326 => x"FF",
		225327 => x"FF",
		225328 => x"FF",
		225399 => x"FF",
		225400 => x"FF",
		225401 => x"FF",
		225402 => x"FF",
		225403 => x"FF",
		225474 => x"FF",
		225475 => x"FF",
		225476 => x"FF",
		225477 => x"FF",
		225478 => x"FF",
		225549 => x"FF",
		225550 => x"FF",
		225551 => x"FF",
		225552 => x"FF",
		225553 => x"FF",
		226348 => x"FF",
		226349 => x"FF",
		226350 => x"FF",
		226351 => x"FF",
		226352 => x"FF",
		226423 => x"FF",
		226424 => x"FF",
		226425 => x"FF",
		226426 => x"FF",
		226427 => x"FF",
		226498 => x"FF",
		226499 => x"FF",
		226500 => x"FF",
		226501 => x"FF",
		226502 => x"FF",
		226573 => x"FF",
		226574 => x"FF",
		226575 => x"FF",
		226576 => x"FF",
		226577 => x"FF",
		227372 => x"FF",
		227373 => x"FF",
		227374 => x"FF",
		227375 => x"FF",
		227376 => x"FF",
		227447 => x"FF",
		227448 => x"FF",
		227449 => x"FF",
		227450 => x"FF",
		227451 => x"FF",
		227522 => x"FF",
		227523 => x"FF",
		227524 => x"FF",
		227525 => x"FF",
		227526 => x"FF",
		227597 => x"FF",
		227598 => x"FF",
		227599 => x"FF",
		227600 => x"FF",
		227601 => x"FF",
		228396 => x"FF",
		228397 => x"FF",
		228398 => x"FF",
		228399 => x"FF",
		228400 => x"FF",
		228471 => x"FF",
		228472 => x"FF",
		228473 => x"FF",
		228474 => x"FF",
		228475 => x"FF",
		228546 => x"FF",
		228547 => x"FF",
		228548 => x"FF",
		228549 => x"FF",
		228550 => x"FF",
		228621 => x"FF",
		228622 => x"FF",
		228623 => x"FF",
		228624 => x"FF",
		228625 => x"FF",
		229420 => x"FF",
		229421 => x"FF",
		229422 => x"FF",
		229423 => x"FF",
		229424 => x"FF",
		229495 => x"FF",
		229496 => x"FF",
		229497 => x"FF",
		229498 => x"FF",
		229499 => x"FF",
		229570 => x"FF",
		229571 => x"FF",
		229572 => x"FF",
		229573 => x"FF",
		229574 => x"FF",
		229645 => x"FF",
		229646 => x"FF",
		229647 => x"FF",
		229648 => x"FF",
		229649 => x"FF",
		230444 => x"FF",
		230445 => x"FF",
		230446 => x"FF",
		230447 => x"FF",
		230448 => x"FF",
		230519 => x"FF",
		230520 => x"FF",
		230521 => x"FF",
		230522 => x"FF",
		230523 => x"FF",
		230594 => x"FF",
		230595 => x"FF",
		230596 => x"FF",
		230597 => x"FF",
		230598 => x"FF",
		230669 => x"FF",
		230670 => x"FF",
		230671 => x"FF",
		230672 => x"FF",
		230673 => x"FF",
		231468 => x"FF",
		231469 => x"FF",
		231470 => x"FF",
		231471 => x"FF",
		231472 => x"FF",
		231543 => x"FF",
		231544 => x"FF",
		231545 => x"FF",
		231546 => x"FF",
		231547 => x"FF",
		231618 => x"FF",
		231619 => x"FF",
		231620 => x"FF",
		231621 => x"FF",
		231622 => x"FF",
		231693 => x"FF",
		231694 => x"FF",
		231695 => x"FF",
		231696 => x"FF",
		231697 => x"FF",
		232492 => x"FF",
		232493 => x"FF",
		232494 => x"FF",
		232495 => x"FF",
		232496 => x"FF",
		232567 => x"FF",
		232568 => x"FF",
		232569 => x"FF",
		232570 => x"FF",
		232571 => x"FF",
		232642 => x"FF",
		232643 => x"FF",
		232644 => x"FF",
		232645 => x"FF",
		232646 => x"FF",
		232717 => x"FF",
		232718 => x"FF",
		232719 => x"FF",
		232720 => x"FF",
		232721 => x"FF",
		233516 => x"FF",
		233517 => x"FF",
		233518 => x"FF",
		233519 => x"FF",
		233520 => x"FF",
		233591 => x"FF",
		233592 => x"FF",
		233593 => x"FF",
		233594 => x"FF",
		233595 => x"FF",
		233666 => x"FF",
		233667 => x"FF",
		233668 => x"FF",
		233669 => x"FF",
		233670 => x"FF",
		233741 => x"FF",
		233742 => x"FF",
		233743 => x"FF",
		233744 => x"FF",
		233745 => x"FF",
		234540 => x"FF",
		234541 => x"FF",
		234542 => x"FF",
		234543 => x"FF",
		234544 => x"FF",
		234545 => x"FF",
		234546 => x"FF",
		234547 => x"FF",
		234548 => x"FF",
		234549 => x"FF",
		234550 => x"FF",
		234551 => x"FF",
		234552 => x"FF",
		234553 => x"FF",
		234554 => x"FF",
		234555 => x"FF",
		234556 => x"FF",
		234557 => x"FF",
		234558 => x"FF",
		234559 => x"FF",
		234560 => x"FF",
		234561 => x"FF",
		234562 => x"FF",
		234563 => x"FF",
		234564 => x"FF",
		234565 => x"FF",
		234566 => x"FF",
		234567 => x"FF",
		234568 => x"FF",
		234569 => x"FF",
		234570 => x"FF",
		234571 => x"FF",
		234572 => x"FF",
		234573 => x"FF",
		234574 => x"FF",
		234575 => x"FF",
		234576 => x"FF",
		234577 => x"FF",
		234578 => x"FF",
		234579 => x"FF",
		234580 => x"FF",
		234581 => x"FF",
		234582 => x"FF",
		234583 => x"FF",
		234584 => x"FF",
		234585 => x"FF",
		234586 => x"FF",
		234587 => x"FF",
		234588 => x"FF",
		234589 => x"FF",
		234590 => x"FF",
		234591 => x"FF",
		234592 => x"FF",
		234593 => x"FF",
		234594 => x"FF",
		234595 => x"FF",
		234596 => x"FF",
		234597 => x"FF",
		234598 => x"FF",
		234599 => x"FF",
		234600 => x"FF",
		234601 => x"FF",
		234602 => x"FF",
		234603 => x"FF",
		234604 => x"FF",
		234605 => x"FF",
		234606 => x"FF",
		234607 => x"FF",
		234608 => x"FF",
		234609 => x"FF",
		234610 => x"FF",
		234611 => x"FF",
		234612 => x"FF",
		234613 => x"FF",
		234614 => x"FF",
		234615 => x"FF",
		234616 => x"FF",
		234617 => x"FF",
		234618 => x"FF",
		234619 => x"FF",
		234620 => x"FF",
		234621 => x"FF",
		234622 => x"FF",
		234623 => x"FF",
		234624 => x"FF",
		234625 => x"FF",
		234626 => x"FF",
		234627 => x"FF",
		234628 => x"FF",
		234629 => x"FF",
		234630 => x"FF",
		234631 => x"FF",
		234632 => x"FF",
		234633 => x"FF",
		234634 => x"FF",
		234635 => x"FF",
		234636 => x"FF",
		234637 => x"FF",
		234638 => x"FF",
		234639 => x"FF",
		234640 => x"FF",
		234641 => x"FF",
		234642 => x"FF",
		234643 => x"FF",
		234644 => x"FF",
		234645 => x"FF",
		234646 => x"FF",
		234647 => x"FF",
		234648 => x"FF",
		234649 => x"FF",
		234650 => x"FF",
		234651 => x"FF",
		234652 => x"FF",
		234653 => x"FF",
		234654 => x"FF",
		234655 => x"FF",
		234656 => x"FF",
		234657 => x"FF",
		234658 => x"FF",
		234659 => x"FF",
		234660 => x"FF",
		234661 => x"FF",
		234662 => x"FF",
		234663 => x"FF",
		234664 => x"FF",
		234665 => x"FF",
		234666 => x"FF",
		234667 => x"FF",
		234668 => x"FF",
		234669 => x"FF",
		234670 => x"FF",
		234671 => x"FF",
		234672 => x"FF",
		234673 => x"FF",
		234674 => x"FF",
		234675 => x"FF",
		234676 => x"FF",
		234677 => x"FF",
		234678 => x"FF",
		234679 => x"FF",
		234680 => x"FF",
		234681 => x"FF",
		234682 => x"FF",
		234683 => x"FF",
		234684 => x"FF",
		234685 => x"FF",
		234686 => x"FF",
		234687 => x"FF",
		234688 => x"FF",
		234689 => x"FF",
		234690 => x"FF",
		234691 => x"FF",
		234692 => x"FF",
		234693 => x"FF",
		234694 => x"FF",
		234695 => x"FF",
		234696 => x"FF",
		234697 => x"FF",
		234698 => x"FF",
		234699 => x"FF",
		234700 => x"FF",
		234701 => x"FF",
		234702 => x"FF",
		234703 => x"FF",
		234704 => x"FF",
		234705 => x"FF",
		234706 => x"FF",
		234707 => x"FF",
		234708 => x"FF",
		234709 => x"FF",
		234710 => x"FF",
		234711 => x"FF",
		234712 => x"FF",
		234713 => x"FF",
		234714 => x"FF",
		234715 => x"FF",
		234716 => x"FF",
		234717 => x"FF",
		234718 => x"FF",
		234719 => x"FF",
		234720 => x"FF",
		234721 => x"FF",
		234722 => x"FF",
		234723 => x"FF",
		234724 => x"FF",
		234725 => x"FF",
		234726 => x"FF",
		234727 => x"FF",
		234728 => x"FF",
		234729 => x"FF",
		234730 => x"FF",
		234731 => x"FF",
		234732 => x"FF",
		234733 => x"FF",
		234734 => x"FF",
		234735 => x"FF",
		234736 => x"FF",
		234737 => x"FF",
		234738 => x"FF",
		234739 => x"FF",
		234740 => x"FF",
		234741 => x"FF",
		234742 => x"FF",
		234743 => x"FF",
		234744 => x"FF",
		234745 => x"FF",
		234746 => x"FF",
		234747 => x"FF",
		234748 => x"FF",
		234749 => x"FF",
		234750 => x"FF",
		234751 => x"FF",
		234752 => x"FF",
		234753 => x"FF",
		234754 => x"FF",
		234755 => x"FF",
		234756 => x"FF",
		234757 => x"FF",
		234758 => x"FF",
		234759 => x"FF",
		234760 => x"FF",
		234761 => x"FF",
		234762 => x"FF",
		234763 => x"FF",
		234764 => x"FF",
		234765 => x"FF",
		234766 => x"FF",
		234767 => x"FF",
		234768 => x"FF",
		234769 => x"FF",
		235564 => x"FF",
		235565 => x"FF",
		235566 => x"FF",
		235567 => x"FF",
		235568 => x"FF",
		235569 => x"FF",
		235570 => x"FF",
		235571 => x"FF",
		235572 => x"FF",
		235573 => x"FF",
		235574 => x"FF",
		235575 => x"FF",
		235576 => x"FF",
		235577 => x"FF",
		235578 => x"FF",
		235579 => x"FF",
		235580 => x"FF",
		235581 => x"FF",
		235582 => x"FF",
		235583 => x"FF",
		235584 => x"FF",
		235585 => x"FF",
		235586 => x"FF",
		235587 => x"FF",
		235588 => x"FF",
		235589 => x"FF",
		235590 => x"FF",
		235591 => x"FF",
		235592 => x"FF",
		235593 => x"FF",
		235594 => x"FF",
		235595 => x"FF",
		235596 => x"FF",
		235597 => x"FF",
		235598 => x"FF",
		235599 => x"FF",
		235600 => x"FF",
		235601 => x"FF",
		235602 => x"FF",
		235603 => x"FF",
		235604 => x"FF",
		235605 => x"FF",
		235606 => x"FF",
		235607 => x"FF",
		235608 => x"FF",
		235609 => x"FF",
		235610 => x"FF",
		235611 => x"FF",
		235612 => x"FF",
		235613 => x"FF",
		235614 => x"FF",
		235615 => x"FF",
		235616 => x"FF",
		235617 => x"FF",
		235618 => x"FF",
		235619 => x"FF",
		235620 => x"FF",
		235621 => x"FF",
		235622 => x"FF",
		235623 => x"FF",
		235624 => x"FF",
		235625 => x"FF",
		235626 => x"FF",
		235627 => x"FF",
		235628 => x"FF",
		235629 => x"FF",
		235630 => x"FF",
		235631 => x"FF",
		235632 => x"FF",
		235633 => x"FF",
		235634 => x"FF",
		235635 => x"FF",
		235636 => x"FF",
		235637 => x"FF",
		235638 => x"FF",
		235639 => x"FF",
		235640 => x"FF",
		235641 => x"FF",
		235642 => x"FF",
		235643 => x"FF",
		235644 => x"FF",
		235645 => x"FF",
		235646 => x"FF",
		235647 => x"FF",
		235648 => x"FF",
		235649 => x"FF",
		235650 => x"FF",
		235651 => x"FF",
		235652 => x"FF",
		235653 => x"FF",
		235654 => x"FF",
		235655 => x"FF",
		235656 => x"FF",
		235657 => x"FF",
		235658 => x"FF",
		235659 => x"FF",
		235660 => x"FF",
		235661 => x"FF",
		235662 => x"FF",
		235663 => x"FF",
		235664 => x"FF",
		235665 => x"FF",
		235666 => x"FF",
		235667 => x"FF",
		235668 => x"FF",
		235669 => x"FF",
		235670 => x"FF",
		235671 => x"FF",
		235672 => x"FF",
		235673 => x"FF",
		235674 => x"FF",
		235675 => x"FF",
		235676 => x"FF",
		235677 => x"FF",
		235678 => x"FF",
		235679 => x"FF",
		235680 => x"FF",
		235681 => x"FF",
		235682 => x"FF",
		235683 => x"FF",
		235684 => x"FF",
		235685 => x"FF",
		235686 => x"FF",
		235687 => x"FF",
		235688 => x"FF",
		235689 => x"FF",
		235690 => x"FF",
		235691 => x"FF",
		235692 => x"FF",
		235693 => x"FF",
		235694 => x"FF",
		235695 => x"FF",
		235696 => x"FF",
		235697 => x"FF",
		235698 => x"FF",
		235699 => x"FF",
		235700 => x"FF",
		235701 => x"FF",
		235702 => x"FF",
		235703 => x"FF",
		235704 => x"FF",
		235705 => x"FF",
		235706 => x"FF",
		235707 => x"FF",
		235708 => x"FF",
		235709 => x"FF",
		235710 => x"FF",
		235711 => x"FF",
		235712 => x"FF",
		235713 => x"FF",
		235714 => x"FF",
		235715 => x"FF",
		235716 => x"FF",
		235717 => x"FF",
		235718 => x"FF",
		235719 => x"FF",
		235720 => x"FF",
		235721 => x"FF",
		235722 => x"FF",
		235723 => x"FF",
		235724 => x"FF",
		235725 => x"FF",
		235726 => x"FF",
		235727 => x"FF",
		235728 => x"FF",
		235729 => x"FF",
		235730 => x"FF",
		235731 => x"FF",
		235732 => x"FF",
		235733 => x"FF",
		235734 => x"FF",
		235735 => x"FF",
		235736 => x"FF",
		235737 => x"FF",
		235738 => x"FF",
		235739 => x"FF",
		235740 => x"FF",
		235741 => x"FF",
		235742 => x"FF",
		235743 => x"FF",
		235744 => x"FF",
		235745 => x"FF",
		235746 => x"FF",
		235747 => x"FF",
		235748 => x"FF",
		235749 => x"FF",
		235750 => x"FF",
		235751 => x"FF",
		235752 => x"FF",
		235753 => x"FF",
		235754 => x"FF",
		235755 => x"FF",
		235756 => x"FF",
		235757 => x"FF",
		235758 => x"FF",
		235759 => x"FF",
		235760 => x"FF",
		235761 => x"FF",
		235762 => x"FF",
		235763 => x"FF",
		235764 => x"FF",
		235765 => x"FF",
		235766 => x"FF",
		235767 => x"FF",
		235768 => x"FF",
		235769 => x"FF",
		235770 => x"FF",
		235771 => x"FF",
		235772 => x"FF",
		235773 => x"FF",
		235774 => x"FF",
		235775 => x"FF",
		235776 => x"FF",
		235777 => x"FF",
		235778 => x"FF",
		235779 => x"FF",
		235780 => x"FF",
		235781 => x"FF",
		235782 => x"FF",
		235783 => x"FF",
		235784 => x"FF",
		235785 => x"FF",
		235786 => x"FF",
		235787 => x"FF",
		235788 => x"FF",
		235789 => x"FF",
		235790 => x"FF",
		235791 => x"FF",
		235792 => x"FF",
		235793 => x"FF",
		236588 => x"FF",
		236589 => x"FF",
		236590 => x"FF",
		236591 => x"FF",
		236592 => x"FF",
		236593 => x"FF",
		236594 => x"FF",
		236595 => x"FF",
		236596 => x"FF",
		236597 => x"FF",
		236598 => x"FF",
		236599 => x"FF",
		236600 => x"FF",
		236601 => x"FF",
		236602 => x"FF",
		236603 => x"FF",
		236604 => x"FF",
		236605 => x"FF",
		236606 => x"FF",
		236607 => x"FF",
		236608 => x"FF",
		236609 => x"FF",
		236610 => x"FF",
		236611 => x"FF",
		236612 => x"FF",
		236613 => x"FF",
		236614 => x"FF",
		236615 => x"FF",
		236616 => x"FF",
		236617 => x"FF",
		236618 => x"FF",
		236619 => x"FF",
		236620 => x"FF",
		236621 => x"FF",
		236622 => x"FF",
		236623 => x"FF",
		236624 => x"FF",
		236625 => x"FF",
		236626 => x"FF",
		236627 => x"FF",
		236628 => x"FF",
		236629 => x"FF",
		236630 => x"FF",
		236631 => x"FF",
		236632 => x"FF",
		236633 => x"FF",
		236634 => x"FF",
		236635 => x"FF",
		236636 => x"FF",
		236637 => x"FF",
		236638 => x"FF",
		236639 => x"FF",
		236640 => x"FF",
		236641 => x"FF",
		236642 => x"FF",
		236643 => x"FF",
		236644 => x"FF",
		236645 => x"FF",
		236646 => x"FF",
		236647 => x"FF",
		236648 => x"FF",
		236649 => x"FF",
		236650 => x"FF",
		236651 => x"FF",
		236652 => x"FF",
		236653 => x"FF",
		236654 => x"FF",
		236655 => x"FF",
		236656 => x"FF",
		236657 => x"FF",
		236658 => x"FF",
		236659 => x"FF",
		236660 => x"FF",
		236661 => x"FF",
		236662 => x"FF",
		236663 => x"FF",
		236664 => x"FF",
		236665 => x"FF",
		236666 => x"FF",
		236667 => x"FF",
		236668 => x"FF",
		236669 => x"FF",
		236670 => x"FF",
		236671 => x"FF",
		236672 => x"FF",
		236673 => x"FF",
		236674 => x"FF",
		236675 => x"FF",
		236676 => x"FF",
		236677 => x"FF",
		236678 => x"FF",
		236679 => x"FF",
		236680 => x"FF",
		236681 => x"FF",
		236682 => x"FF",
		236683 => x"FF",
		236684 => x"FF",
		236685 => x"FF",
		236686 => x"FF",
		236687 => x"FF",
		236688 => x"FF",
		236689 => x"FF",
		236690 => x"FF",
		236691 => x"FF",
		236692 => x"FF",
		236693 => x"FF",
		236694 => x"FF",
		236695 => x"FF",
		236696 => x"FF",
		236697 => x"FF",
		236698 => x"FF",
		236699 => x"FF",
		236700 => x"FF",
		236701 => x"FF",
		236702 => x"FF",
		236703 => x"FF",
		236704 => x"FF",
		236705 => x"FF",
		236706 => x"FF",
		236707 => x"FF",
		236708 => x"FF",
		236709 => x"FF",
		236710 => x"FF",
		236711 => x"FF",
		236712 => x"FF",
		236713 => x"FF",
		236714 => x"FF",
		236715 => x"FF",
		236716 => x"FF",
		236717 => x"FF",
		236718 => x"FF",
		236719 => x"FF",
		236720 => x"FF",
		236721 => x"FF",
		236722 => x"FF",
		236723 => x"FF",
		236724 => x"FF",
		236725 => x"FF",
		236726 => x"FF",
		236727 => x"FF",
		236728 => x"FF",
		236729 => x"FF",
		236730 => x"FF",
		236731 => x"FF",
		236732 => x"FF",
		236733 => x"FF",
		236734 => x"FF",
		236735 => x"FF",
		236736 => x"FF",
		236737 => x"FF",
		236738 => x"FF",
		236739 => x"FF",
		236740 => x"FF",
		236741 => x"FF",
		236742 => x"FF",
		236743 => x"FF",
		236744 => x"FF",
		236745 => x"FF",
		236746 => x"FF",
		236747 => x"FF",
		236748 => x"FF",
		236749 => x"FF",
		236750 => x"FF",
		236751 => x"FF",
		236752 => x"FF",
		236753 => x"FF",
		236754 => x"FF",
		236755 => x"FF",
		236756 => x"FF",
		236757 => x"FF",
		236758 => x"FF",
		236759 => x"FF",
		236760 => x"FF",
		236761 => x"FF",
		236762 => x"FF",
		236763 => x"FF",
		236764 => x"FF",
		236765 => x"FF",
		236766 => x"FF",
		236767 => x"FF",
		236768 => x"FF",
		236769 => x"FF",
		236770 => x"FF",
		236771 => x"FF",
		236772 => x"FF",
		236773 => x"FF",
		236774 => x"FF",
		236775 => x"FF",
		236776 => x"FF",
		236777 => x"FF",
		236778 => x"FF",
		236779 => x"FF",
		236780 => x"FF",
		236781 => x"FF",
		236782 => x"FF",
		236783 => x"FF",
		236784 => x"FF",
		236785 => x"FF",
		236786 => x"FF",
		236787 => x"FF",
		236788 => x"FF",
		236789 => x"FF",
		236790 => x"FF",
		236791 => x"FF",
		236792 => x"FF",
		236793 => x"FF",
		236794 => x"FF",
		236795 => x"FF",
		236796 => x"FF",
		236797 => x"FF",
		236798 => x"FF",
		236799 => x"FF",
		236800 => x"FF",
		236801 => x"FF",
		236802 => x"FF",
		236803 => x"FF",
		236804 => x"FF",
		236805 => x"FF",
		236806 => x"FF",
		236807 => x"FF",
		236808 => x"FF",
		236809 => x"FF",
		236810 => x"FF",
		236811 => x"FF",
		236812 => x"FF",
		236813 => x"FF",
		236814 => x"FF",
		236815 => x"FF",
		236816 => x"FF",
		236817 => x"FF",
		237612 => x"FF",
		237613 => x"FF",
		237614 => x"FF",
		237615 => x"FF",
		237616 => x"FF",
		237617 => x"FF",
		237618 => x"FF",
		237619 => x"FF",
		237620 => x"FF",
		237621 => x"FF",
		237622 => x"FF",
		237623 => x"FF",
		237624 => x"FF",
		237625 => x"FF",
		237626 => x"FF",
		237627 => x"FF",
		237628 => x"FF",
		237629 => x"FF",
		237630 => x"FF",
		237631 => x"FF",
		237632 => x"FF",
		237633 => x"FF",
		237634 => x"FF",
		237635 => x"FF",
		237636 => x"FF",
		237637 => x"FF",
		237638 => x"FF",
		237639 => x"FF",
		237640 => x"FF",
		237641 => x"FF",
		237642 => x"FF",
		237643 => x"FF",
		237644 => x"FF",
		237645 => x"FF",
		237646 => x"FF",
		237647 => x"FF",
		237648 => x"FF",
		237649 => x"FF",
		237650 => x"FF",
		237651 => x"FF",
		237652 => x"FF",
		237653 => x"FF",
		237654 => x"FF",
		237655 => x"FF",
		237656 => x"FF",
		237657 => x"FF",
		237658 => x"FF",
		237659 => x"FF",
		237660 => x"FF",
		237661 => x"FF",
		237662 => x"FF",
		237663 => x"FF",
		237664 => x"FF",
		237665 => x"FF",
		237666 => x"FF",
		237667 => x"FF",
		237668 => x"FF",
		237669 => x"FF",
		237670 => x"FF",
		237671 => x"FF",
		237672 => x"FF",
		237673 => x"FF",
		237674 => x"FF",
		237675 => x"FF",
		237676 => x"FF",
		237677 => x"FF",
		237678 => x"FF",
		237679 => x"FF",
		237680 => x"FF",
		237681 => x"FF",
		237682 => x"FF",
		237683 => x"FF",
		237684 => x"FF",
		237685 => x"FF",
		237686 => x"FF",
		237687 => x"FF",
		237688 => x"FF",
		237689 => x"FF",
		237690 => x"FF",
		237691 => x"FF",
		237692 => x"FF",
		237693 => x"FF",
		237694 => x"FF",
		237695 => x"FF",
		237696 => x"FF",
		237697 => x"FF",
		237698 => x"FF",
		237699 => x"FF",
		237700 => x"FF",
		237701 => x"FF",
		237702 => x"FF",
		237703 => x"FF",
		237704 => x"FF",
		237705 => x"FF",
		237706 => x"FF",
		237707 => x"FF",
		237708 => x"FF",
		237709 => x"FF",
		237710 => x"FF",
		237711 => x"FF",
		237712 => x"FF",
		237713 => x"FF",
		237714 => x"FF",
		237715 => x"FF",
		237716 => x"FF",
		237717 => x"FF",
		237718 => x"FF",
		237719 => x"FF",
		237720 => x"FF",
		237721 => x"FF",
		237722 => x"FF",
		237723 => x"FF",
		237724 => x"FF",
		237725 => x"FF",
		237726 => x"FF",
		237727 => x"FF",
		237728 => x"FF",
		237729 => x"FF",
		237730 => x"FF",
		237731 => x"FF",
		237732 => x"FF",
		237733 => x"FF",
		237734 => x"FF",
		237735 => x"FF",
		237736 => x"FF",
		237737 => x"FF",
		237738 => x"FF",
		237739 => x"FF",
		237740 => x"FF",
		237741 => x"FF",
		237742 => x"FF",
		237743 => x"FF",
		237744 => x"FF",
		237745 => x"FF",
		237746 => x"FF",
		237747 => x"FF",
		237748 => x"FF",
		237749 => x"FF",
		237750 => x"FF",
		237751 => x"FF",
		237752 => x"FF",
		237753 => x"FF",
		237754 => x"FF",
		237755 => x"FF",
		237756 => x"FF",
		237757 => x"FF",
		237758 => x"FF",
		237759 => x"FF",
		237760 => x"FF",
		237761 => x"FF",
		237762 => x"FF",
		237763 => x"FF",
		237764 => x"FF",
		237765 => x"FF",
		237766 => x"FF",
		237767 => x"FF",
		237768 => x"FF",
		237769 => x"FF",
		237770 => x"FF",
		237771 => x"FF",
		237772 => x"FF",
		237773 => x"FF",
		237774 => x"FF",
		237775 => x"FF",
		237776 => x"FF",
		237777 => x"FF",
		237778 => x"FF",
		237779 => x"FF",
		237780 => x"FF",
		237781 => x"FF",
		237782 => x"FF",
		237783 => x"FF",
		237784 => x"FF",
		237785 => x"FF",
		237786 => x"FF",
		237787 => x"FF",
		237788 => x"FF",
		237789 => x"FF",
		237790 => x"FF",
		237791 => x"FF",
		237792 => x"FF",
		237793 => x"FF",
		237794 => x"FF",
		237795 => x"FF",
		237796 => x"FF",
		237797 => x"FF",
		237798 => x"FF",
		237799 => x"FF",
		237800 => x"FF",
		237801 => x"FF",
		237802 => x"FF",
		237803 => x"FF",
		237804 => x"FF",
		237805 => x"FF",
		237806 => x"FF",
		237807 => x"FF",
		237808 => x"FF",
		237809 => x"FF",
		237810 => x"FF",
		237811 => x"FF",
		237812 => x"FF",
		237813 => x"FF",
		237814 => x"FF",
		237815 => x"FF",
		237816 => x"FF",
		237817 => x"FF",
		237818 => x"FF",
		237819 => x"FF",
		237820 => x"FF",
		237821 => x"FF",
		237822 => x"FF",
		237823 => x"FF",
		237824 => x"FF",
		237825 => x"FF",
		237826 => x"FF",
		237827 => x"FF",
		237828 => x"FF",
		237829 => x"FF",
		237830 => x"FF",
		237831 => x"FF",
		237832 => x"FF",
		237833 => x"FF",
		237834 => x"FF",
		237835 => x"FF",
		237836 => x"FF",
		237837 => x"FF",
		237838 => x"FF",
		237839 => x"FF",
		237840 => x"FF",
		237841 => x"FF",
		238636 => x"FF",
		238637 => x"FF",
		238638 => x"FF",
		238639 => x"FF",
		238640 => x"FF",
		238641 => x"FF",
		238642 => x"FF",
		238643 => x"FF",
		238644 => x"FF",
		238645 => x"FF",
		238646 => x"FF",
		238647 => x"FF",
		238648 => x"FF",
		238649 => x"FF",
		238650 => x"FF",
		238651 => x"FF",
		238652 => x"FF",
		238653 => x"FF",
		238654 => x"FF",
		238655 => x"FF",
		238656 => x"FF",
		238657 => x"FF",
		238658 => x"FF",
		238659 => x"FF",
		238660 => x"FF",
		238661 => x"FF",
		238662 => x"FF",
		238663 => x"FF",
		238664 => x"FF",
		238665 => x"FF",
		238666 => x"FF",
		238667 => x"FF",
		238668 => x"FF",
		238669 => x"FF",
		238670 => x"FF",
		238671 => x"FF",
		238672 => x"FF",
		238673 => x"FF",
		238674 => x"FF",
		238675 => x"FF",
		238676 => x"FF",
		238677 => x"FF",
		238678 => x"FF",
		238679 => x"FF",
		238680 => x"FF",
		238681 => x"FF",
		238682 => x"FF",
		238683 => x"FF",
		238684 => x"FF",
		238685 => x"FF",
		238686 => x"FF",
		238687 => x"FF",
		238688 => x"FF",
		238689 => x"FF",
		238690 => x"FF",
		238691 => x"FF",
		238692 => x"FF",
		238693 => x"FF",
		238694 => x"FF",
		238695 => x"FF",
		238696 => x"FF",
		238697 => x"FF",
		238698 => x"FF",
		238699 => x"FF",
		238700 => x"FF",
		238701 => x"FF",
		238702 => x"FF",
		238703 => x"FF",
		238704 => x"FF",
		238705 => x"FF",
		238706 => x"FF",
		238707 => x"FF",
		238708 => x"FF",
		238709 => x"FF",
		238710 => x"FF",
		238711 => x"FF",
		238712 => x"FF",
		238713 => x"FF",
		238714 => x"FF",
		238715 => x"FF",
		238716 => x"FF",
		238717 => x"FF",
		238718 => x"FF",
		238719 => x"FF",
		238720 => x"FF",
		238721 => x"FF",
		238722 => x"FF",
		238723 => x"FF",
		238724 => x"FF",
		238725 => x"FF",
		238726 => x"FF",
		238727 => x"FF",
		238728 => x"FF",
		238729 => x"FF",
		238730 => x"FF",
		238731 => x"FF",
		238732 => x"FF",
		238733 => x"FF",
		238734 => x"FF",
		238735 => x"FF",
		238736 => x"FF",
		238737 => x"FF",
		238738 => x"FF",
		238739 => x"FF",
		238740 => x"FF",
		238741 => x"FF",
		238742 => x"FF",
		238743 => x"FF",
		238744 => x"FF",
		238745 => x"FF",
		238746 => x"FF",
		238747 => x"FF",
		238748 => x"FF",
		238749 => x"FF",
		238750 => x"FF",
		238751 => x"FF",
		238752 => x"FF",
		238753 => x"FF",
		238754 => x"FF",
		238755 => x"FF",
		238756 => x"FF",
		238757 => x"FF",
		238758 => x"FF",
		238759 => x"FF",
		238760 => x"FF",
		238761 => x"FF",
		238762 => x"FF",
		238763 => x"FF",
		238764 => x"FF",
		238765 => x"FF",
		238766 => x"FF",
		238767 => x"FF",
		238768 => x"FF",
		238769 => x"FF",
		238770 => x"FF",
		238771 => x"FF",
		238772 => x"FF",
		238773 => x"FF",
		238774 => x"FF",
		238775 => x"FF",
		238776 => x"FF",
		238777 => x"FF",
		238778 => x"FF",
		238779 => x"FF",
		238780 => x"FF",
		238781 => x"FF",
		238782 => x"FF",
		238783 => x"FF",
		238784 => x"FF",
		238785 => x"FF",
		238786 => x"FF",
		238787 => x"FF",
		238788 => x"FF",
		238789 => x"FF",
		238790 => x"FF",
		238791 => x"FF",
		238792 => x"FF",
		238793 => x"FF",
		238794 => x"FF",
		238795 => x"FF",
		238796 => x"FF",
		238797 => x"FF",
		238798 => x"FF",
		238799 => x"FF",
		238800 => x"FF",
		238801 => x"FF",
		238802 => x"FF",
		238803 => x"FF",
		238804 => x"FF",
		238805 => x"FF",
		238806 => x"FF",
		238807 => x"FF",
		238808 => x"FF",
		238809 => x"FF",
		238810 => x"FF",
		238811 => x"FF",
		238812 => x"FF",
		238813 => x"FF",
		238814 => x"FF",
		238815 => x"FF",
		238816 => x"FF",
		238817 => x"FF",
		238818 => x"FF",
		238819 => x"FF",
		238820 => x"FF",
		238821 => x"FF",
		238822 => x"FF",
		238823 => x"FF",
		238824 => x"FF",
		238825 => x"FF",
		238826 => x"FF",
		238827 => x"FF",
		238828 => x"FF",
		238829 => x"FF",
		238830 => x"FF",
		238831 => x"FF",
		238832 => x"FF",
		238833 => x"FF",
		238834 => x"FF",
		238835 => x"FF",
		238836 => x"FF",
		238837 => x"FF",
		238838 => x"FF",
		238839 => x"FF",
		238840 => x"FF",
		238841 => x"FF",
		238842 => x"FF",
		238843 => x"FF",
		238844 => x"FF",
		238845 => x"FF",
		238846 => x"FF",
		238847 => x"FF",
		238848 => x"FF",
		238849 => x"FF",
		238850 => x"FF",
		238851 => x"FF",
		238852 => x"FF",
		238853 => x"FF",
		238854 => x"FF",
		238855 => x"FF",
		238856 => x"FF",
		238857 => x"FF",
		238858 => x"FF",
		238859 => x"FF",
		238860 => x"FF",
		238861 => x"FF",
		238862 => x"FF",
		238863 => x"FF",
		238864 => x"FF",
		238865 => x"FF",
