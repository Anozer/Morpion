0 => "00000000",
1 => "00000000",
2 => "00000000",
3 => "00000000",
4 => "00000000",
5 => "00000000",
6 => "00000000",
7 => "00000000",
8 => "00000000",
9 => "00000000",
10 => "00000000",
11 => "00000000",
12 => "00000000",
13 => "00000000",
14 => "00000000",
15 => "00000000",
16 => "00000000",
17 => "00000000",
18 => "00000000",
19 => "00000000",
20 => "00000000",
21 => "00000000",
22 => "00000000",
23 => "00000000",
24 => "00000000",
25 => "00000000",
26 => "00000000",
27 => "00001000",
28 => "00000000",
29 => "00000000",
30 => "00000000",
31 => "00000000",
32 => "00000000",
33 => "00000000",
34 => "00000000",
35 => "00000000",
36 => "00000000",
37 => "00000000",
38 => "00000000",
39 => "00000000",
40 => "00000000",
41 => "00000000",
42 => "00000000",
43 => "00000000",
44 => "00000000",
45 => "00000000",
46 => "00000000",
47 => "00000000",
48 => "00000000",
49 => "00000000",
50 => "00000000",
51 => "00000000",
52 => "00000000",
53 => "00000000",
54 => "00000000",
55 => "00000000",
56 => "00000000",
57 => "00000000",
58 => "00000000",
59 => "00000000",
60 => "00000000",
61 => "00000000",
62 => "00000000",
63 => "00000000",
64 => "00000000",
65 => "00000000",
66 => "00000000",
67 => "00000000",
68 => "00000000",
69 => "00000000",
70 => "00001000",
71 => "00000000",
72 => "00000000",
73 => "00000000",
74 => "00000000",
75 => "00000000",
76 => "00000000",
77 => "00001000",
78 => "00001000",
79 => "00000000",
80 => "00000000",
81 => "00000000",
82 => "00000000",
83 => "00000000",
84 => "00000000",
85 => "00000000",
86 => "00000000",
87 => "00000000",
88 => "00000000",
89 => "00000000",
90 => "00000000",
91 => "00000000",
92 => "00000000",
93 => "00000000",
94 => "00000000",
95 => "00000000",
96 => "00000000",
97 => "00000000",
98 => "00000000",
99 => "00000000",
100 => "00000000",
101 => "00000000",
102 => "00000000",
103 => "00000000",
104 => "00000000",
105 => "00000000",
106 => "00000000",
107 => "00000000",
108 => "00000000",
109 => "00000000",
110 => "00000000",
111 => "00000000",
112 => "00000000",
113 => "00000000",
114 => "00000000",
115 => "00000000",
116 => "00000000",
128 => "00000000",
129 => "00000000",
130 => "00000000",
131 => "00000000",
132 => "00000000",
133 => "00000000",
134 => "00000000",
135 => "00000000",
136 => "00000000",
137 => "00000000",
138 => "00000000",
139 => "00000000",
140 => "00000000",
141 => "00000000",
142 => "00000000",
143 => "00000000",
144 => "00000000",
145 => "00000000",
146 => "00000000",
147 => "00000000",
148 => "00000000",
149 => "00000000",
150 => "00000000",
151 => "00000000",
152 => "00000000",
153 => "00000000",
154 => "00000000",
155 => "00000000",
156 => "00000000",
157 => "00000000",
158 => "00000000",
159 => "00000000",
160 => "00000000",
161 => "00000000",
162 => "00000000",
163 => "00000000",
164 => "00000000",
165 => "00000000",
166 => "00000000",
167 => "00000000",
168 => "00000000",
169 => "00000000",
170 => "00000000",
171 => "00000000",
172 => "00000000",
173 => "00000000",
174 => "00000000",
175 => "00000000",
176 => "00000000",
177 => "00000000",
178 => "00000000",
179 => "00000000",
180 => "00000000",
181 => "00000000",
182 => "00000000",
183 => "00000000",
184 => "00000000",
185 => "00000000",
186 => "00000000",
187 => "00000000",
188 => "00000000",
189 => "00000000",
190 => "00000000",
191 => "00000000",
192 => "00000000",
193 => "00000000",
194 => "00000000",
195 => "00000000",
196 => "00000000",
197 => "00000000",
198 => "00000000",
199 => "00000000",
200 => "00000000",
201 => "00000000",
202 => "00000000",
203 => "00000000",
204 => "00000000",
205 => "00000000",
206 => "00000000",
207 => "00000000",
208 => "00000000",
209 => "00000000",
210 => "00000000",
211 => "00000000",
212 => "00000000",
213 => "00000000",
214 => "00000000",
215 => "00000000",
216 => "00000000",
217 => "00000000",
218 => "00000000",
219 => "00000000",
220 => "00000000",
221 => "00000000",
222 => "00000000",
223 => "00000000",
224 => "00000000",
225 => "00000000",
226 => "00000000",
227 => "00000000",
228 => "00000000",
229 => "00000000",
230 => "00000000",
231 => "00000000",
232 => "00000000",
233 => "00000000",
234 => "00000000",
235 => "00000000",
236 => "00000000",
237 => "00000000",
238 => "00000000",
239 => "00000000",
240 => "00000000",
241 => "00000000",
242 => "00000000",
243 => "00000000",
244 => "00000000",
256 => "00000000",
257 => "00000000",
258 => "00000000",
259 => "00000000",
260 => "00000000",
261 => "00000000",
262 => "00000000",
263 => "00000000",
264 => "00000000",
265 => "00000000",
266 => "00000000",
267 => "00000000",
268 => "00000000",
269 => "00000000",
270 => "00000000",
271 => "00000000",
272 => "00000000",
273 => "00000000",
274 => "00000000",
275 => "00000000",
276 => "00000000",
277 => "00000000",
278 => "00000000",
279 => "00000000",
280 => "00000000",
281 => "00000000",
282 => "00000000",
283 => "00000000",
284 => "00000000",
285 => "00000000",
286 => "00000000",
287 => "00000000",
288 => "00000000",
289 => "00000000",
290 => "00000000",
291 => "00000000",
292 => "00000000",
293 => "00000000",
294 => "00000000",
295 => "00000000",
296 => "00000000",
297 => "00000000",
298 => "00000000",
299 => "00000000",
300 => "00000000",
301 => "00000000",
302 => "00000000",
303 => "00000000",
304 => "00000000",
305 => "00000000",
306 => "00000000",
307 => "00000000",
308 => "00000000",
309 => "00000000",
310 => "00000000",
311 => "00000000",
312 => "00000000",
313 => "00000000",
314 => "00000000",
315 => "00000000",
316 => "00000000",
317 => "00000000",
318 => "00000000",
319 => "00000000",
320 => "00000000",
321 => "00000000",
322 => "00000000",
323 => "00000000",
324 => "00000000",
325 => "00000000",
326 => "00000000",
327 => "00000000",
328 => "00000000",
329 => "00000000",
330 => "00000000",
331 => "00000000",
332 => "00000000",
333 => "00000000",
334 => "00000000",
335 => "00000000",
336 => "00000000",
337 => "00000000",
338 => "00000000",
339 => "00000000",
340 => "00000000",
341 => "00000000",
342 => "00000000",
343 => "00000000",
344 => "00000000",
345 => "00000000",
346 => "00000000",
347 => "00000000",
348 => "00000000",
349 => "00000000",
350 => "00000000",
351 => "00000000",
352 => "00000000",
353 => "00000000",
354 => "00000000",
355 => "00000000",
356 => "00000000",
357 => "00000000",
358 => "00000000",
359 => "00000000",
360 => "00000000",
361 => "00000000",
362 => "00000000",
363 => "00000000",
364 => "00000000",
365 => "00000000",
366 => "00000000",
367 => "00000000",
368 => "00000000",
369 => "00000000",
370 => "00000000",
371 => "00000000",
372 => "00000000",
384 => "00000000",
385 => "00000000",
386 => "00000000",
387 => "00000000",
388 => "00000000",
389 => "00000000",
390 => "00000000",
391 => "00000000",
392 => "00000000",
393 => "00000000",
394 => "00000000",
395 => "00000000",
396 => "00000000",
397 => "00000000",
398 => "00000000",
399 => "00000000",
400 => "00000000",
401 => "00000000",
402 => "00000000",
403 => "00000000",
404 => "00000000",
405 => "00000000",
406 => "00000000",
407 => "00000000",
408 => "00000000",
409 => "00000000",
410 => "00000000",
411 => "00000000",
412 => "00000000",
413 => "00000000",
414 => "00000000",
415 => "00000000",
416 => "00000000",
417 => "00000000",
418 => "00000000",
419 => "00000000",
420 => "00000000",
421 => "00000000",
422 => "00000000",
423 => "00000000",
424 => "00000000",
425 => "00000000",
426 => "00000000",
427 => "00000000",
428 => "00000000",
429 => "00000000",
430 => "00000000",
431 => "00000000",
432 => "00000000",
433 => "00000000",
434 => "00000000",
435 => "00000000",
436 => "00000000",
437 => "00000000",
438 => "00000000",
439 => "00000000",
440 => "00000000",
441 => "00000000",
442 => "00000000",
443 => "00000000",
444 => "00000000",
445 => "00000000",
446 => "00000000",
447 => "00000000",
448 => "00000000",
449 => "00000000",
450 => "00001000",
451 => "00000000",
452 => "00000000",
453 => "00000000",
454 => "00000000",
455 => "00000000",
456 => "00000000",
457 => "00000000",
458 => "00000000",
459 => "00000000",
460 => "00000000",
461 => "00000000",
462 => "00000000",
463 => "00000000",
464 => "00000000",
465 => "00000000",
466 => "00000000",
467 => "00000000",
468 => "00000000",
469 => "00000000",
470 => "00000000",
471 => "00000000",
472 => "00000000",
473 => "00000000",
474 => "00000000",
475 => "00000000",
476 => "00000000",
477 => "00000000",
478 => "00000000",
479 => "00000000",
480 => "00000000",
481 => "00000000",
482 => "00000000",
483 => "00000000",
484 => "00000000",
485 => "00000000",
486 => "00000000",
487 => "00000000",
488 => "00000000",
489 => "00000000",
490 => "00000000",
491 => "00000000",
492 => "00000000",
493 => "00000000",
494 => "00000000",
495 => "00000000",
496 => "00000000",
497 => "00000000",
498 => "00000000",
499 => "00000000",
500 => "00000000",
512 => "00000000",
513 => "00000000",
514 => "00000000",
515 => "00000000",
516 => "00000000",
517 => "00000000",
518 => "00000000",
519 => "00000000",
520 => "00000000",
521 => "00000000",
522 => "00000000",
523 => "00000000",
524 => "00000000",
525 => "00000000",
526 => "00000000",
527 => "00000000",
528 => "00000000",
529 => "00000000",
530 => "00000000",
531 => "00000000",
532 => "00000000",
533 => "00000000",
534 => "00000000",
535 => "00000000",
536 => "00000000",
537 => "00000000",
538 => "00000000",
539 => "00000000",
540 => "00000000",
541 => "00000000",
542 => "00000000",
543 => "00000000",
544 => "00000000",
545 => "00000000",
546 => "00000000",
547 => "00000000",
548 => "00000000",
549 => "00000000",
550 => "00000000",
551 => "00000000",
552 => "00000000",
553 => "00000000",
554 => "00000000",
555 => "00000000",
556 => "00000000",
557 => "00000000",
558 => "00000000",
559 => "00000000",
560 => "00000000",
561 => "00000000",
562 => "00000000",
563 => "00000000",
564 => "00000000",
565 => "00000000",
566 => "00000000",
567 => "00000000",
568 => "00000000",
569 => "00000000",
570 => "00000000",
571 => "00000000",
572 => "00000000",
573 => "00000000",
574 => "00000000",
575 => "00000000",
576 => "00000000",
577 => "00000000",
578 => "00000000",
579 => "00000000",
580 => "00000000",
581 => "00000000",
582 => "00000000",
583 => "00000000",
584 => "00000000",
585 => "00000000",
586 => "00000000",
587 => "00000000",
588 => "00000000",
589 => "00000000",
590 => "00000000",
591 => "00000000",
592 => "00000000",
593 => "00000000",
594 => "00000000",
595 => "00000000",
596 => "00000000",
597 => "00000000",
598 => "00000000",
599 => "00000000",
600 => "00000000",
601 => "00000000",
602 => "00000000",
603 => "00000000",
604 => "00000000",
605 => "00000000",
606 => "00000000",
607 => "00000000",
608 => "00000000",
609 => "00000000",
610 => "00000000",
611 => "00000000",
612 => "00000000",
613 => "00000000",
614 => "00000000",
615 => "00000000",
616 => "00000000",
617 => "00000000",
618 => "00000000",
619 => "00000000",
620 => "00000000",
621 => "00000000",
622 => "00000000",
623 => "00000000",
624 => "00000000",
625 => "00000000",
626 => "00000000",
627 => "00000000",
628 => "00000000",
640 => "00000000",
641 => "00000000",
642 => "00000000",
643 => "00000000",
644 => "00000000",
645 => "00000000",
646 => "00000000",
647 => "00000000",
648 => "00000000",
649 => "00000000",
650 => "00000000",
651 => "00000000",
652 => "00000000",
653 => "00000000",
654 => "00000000",
655 => "00000000",
656 => "00000000",
657 => "00000000",
658 => "00000000",
659 => "00000000",
660 => "00000000",
661 => "00000000",
662 => "00000000",
663 => "00000000",
664 => "00000000",
665 => "00000000",
666 => "00000000",
667 => "00000000",
668 => "00000000",
669 => "00000000",
670 => "00000000",
671 => "00000000",
672 => "00000000",
673 => "00000000",
674 => "00000000",
675 => "00000000",
676 => "00000000",
677 => "00000000",
678 => "00000000",
679 => "00000000",
680 => "00000000",
681 => "00000000",
682 => "00000000",
683 => "00000000",
684 => "00000000",
685 => "00000000",
686 => "00000000",
687 => "00000000",
688 => "00000000",
689 => "00000000",
690 => "00000000",
691 => "00000000",
692 => "00000000",
693 => "00000000",
694 => "00000000",
695 => "00000000",
696 => "00000000",
697 => "00000000",
698 => "00000000",
699 => "00000000",
700 => "00000000",
701 => "00000000",
702 => "00000000",
703 => "00000000",
704 => "00000000",
705 => "00000000",
706 => "00000000",
707 => "00000000",
708 => "00000000",
709 => "00000000",
710 => "00000000",
711 => "00000000",
712 => "00000000",
713 => "00000000",
714 => "00000000",
715 => "00000000",
716 => "00000000",
717 => "00000000",
718 => "00000000",
719 => "00000000",
720 => "00000000",
721 => "00000000",
722 => "00000000",
723 => "00000000",
724 => "00000000",
725 => "00000000",
726 => "00000000",
727 => "00000000",
728 => "00000000",
729 => "00000000",
730 => "00000000",
731 => "00000000",
732 => "00000000",
733 => "00000000",
734 => "00000000",
735 => "00000000",
736 => "00000000",
737 => "00000000",
738 => "00000000",
739 => "00000000",
740 => "00000000",
741 => "00000000",
742 => "00000000",
743 => "00000000",
744 => "00000000",
745 => "00000000",
746 => "00000000",
747 => "00000000",
748 => "00000000",
749 => "00000000",
750 => "00000000",
751 => "00000000",
752 => "00000000",
753 => "00000000",
754 => "00000000",
755 => "00000000",
756 => "00000000",
768 => "00000000",
769 => "00000000",
770 => "00000000",
771 => "00000000",
772 => "00000000",
773 => "00000000",
774 => "00000000",
775 => "00000000",
776 => "00000000",
777 => "00000000",
778 => "00000000",
779 => "00000000",
780 => "00000000",
781 => "00000000",
782 => "00000000",
783 => "00000000",
784 => "00000000",
785 => "00000000",
786 => "00000000",
787 => "00000000",
788 => "00000000",
789 => "00000000",
790 => "00000000",
791 => "00000000",
792 => "00000000",
793 => "00000000",
794 => "00000000",
795 => "00000000",
796 => "00000000",
797 => "00000000",
798 => "00000000",
799 => "00000000",
800 => "00000000",
801 => "00000000",
802 => "00000000",
803 => "00000000",
804 => "00000000",
805 => "00000000",
806 => "00000000",
807 => "00000000",
808 => "00000000",
809 => "00000000",
810 => "00000000",
811 => "00000000",
812 => "00000000",
813 => "00000000",
814 => "00000000",
815 => "00000000",
816 => "00000000",
817 => "00000000",
818 => "00000000",
819 => "00000000",
820 => "00000000",
821 => "00000000",
822 => "00000000",
823 => "00000000",
824 => "00000000",
825 => "00000000",
826 => "00000000",
827 => "00000000",
828 => "00000000",
829 => "00000000",
830 => "00000000",
831 => "00000000",
832 => "00000000",
833 => "00000000",
834 => "00000000",
835 => "00000000",
836 => "00000000",
837 => "00000000",
838 => "00000000",
839 => "00000000",
840 => "00000000",
841 => "00000000",
842 => "00000000",
843 => "00000000",
844 => "00000000",
845 => "00000000",
846 => "00000000",
847 => "00000000",
848 => "00000000",
849 => "00000000",
850 => "00000000",
851 => "00000000",
852 => "00000000",
853 => "00000000",
854 => "00000000",
855 => "00000000",
856 => "00000000",
857 => "00000000",
858 => "00000000",
859 => "00000000",
860 => "00000000",
861 => "00000000",
862 => "00000000",
863 => "00000000",
864 => "00000000",
865 => "00000000",
866 => "00000000",
867 => "00000000",
868 => "00000000",
869 => "00000000",
870 => "00000000",
871 => "00000000",
872 => "00000000",
873 => "00000000",
874 => "00000000",
875 => "00000000",
876 => "00000000",
877 => "00000000",
878 => "00000000",
879 => "00000000",
880 => "00000000",
881 => "00000000",
882 => "00000000",
883 => "00000000",
884 => "00000000",
896 => "00000000",
897 => "00000000",
898 => "00000000",
899 => "00000000",
900 => "00000000",
901 => "00000000",
902 => "00000000",
903 => "00000000",
904 => "00000000",
905 => "00000000",
906 => "00000000",
907 => "00000000",
908 => "00000000",
909 => "00000000",
910 => "00000000",
911 => "00000000",
912 => "00000000",
913 => "00000000",
914 => "00000000",
915 => "00000000",
916 => "00000000",
917 => "00000000",
918 => "00000000",
919 => "00000000",
920 => "00000000",
921 => "00000000",
922 => "00000000",
923 => "00000000",
924 => "00000000",
925 => "00000000",
926 => "00000000",
927 => "00000000",
928 => "00000000",
929 => "00000000",
930 => "00000000",
931 => "00000000",
932 => "00000000",
933 => "00000000",
934 => "00000000",
935 => "00000000",
936 => "00000000",
937 => "00000000",
938 => "00000000",
939 => "00000000",
940 => "00000000",
941 => "00000000",
942 => "00000000",
943 => "00000000",
944 => "00000000",
945 => "00000000",
946 => "00000000",
947 => "00000000",
948 => "00000000",
949 => "00000000",
950 => "00000000",
951 => "00000000",
952 => "00000000",
953 => "00000000",
954 => "00000000",
955 => "00000000",
956 => "00000000",
957 => "00000000",
958 => "00000000",
959 => "00000000",
960 => "00000000",
961 => "00000000",
962 => "00000000",
963 => "00000000",
964 => "00000000",
965 => "00000000",
966 => "00000000",
967 => "00000000",
968 => "00000000",
969 => "00000000",
970 => "00000000",
971 => "00000000",
972 => "00000000",
973 => "00000000",
974 => "00000000",
975 => "00000000",
976 => "00000000",
977 => "00000000",
978 => "00000000",
979 => "00000000",
980 => "00000000",
981 => "00000000",
982 => "00000000",
983 => "00000000",
984 => "00000000",
985 => "00000000",
986 => "00000000",
987 => "00000000",
988 => "00000000",
989 => "00000000",
990 => "00000000",
991 => "00000000",
992 => "00000000",
993 => "00000000",
994 => "00000000",
995 => "00000000",
996 => "00000000",
997 => "00000000",
998 => "00000000",
999 => "00000000",
1000 => "00000000",
1001 => "00000000",
1002 => "00000000",
1003 => "00000000",
1004 => "00000000",
1005 => "00000000",
1006 => "00000000",
1007 => "00000000",
1008 => "00000000",
1009 => "00000000",
1010 => "00000000",
1011 => "00000000",
1012 => "00000000",
1024 => "00000000",
1025 => "00000000",
1026 => "00000000",
1027 => "00000000",
1028 => "00000000",
1029 => "00000000",
1030 => "00000000",
1031 => "00000000",
1032 => "00000000",
1033 => "00000000",
1034 => "00000000",
1035 => "00000000",
1036 => "00000000",
1037 => "00000000",
1038 => "00000000",
1039 => "00000000",
1040 => "00000000",
1041 => "00000000",
1042 => "00000000",
1043 => "00000000",
1044 => "00000000",
1045 => "00000000",
1046 => "00000000",
1047 => "00000000",
1048 => "00000000",
1049 => "00000000",
1050 => "00000000",
1051 => "00000000",
1052 => "00000000",
1053 => "00000000",
1054 => "00000000",
1055 => "00000000",
1056 => "00000000",
1057 => "00000000",
1058 => "00000000",
1059 => "00000000",
1060 => "00000000",
1061 => "00000000",
1062 => "00000000",
1063 => "00000000",
1064 => "00000000",
1065 => "00000000",
1066 => "00000000",
1067 => "00000000",
1068 => "00000000",
1069 => "00000000",
1070 => "00000000",
1071 => "00000000",
1072 => "00000000",
1073 => "00000000",
1074 => "00000000",
1075 => "00000000",
1076 => "00000000",
1077 => "00000000",
1078 => "00000000",
1079 => "00000000",
1080 => "00000000",
1081 => "00000000",
1082 => "00000000",
1083 => "00000000",
1084 => "00000000",
1085 => "00000000",
1086 => "00000000",
1087 => "00000000",
1088 => "00000000",
1089 => "00000000",
1090 => "00000000",
1091 => "00000000",
1092 => "00000000",
1093 => "00000000",
1094 => "00000000",
1095 => "00000000",
1096 => "00000000",
1097 => "00000000",
1098 => "00000000",
1099 => "00000000",
1100 => "00000000",
1101 => "00000000",
1102 => "00000000",
1103 => "00000000",
1104 => "00000000",
1105 => "00000000",
1106 => "00000000",
1107 => "00000000",
1108 => "00000000",
1109 => "00000000",
1110 => "00000000",
1111 => "00000000",
1112 => "00000000",
1113 => "00000000",
1114 => "00000000",
1115 => "00000000",
1116 => "00000000",
1117 => "00000000",
1118 => "00000000",
1119 => "00000000",
1120 => "00000000",
1121 => "00000000",
1122 => "00000000",
1123 => "00000000",
1124 => "00000000",
1125 => "00000000",
1126 => "00000000",
1127 => "00000000",
1128 => "00000000",
1129 => "00000000",
1130 => "00000000",
1131 => "00000000",
1132 => "00000000",
1133 => "00000000",
1134 => "00000000",
1135 => "00000000",
1136 => "00000000",
1137 => "00000000",
1138 => "00000000",
1139 => "00000000",
1140 => "00000000",
1152 => "00000000",
1153 => "00000000",
1154 => "00000000",
1155 => "00000000",
1156 => "00000000",
1157 => "00000000",
1158 => "00000000",
1159 => "00000000",
1160 => "00000000",
1161 => "00000000",
1162 => "00000000",
1163 => "00000000",
1164 => "00000000",
1165 => "00000000",
1166 => "00000000",
1167 => "00000000",
1168 => "00000000",
1169 => "00000000",
1170 => "00000000",
1171 => "00000000",
1172 => "00000000",
1173 => "00000000",
1174 => "00000000",
1175 => "00000000",
1176 => "00000000",
1177 => "00000000",
1178 => "00000000",
1179 => "00000000",
1180 => "00000000",
1181 => "00000000",
1182 => "00000000",
1183 => "00000000",
1184 => "00000000",
1185 => "00000000",
1186 => "00000000",
1187 => "00000000",
1188 => "00000000",
1189 => "00000000",
1190 => "00000000",
1191 => "00000000",
1192 => "00000000",
1193 => "00000000",
1194 => "00000000",
1195 => "00000000",
1196 => "00000000",
1197 => "00000000",
1198 => "00000000",
1199 => "00000000",
1200 => "00000000",
1201 => "00000000",
1202 => "00000000",
1203 => "00000000",
1204 => "00000000",
1205 => "00000000",
1206 => "00000000",
1207 => "00000000",
1208 => "00000000",
1209 => "00000000",
1210 => "00000000",
1211 => "00000000",
1212 => "00000000",
1213 => "00000000",
1214 => "00000000",
1215 => "00000000",
1216 => "00000000",
1217 => "00000000",
1218 => "00000000",
1219 => "00000000",
1220 => "00000000",
1221 => "00000000",
1222 => "00000000",
1223 => "00000000",
1224 => "00000000",
1225 => "00000000",
1226 => "00000000",
1227 => "00000000",
1228 => "00000000",
1229 => "00000000",
1230 => "00000000",
1231 => "00000000",
1232 => "00000000",
1233 => "00000000",
1234 => "00000000",
1235 => "00000000",
1236 => "00000000",
1237 => "00000000",
1238 => "00000000",
1239 => "00000000",
1240 => "00000000",
1241 => "00000000",
1242 => "00000000",
1243 => "00000000",
1244 => "00000000",
1245 => "00000000",
1246 => "00000000",
1247 => "00000000",
1248 => "00000000",
1249 => "00000000",
1250 => "00000000",
1251 => "00000000",
1252 => "00000000",
1253 => "00000000",
1254 => "00000000",
1255 => "00000000",
1256 => "00000000",
1257 => "00000000",
1258 => "00000000",
1259 => "00000000",
1260 => "00000000",
1261 => "00000000",
1262 => "00000000",
1263 => "00000000",
1264 => "00000000",
1265 => "00000000",
1266 => "00000000",
1267 => "00000000",
1268 => "00000000",
1280 => "00000000",
1281 => "00000000",
1282 => "00000000",
1283 => "00000000",
1284 => "00000000",
1285 => "00000000",
1286 => "00000000",
1287 => "00000000",
1288 => "00000000",
1289 => "00000000",
1290 => "00000000",
1291 => "00000000",
1292 => "00000000",
1293 => "00000000",
1294 => "00000000",
1295 => "00000000",
1296 => "00000000",
1297 => "00000000",
1298 => "00000000",
1299 => "00000000",
1300 => "00000000",
1301 => "00000000",
1302 => "00000000",
1303 => "00000000",
1304 => "00000000",
1305 => "00000000",
1306 => "00000000",
1307 => "00000000",
1308 => "00000000",
1309 => "00000000",
1310 => "00000000",
1311 => "00000000",
1312 => "00000000",
1313 => "00000000",
1314 => "00000000",
1315 => "00000000",
1316 => "00000000",
1317 => "00000000",
1318 => "00000000",
1319 => "00000000",
1320 => "00000000",
1321 => "00000000",
1322 => "00000000",
1323 => "00000000",
1324 => "00000000",
1325 => "00000000",
1326 => "00000000",
1327 => "00000000",
1328 => "00000000",
1329 => "00000000",
1330 => "00000000",
1331 => "00000000",
1332 => "00000000",
1333 => "00000000",
1334 => "00000000",
1335 => "00000000",
1336 => "00000000",
1337 => "00000000",
1338 => "00000000",
1339 => "00000000",
1340 => "00000000",
1341 => "00000000",
1342 => "00000000",
1343 => "00000000",
1344 => "00000000",
1345 => "00000000",
1346 => "00000000",
1347 => "00000000",
1348 => "00000000",
1349 => "00000000",
1350 => "00000000",
1351 => "00000000",
1352 => "00000000",
1353 => "00000000",
1354 => "00000000",
1355 => "00000000",
1356 => "00000000",
1357 => "00000000",
1358 => "00000000",
1359 => "00000000",
1360 => "00000000",
1361 => "00000000",
1362 => "00000000",
1363 => "00000000",
1364 => "00000000",
1365 => "00000000",
1366 => "00000000",
1367 => "00000000",
1368 => "00000000",
1369 => "00000000",
1370 => "00000000",
1371 => "00000000",
1372 => "00000000",
1373 => "00000000",
1374 => "00000000",
1375 => "00000000",
1376 => "00000000",
1377 => "00000000",
1378 => "00000000",
1379 => "00000000",
1380 => "00000000",
1381 => "00000000",
1382 => "00000000",
1383 => "00000000",
1384 => "00000000",
1385 => "00000000",
1386 => "00000000",
1387 => "00000000",
1388 => "00000000",
1389 => "00000000",
1390 => "00000000",
1391 => "00000000",
1392 => "00000000",
1393 => "00000000",
1394 => "00000000",
1395 => "00000000",
1396 => "00000000",
1408 => "00000000",
1409 => "00000000",
1410 => "00000000",
1411 => "00000000",
1412 => "00000000",
1413 => "00000000",
1414 => "00000000",
1415 => "00000000",
1416 => "00000000",
1417 => "00000000",
1418 => "00000000",
1419 => "00000000",
1420 => "00000000",
1421 => "00000000",
1422 => "00000000",
1423 => "00000000",
1424 => "00000000",
1425 => "00000000",
1426 => "00000000",
1427 => "00000000",
1428 => "00000000",
1429 => "00000000",
1430 => "00000000",
1431 => "00000000",
1432 => "00000000",
1433 => "00000000",
1434 => "00000000",
1435 => "00000000",
1436 => "00000000",
1437 => "00000000",
1438 => "00000000",
1439 => "00000000",
1440 => "00000000",
1441 => "00000000",
1442 => "00000000",
1443 => "00000000",
1444 => "00000000",
1445 => "00000000",
1446 => "00000000",
1447 => "00000000",
1448 => "00000000",
1449 => "00000000",
1450 => "00000000",
1451 => "00000000",
1452 => "00000000",
1453 => "00000000",
1454 => "00000000",
1455 => "00000000",
1456 => "00000000",
1457 => "00000000",
1458 => "00000000",
1459 => "00000000",
1460 => "00000000",
1461 => "00000000",
1462 => "00000000",
1463 => "00000000",
1464 => "00000000",
1465 => "00000000",
1466 => "00000000",
1467 => "00000000",
1468 => "00000000",
1469 => "00000000",
1470 => "00000000",
1471 => "00000000",
1472 => "00000000",
1473 => "00000000",
1474 => "00000000",
1475 => "00000000",
1476 => "00000000",
1477 => "00000000",
1478 => "00000000",
1479 => "00000000",
1480 => "00000000",
1481 => "00000000",
1482 => "00000000",
1483 => "00000000",
1484 => "00000000",
1485 => "00000000",
1486 => "00000000",
1487 => "00000000",
1488 => "00000000",
1489 => "00000000",
1490 => "00000000",
1491 => "00000000",
1492 => "00000000",
1493 => "00000000",
1494 => "00000000",
1495 => "00000000",
1496 => "00000000",
1497 => "00000000",
1498 => "00000000",
1499 => "00000000",
1500 => "00000000",
1501 => "00000000",
1502 => "00000000",
1503 => "00000000",
1504 => "00000000",
1505 => "00000000",
1506 => "00000000",
1507 => "00000000",
1508 => "00000000",
1509 => "00000000",
1510 => "00000000",
1511 => "00000000",
1512 => "00000000",
1513 => "00000000",
1514 => "00000000",
1515 => "00000000",
1516 => "00000000",
1517 => "00000000",
1518 => "00000000",
1519 => "00000000",
1520 => "00000000",
1521 => "00000000",
1522 => "00000000",
1523 => "00000000",
1524 => "00000000",
1536 => "00000000",
1537 => "00000000",
1538 => "00000000",
1539 => "00000000",
1540 => "00000000",
1541 => "00000000",
1542 => "00000000",
1543 => "00000000",
1544 => "00000000",
1545 => "00000000",
1546 => "00000000",
1547 => "00000000",
1548 => "00000000",
1549 => "00000000",
1550 => "00000000",
1551 => "00000000",
1552 => "00000000",
1553 => "00000000",
1554 => "00000000",
1555 => "00000000",
1556 => "00000000",
1557 => "00000000",
1558 => "00000000",
1559 => "00000000",
1560 => "00000000",
1561 => "00000000",
1562 => "00000000",
1563 => "00000000",
1564 => "00000000",
1565 => "00000000",
1566 => "00000000",
1567 => "00000000",
1568 => "00000000",
1569 => "00000000",
1570 => "00000000",
1571 => "00000000",
1572 => "00000000",
1573 => "00000000",
1574 => "00000000",
1575 => "00000000",
1576 => "00000000",
1577 => "00000000",
1578 => "00000000",
1579 => "00000000",
1580 => "00000000",
1581 => "00000000",
1582 => "00000000",
1583 => "00000000",
1584 => "00000000",
1585 => "00000000",
1586 => "00000000",
1587 => "00000000",
1588 => "00000000",
1589 => "00000000",
1590 => "00000000",
1591 => "00000000",
1592 => "00000000",
1593 => "00000000",
1594 => "00000000",
1595 => "00000000",
1596 => "00000000",
1597 => "00000000",
1598 => "00000000",
1599 => "00000000",
1600 => "00000000",
1601 => "00000000",
1602 => "00000000",
1603 => "00000000",
1604 => "00000000",
1605 => "00000000",
1606 => "00000000",
1607 => "00000000",
1608 => "00000000",
1609 => "00000000",
1610 => "00000000",
1611 => "00000000",
1612 => "00000000",
1613 => "00000000",
1614 => "00000000",
1615 => "00000000",
1616 => "00000000",
1617 => "00000000",
1618 => "00000000",
1619 => "00000000",
1620 => "00000000",
1621 => "00000000",
1622 => "00000000",
1623 => "00000000",
1624 => "00000000",
1625 => "00000000",
1626 => "00000000",
1627 => "00000000",
1628 => "00000000",
1629 => "00000000",
1630 => "00000000",
1631 => "00000000",
1632 => "00000000",
1633 => "00000000",
1634 => "00000000",
1635 => "00000000",
1636 => "00000000",
1637 => "00000000",
1638 => "00000000",
1639 => "00000000",
1640 => "00000000",
1641 => "00000000",
1642 => "00000000",
1643 => "00000000",
1644 => "00000000",
1645 => "00000000",
1646 => "00000000",
1647 => "00000000",
1648 => "00000000",
1649 => "00000000",
1650 => "00000000",
1651 => "00000000",
1652 => "00000000",
1664 => "00000000",
1665 => "00000000",
1666 => "00000000",
1667 => "00000000",
1668 => "00000000",
1669 => "00000000",
1670 => "00000000",
1671 => "00000000",
1672 => "00000000",
1673 => "00000000",
1674 => "00000000",
1675 => "00000000",
1676 => "00000000",
1677 => "00000000",
1678 => "00000000",
1679 => "00000000",
1680 => "00000000",
1681 => "00000000",
1682 => "00000000",
1683 => "00000000",
1684 => "00000000",
1685 => "00000000",
1686 => "00000000",
1687 => "00000000",
1688 => "00000000",
1689 => "00000000",
1690 => "00000000",
1691 => "00000000",
1692 => "00000000",
1693 => "00000000",
1694 => "00000000",
1695 => "00000000",
1696 => "00000000",
1697 => "00000000",
1698 => "00000000",
1699 => "00000000",
1700 => "00000000",
1701 => "00000000",
1702 => "00000000",
1703 => "00000000",
1704 => "00000000",
1705 => "00000000",
1706 => "00000000",
1707 => "00000000",
1708 => "00000000",
1709 => "00000000",
1710 => "00000000",
1711 => "00000000",
1712 => "00000000",
1713 => "00000000",
1714 => "00000000",
1715 => "00000000",
1716 => "00000000",
1717 => "00000000",
1718 => "00000000",
1719 => "00000000",
1720 => "00000000",
1721 => "00000000",
1722 => "00000000",
1723 => "00000000",
1724 => "00000000",
1725 => "00000000",
1726 => "00000000",
1727 => "00000000",
1728 => "00000000",
1729 => "00000000",
1730 => "00000000",
1731 => "00000000",
1732 => "00000000",
1733 => "00000000",
1734 => "00000000",
1735 => "00000000",
1736 => "00000000",
1737 => "00000000",
1738 => "00000000",
1739 => "00000000",
1740 => "00000000",
1741 => "00000000",
1742 => "00000000",
1743 => "00000000",
1744 => "00000000",
1745 => "00000000",
1746 => "00000000",
1747 => "00000000",
1748 => "00000000",
1749 => "00000000",
1750 => "00000000",
1751 => "00000000",
1752 => "00000000",
1753 => "00000000",
1754 => "00000000",
1755 => "00000000",
1756 => "00000000",
1757 => "00000000",
1758 => "00000000",
1759 => "00000000",
1760 => "00000000",
1761 => "00000000",
1762 => "00000000",
1763 => "00000000",
1764 => "00000000",
1765 => "00000000",
1766 => "00000000",
1767 => "00000000",
1768 => "00000000",
1769 => "00000000",
1770 => "00000000",
1771 => "00000000",
1772 => "00000000",
1773 => "00000000",
1774 => "00000000",
1775 => "00000000",
1776 => "00000000",
1777 => "00000000",
1778 => "00000000",
1779 => "00000000",
1780 => "00000000",
1792 => "00000000",
1793 => "00000000",
1794 => "00000000",
1795 => "00000000",
1796 => "00000000",
1797 => "00000000",
1798 => "00000000",
1799 => "00000000",
1800 => "00000000",
1801 => "00000000",
1802 => "00000000",
1803 => "00000000",
1804 => "00000000",
1805 => "00000000",
1806 => "00000000",
1807 => "00000000",
1808 => "00000000",
1809 => "00000000",
1810 => "00000000",
1811 => "00000000",
1812 => "00000000",
1813 => "00000000",
1814 => "00000000",
1815 => "00000000",
1816 => "00000000",
1817 => "00000000",
1818 => "00000000",
1819 => "00000000",
1820 => "00000000",
1821 => "00000000",
1822 => "00000000",
1823 => "00000000",
1824 => "00000000",
1825 => "00000000",
1826 => "00000000",
1827 => "00000000",
1828 => "00000000",
1829 => "00000000",
1830 => "00000000",
1831 => "00000000",
1832 => "00000000",
1833 => "00000000",
1834 => "00000000",
1835 => "00000000",
1836 => "00000000",
1837 => "00000000",
1838 => "00000000",
1839 => "00000000",
1840 => "00000000",
1841 => "00000000",
1842 => "00000000",
1843 => "00000000",
1844 => "00000000",
1845 => "00000000",
1846 => "00000000",
1847 => "00000000",
1848 => "00000000",
1849 => "00000000",
1850 => "00000000",
1851 => "00000000",
1852 => "00000000",
1853 => "00000000",
1854 => "00000000",
1855 => "00000000",
1856 => "00000000",
1857 => "00000000",
1858 => "00000000",
1859 => "00000000",
1860 => "00000000",
1861 => "00000000",
1862 => "00000000",
1863 => "00000000",
1864 => "00000000",
1865 => "00000000",
1866 => "00000000",
1867 => "00000000",
1868 => "00000000",
1869 => "00000000",
1870 => "00000000",
1871 => "00000000",
1872 => "00000000",
1873 => "00000000",
1874 => "00000000",
1875 => "00000000",
1876 => "00000000",
1877 => "00000000",
1878 => "00000000",
1879 => "00000000",
1880 => "00000000",
1881 => "00000000",
1882 => "00000000",
1883 => "00000000",
1884 => "00000000",
1885 => "00000000",
1886 => "00000000",
1887 => "00000000",
1888 => "00000000",
1889 => "00000000",
1890 => "00000000",
1891 => "00000000",
1892 => "00000000",
1893 => "00000000",
1894 => "00000000",
1895 => "00000000",
1896 => "00000000",
1897 => "00000000",
1898 => "00000000",
1899 => "00000000",
1900 => "00000000",
1901 => "00000000",
1902 => "00000000",
1903 => "00000000",
1904 => "00000000",
1905 => "00000000",
1906 => "00000000",
1907 => "00000000",
1908 => "00000000",
1920 => "00000000",
1921 => "00000000",
1922 => "00000000",
1923 => "00000000",
1924 => "00000000",
1925 => "00000000",
1926 => "00000000",
1927 => "00000000",
1928 => "00000000",
1929 => "00000000",
1930 => "00000000",
1931 => "00000000",
1932 => "00000000",
1933 => "00000000",
1934 => "00000000",
1935 => "00000000",
1936 => "00000000",
1937 => "00000000",
1938 => "00000000",
1939 => "00000000",
1940 => "00000000",
1941 => "00000000",
1942 => "00000000",
1943 => "00000000",
1944 => "00000000",
1945 => "00000000",
1946 => "00000000",
1947 => "00000000",
1948 => "00000000",
1949 => "00000000",
1950 => "00000000",
1951 => "00000000",
1952 => "00000000",
1953 => "00000000",
1954 => "00000000",
1955 => "00000000",
1956 => "00000000",
1957 => "00000000",
1958 => "00000000",
1959 => "00000000",
1960 => "00000000",
1961 => "00000000",
1962 => "00000000",
1963 => "00000000",
1964 => "00000000",
1965 => "00000000",
1966 => "00000000",
1967 => "00000000",
1968 => "00000000",
1969 => "00000000",
1970 => "00000000",
1971 => "00000000",
1972 => "00000000",
1973 => "00000000",
1974 => "00000000",
1975 => "00000000",
1976 => "00000000",
1977 => "00000000",
1978 => "00000000",
1979 => "00000000",
1980 => "00000000",
1981 => "00000000",
1982 => "00000000",
1983 => "00000000",
1984 => "00000000",
1985 => "00000000",
1986 => "00000000",
1987 => "00000000",
1988 => "00000000",
1989 => "00000000",
1990 => "00000000",
1991 => "00000000",
1992 => "00000000",
1993 => "00000000",
1994 => "00000000",
1995 => "00000000",
1996 => "00000000",
1997 => "00000000",
1998 => "00000000",
1999 => "00000000",
2000 => "00000000",
2001 => "00000000",
2002 => "00000000",
2003 => "00000000",
2004 => "00000000",
2005 => "00000000",
2006 => "00000000",
2007 => "00000000",
2008 => "00000000",
2009 => "00000000",
2010 => "00000000",
2011 => "00000000",
2012 => "00000000",
2013 => "00000000",
2014 => "00000000",
2015 => "00000000",
2016 => "00000000",
2017 => "00000000",
2018 => "00000000",
2019 => "00000000",
2020 => "00000000",
2021 => "00000000",
2022 => "00000000",
2023 => "00000000",
2024 => "00000000",
2025 => "00000000",
2026 => "00000000",
2027 => "00000000",
2028 => "00000000",
2029 => "00000000",
2030 => "00000000",
2031 => "00000000",
2032 => "00000000",
2033 => "00000000",
2034 => "00000000",
2035 => "00000000",
2036 => "00000000",
2048 => "00000000",
2049 => "00000000",
2050 => "00000000",
2051 => "00000000",
2052 => "00000000",
2053 => "00000000",
2054 => "00000000",
2055 => "00000000",
2056 => "00000000",
2057 => "00000000",
2058 => "00000000",
2059 => "00000000",
2060 => "00000000",
2061 => "00000000",
2062 => "00000000",
2063 => "00000000",
2064 => "00000000",
2065 => "00000000",
2066 => "00000000",
2067 => "00000000",
2068 => "00000000",
2069 => "00000000",
2070 => "00000000",
2071 => "00000000",
2072 => "00000000",
2073 => "00000000",
2074 => "00000000",
2075 => "00000000",
2076 => "00000000",
2077 => "00000000",
2078 => "00000000",
2079 => "00000000",
2080 => "00000000",
2081 => "00000000",
2082 => "00000000",
2083 => "00000000",
2084 => "00000000",
2085 => "00000000",
2086 => "00000000",
2087 => "00000000",
2088 => "00000000",
2089 => "00000000",
2090 => "00000000",
2091 => "00000000",
2092 => "00000000",
2093 => "00000000",
2094 => "00000000",
2095 => "00000000",
2096 => "00000000",
2097 => "00000000",
2098 => "00000000",
2099 => "00000000",
2100 => "00000000",
2101 => "00000000",
2102 => "00000000",
2103 => "00000000",
2104 => "00000000",
2105 => "00000000",
2106 => "00000000",
2107 => "00000000",
2108 => "00000000",
2109 => "00000000",
2110 => "00000000",
2111 => "00000000",
2112 => "00000000",
2113 => "00000000",
2114 => "00000000",
2115 => "00000000",
2116 => "00000000",
2117 => "00000000",
2118 => "00000000",
2119 => "00000000",
2120 => "00000000",
2121 => "00000000",
2122 => "00000000",
2123 => "00000000",
2124 => "00000000",
2125 => "00000000",
2126 => "00000000",
2127 => "00000000",
2128 => "00000000",
2129 => "00000000",
2130 => "00000000",
2131 => "00000000",
2132 => "00000000",
2133 => "00000000",
2134 => "00000000",
2135 => "00000000",
2136 => "00000000",
2137 => "00000000",
2138 => "00000000",
2139 => "00000000",
2140 => "00000000",
2141 => "00000000",
2142 => "00000000",
2143 => "00000000",
2144 => "00000000",
2145 => "00000000",
2146 => "00000000",
2147 => "00000000",
2148 => "00000000",
2149 => "00000000",
2150 => "00000000",
2151 => "00000000",
2152 => "00000000",
2153 => "00000000",
2154 => "00000000",
2155 => "00000000",
2156 => "00000000",
2157 => "00000000",
2158 => "00000000",
2159 => "00000000",
2160 => "00000000",
2161 => "00000000",
2162 => "00000000",
2163 => "00000000",
2164 => "00000000",
2176 => "00000000",
2177 => "00000000",
2178 => "00000000",
2179 => "00000000",
2180 => "00000000",
2181 => "00000000",
2182 => "00000000",
2183 => "00000000",
2184 => "00000000",
2185 => "00000000",
2186 => "00000000",
2187 => "00000000",
2188 => "00000000",
2189 => "00000000",
2190 => "00000000",
2191 => "00000000",
2192 => "00000000",
2193 => "00000000",
2194 => "00000000",
2195 => "00000000",
2196 => "00000000",
2197 => "00000000",
2198 => "00000000",
2199 => "00000000",
2200 => "00000000",
2201 => "00000000",
2202 => "00000000",
2203 => "00000000",
2204 => "00000000",
2205 => "00000000",
2206 => "00000000",
2207 => "00000000",
2208 => "00000000",
2209 => "00000000",
2210 => "00000000",
2211 => "00000000",
2212 => "00000000",
2213 => "00000000",
2214 => "00000000",
2215 => "00000000",
2216 => "00000000",
2217 => "00000000",
2218 => "00000000",
2219 => "00000000",
2220 => "00000000",
2221 => "00000000",
2222 => "00000000",
2223 => "00000000",
2224 => "00000000",
2225 => "00000000",
2226 => "00000000",
2227 => "00000000",
2228 => "00000000",
2229 => "00000000",
2230 => "00000000",
2231 => "00000000",
2232 => "00000000",
2233 => "00000000",
2234 => "00000000",
2235 => "00000000",
2236 => "00000000",
2237 => "00000000",
2238 => "00000000",
2239 => "00000000",
2240 => "00000000",
2241 => "00000000",
2242 => "00000000",
2243 => "00000000",
2244 => "00000000",
2245 => "00000000",
2246 => "00000000",
2247 => "00000000",
2248 => "00000000",
2249 => "00000000",
2250 => "00000000",
2251 => "00000000",
2252 => "00000000",
2253 => "00000000",
2254 => "00000000",
2255 => "00000000",
2256 => "00000000",
2257 => "00000000",
2258 => "00000000",
2259 => "00000000",
2260 => "00000000",
2261 => "00000000",
2262 => "00000000",
2263 => "00000000",
2264 => "00000000",
2265 => "00000000",
2266 => "00000000",
2267 => "00000000",
2268 => "00000000",
2269 => "00000000",
2270 => "00000000",
2271 => "00000000",
2272 => "00000000",
2273 => "00000000",
2274 => "00000000",
2275 => "00000000",
2276 => "00000000",
2277 => "00000000",
2278 => "00000000",
2279 => "00000000",
2280 => "00000000",
2281 => "00000000",
2282 => "00000000",
2283 => "00000000",
2284 => "00000000",
2285 => "00000000",
2286 => "00000000",
2287 => "00000000",
2288 => "00000000",
2289 => "00000000",
2290 => "00000000",
2291 => "00000000",
2292 => "00000000",
2304 => "00000000",
2305 => "00000000",
2306 => "00000000",
2307 => "00000000",
2308 => "00000000",
2309 => "00000000",
2310 => "00000000",
2311 => "00000000",
2312 => "00000000",
2313 => "00000000",
2314 => "00000000",
2315 => "00000000",
2316 => "00000000",
2317 => "00000000",
2318 => "00000000",
2319 => "00000000",
2320 => "00000000",
2321 => "00000000",
2322 => "00000000",
2323 => "00000000",
2324 => "00000000",
2325 => "00000000",
2326 => "00000000",
2327 => "00000000",
2328 => "00000000",
2329 => "00000000",
2330 => "00000000",
2331 => "00000000",
2332 => "00000000",
2333 => "00000000",
2334 => "00000000",
2335 => "00000000",
2336 => "00000000",
2337 => "00000000",
2338 => "00000000",
2339 => "00000000",
2340 => "00000000",
2341 => "00000000",
2342 => "00000000",
2343 => "00000000",
2344 => "00000000",
2345 => "00000000",
2346 => "00000000",
2347 => "00000000",
2348 => "00000000",
2349 => "00000000",
2350 => "00000000",
2351 => "00000000",
2352 => "00000000",
2353 => "00000000",
2354 => "00000000",
2355 => "00000000",
2356 => "00000000",
2357 => "00000000",
2358 => "00000000",
2359 => "00000000",
2360 => "00000000",
2361 => "00000000",
2362 => "00000000",
2363 => "00000000",
2364 => "00000000",
2365 => "00000000",
2366 => "00000000",
2367 => "00000000",
2368 => "00000000",
2369 => "00000000",
2370 => "00000000",
2371 => "00000000",
2372 => "00000000",
2373 => "00000000",
2374 => "00000000",
2375 => "00000000",
2376 => "00000000",
2377 => "00000000",
2378 => "00000000",
2379 => "00000000",
2380 => "00000000",
2381 => "00000000",
2382 => "00000000",
2383 => "00000000",
2384 => "00000000",
2385 => "00000000",
2386 => "00000000",
2387 => "00000000",
2388 => "00000000",
2389 => "00000000",
2390 => "00000000",
2391 => "00000000",
2392 => "00000000",
2393 => "00000000",
2394 => "00000000",
2395 => "00000000",
2396 => "00000000",
2397 => "00000000",
2398 => "00000000",
2399 => "00000000",
2400 => "00000000",
2401 => "00000000",
2402 => "00000000",
2403 => "00000000",
2404 => "00000000",
2405 => "00000000",
2406 => "00000000",
2407 => "00000000",
2408 => "00000000",
2409 => "00000000",
2410 => "00000000",
2411 => "00000000",
2412 => "00000000",
2413 => "00000000",
2414 => "00000000",
2415 => "00000000",
2416 => "00000000",
2417 => "00000000",
2418 => "00000000",
2419 => "00000000",
2420 => "00000000",
2432 => "00000000",
2433 => "00000000",
2434 => "00000000",
2435 => "00000000",
2436 => "00000000",
2437 => "00000000",
2438 => "00000000",
2439 => "00000000",
2440 => "00000000",
2441 => "00000000",
2442 => "00000000",
2443 => "00000000",
2444 => "00000000",
2445 => "00000000",
2446 => "00000000",
2447 => "00000000",
2448 => "00000000",
2449 => "00000000",
2450 => "00000000",
2451 => "00000000",
2452 => "00000000",
2453 => "00000000",
2454 => "00000000",
2455 => "00000000",
2456 => "00000000",
2457 => "00000000",
2458 => "00000000",
2459 => "00000000",
2460 => "00000000",
2461 => "00000000",
2462 => "00000000",
2463 => "00000000",
2464 => "00000000",
2465 => "00000000",
2466 => "00000000",
2467 => "00000000",
2468 => "00000000",
2469 => "00000000",
2470 => "00000000",
2471 => "00000000",
2472 => "00000000",
2473 => "00000000",
2474 => "00000000",
2475 => "00000000",
2476 => "00000000",
2477 => "00000000",
2478 => "00000000",
2479 => "00000000",
2480 => "00000000",
2481 => "00000000",
2482 => "00000000",
2483 => "00000000",
2484 => "00000000",
2485 => "00000000",
2486 => "00000000",
2487 => "00000000",
2488 => "00000000",
2489 => "00000000",
2490 => "00000000",
2491 => "00000000",
2492 => "00000000",
2493 => "00000000",
2494 => "00000000",
2495 => "00000000",
2496 => "00000000",
2497 => "00000000",
2498 => "00000000",
2499 => "00000000",
2500 => "00000000",
2501 => "00000000",
2502 => "00000000",
2503 => "00000000",
2504 => "00000000",
2505 => "00000000",
2506 => "00000000",
2507 => "00000000",
2508 => "00000000",
2509 => "00000000",
2510 => "00000000",
2511 => "00000000",
2512 => "00000000",
2513 => "00000000",
2514 => "00000000",
2515 => "00000000",
2516 => "00000000",
2517 => "00000000",
2518 => "00000000",
2519 => "00000000",
2520 => "00000000",
2521 => "00000000",
2522 => "00000000",
2523 => "00000000",
2524 => "00000000",
2525 => "00000000",
2526 => "00000000",
2527 => "00000000",
2528 => "00000000",
2529 => "00000000",
2530 => "00000000",
2531 => "00000000",
2532 => "00000000",
2533 => "00000000",
2534 => "00000000",
2535 => "00000000",
2536 => "00000000",
2537 => "00000000",
2538 => "00000000",
2539 => "00000000",
2540 => "00000000",
2541 => "00000000",
2542 => "00000000",
2543 => "00000000",
2544 => "00000000",
2545 => "00000000",
2546 => "00000000",
2547 => "00000000",
2548 => "00000000",
2560 => "00000000",
2561 => "00000000",
2562 => "00000000",
2563 => "00000000",
2564 => "00000000",
2565 => "00000000",
2566 => "00000000",
2567 => "00000000",
2568 => "00000000",
2569 => "00000000",
2570 => "00000000",
2571 => "00000000",
2572 => "00000000",
2573 => "00000000",
2574 => "00000000",
2575 => "00000000",
2576 => "00000000",
2577 => "00000000",
2578 => "00000000",
2579 => "00000000",
2580 => "00000000",
2581 => "00000000",
2582 => "00000000",
2583 => "00000000",
2584 => "00000000",
2585 => "00000000",
2586 => "00000000",
2587 => "00000000",
2588 => "00000000",
2589 => "00000000",
2590 => "00000000",
2591 => "00000000",
2592 => "00000000",
2593 => "00000000",
2594 => "00000000",
2595 => "00000000",
2596 => "00000000",
2597 => "00000000",
2598 => "00000000",
2599 => "00000000",
2600 => "00000000",
2601 => "00000000",
2602 => "00000000",
2603 => "00000000",
2604 => "00000000",
2605 => "00000000",
2606 => "00000000",
2607 => "00000000",
2608 => "00000000",
2609 => "00000000",
2610 => "00000000",
2611 => "00000000",
2612 => "00000000",
2613 => "00000000",
2614 => "00000000",
2615 => "00000000",
2616 => "00000000",
2617 => "00000000",
2618 => "00000000",
2619 => "00000000",
2620 => "00000000",
2621 => "00000000",
2622 => "00000000",
2623 => "00000000",
2624 => "00000000",
2625 => "00000000",
2626 => "00000000",
2627 => "00000000",
2628 => "00000000",
2629 => "00000000",
2630 => "00000000",
2631 => "00000000",
2632 => "00000000",
2633 => "00000000",
2634 => "00000000",
2635 => "00000000",
2636 => "00000000",
2637 => "00000000",
2638 => "00000000",
2639 => "00000000",
2640 => "00000000",
2641 => "00000000",
2642 => "00000000",
2643 => "00000000",
2644 => "00000000",
2645 => "00000000",
2646 => "00000000",
2647 => "00000000",
2648 => "00000000",
2649 => "00000000",
2650 => "00000000",
2651 => "00000000",
2652 => "00000000",
2653 => "00000000",
2654 => "00000000",
2655 => "00000000",
2656 => "00000000",
2657 => "00000000",
2658 => "00000000",
2659 => "00000000",
2660 => "00000000",
2661 => "00000000",
2662 => "00000000",
2663 => "00000000",
2664 => "00000000",
2665 => "00000000",
2666 => "00000000",
2667 => "00000000",
2668 => "00000000",
2669 => "00000000",
2670 => "00000000",
2671 => "00000000",
2672 => "00000000",
2673 => "00000000",
2674 => "00000000",
2675 => "00000000",
2676 => "00000000",
2688 => "00000000",
2689 => "00000000",
2690 => "00000000",
2691 => "00000000",
2692 => "00000000",
2693 => "00000000",
2694 => "00000000",
2695 => "00000000",
2696 => "00000000",
2697 => "00000000",
2698 => "00000000",
2699 => "00000000",
2700 => "00000000",
2701 => "00000000",
2702 => "00000000",
2703 => "00000000",
2704 => "00000000",
2705 => "00000000",
2706 => "00000000",
2707 => "00000000",
2708 => "00000000",
2709 => "00000000",
2710 => "00000000",
2711 => "00000000",
2712 => "00000000",
2713 => "00000000",
2714 => "00000000",
2715 => "00000000",
2716 => "00000000",
2717 => "00000000",
2718 => "00000000",
2719 => "00000000",
2720 => "00000000",
2721 => "00000000",
2722 => "00000000",
2723 => "00000000",
2724 => "00000000",
2725 => "00000000",
2726 => "00000000",
2727 => "00000000",
2728 => "00000000",
2729 => "00000000",
2730 => "00000000",
2731 => "00000000",
2732 => "00000000",
2733 => "00000000",
2734 => "00000000",
2735 => "00000000",
2736 => "00000000",
2737 => "00000000",
2738 => "00000000",
2739 => "00000000",
2740 => "00000000",
2741 => "00000000",
2742 => "00000000",
2743 => "00000000",
2744 => "00000000",
2745 => "00000000",
2746 => "00000000",
2747 => "00000000",
2748 => "00000000",
2749 => "00000000",
2750 => "00000000",
2751 => "00000000",
2752 => "00000000",
2753 => "00000000",
2754 => "00000000",
2755 => "00000000",
2756 => "00000000",
2757 => "00000000",
2758 => "00000000",
2759 => "00000000",
2760 => "00000000",
2761 => "00000000",
2762 => "00000000",
2763 => "00000000",
2764 => "00000000",
2765 => "00000000",
2766 => "00000000",
2767 => "00000000",
2768 => "00000000",
2769 => "00000000",
2770 => "00000000",
2771 => "00000000",
2772 => "00000000",
2773 => "00000000",
2774 => "00000000",
2775 => "00000000",
2776 => "00000000",
2777 => "00000000",
2778 => "00000000",
2779 => "00000000",
2780 => "00000000",
2781 => "00000000",
2782 => "00000000",
2783 => "00000000",
2784 => "00000000",
2785 => "00000000",
2786 => "00000000",
2787 => "00000000",
2788 => "00000000",
2789 => "00000000",
2790 => "00000000",
2791 => "00000000",
2792 => "00000000",
2793 => "00000000",
2794 => "00000000",
2795 => "00000000",
2796 => "00000000",
2797 => "00000000",
2798 => "00000000",
2799 => "00000000",
2800 => "00000000",
2801 => "00000000",
2802 => "00000000",
2803 => "00000000",
2804 => "00000000",
2816 => "00000000",
2817 => "00000000",
2818 => "00000000",
2819 => "00000000",
2820 => "00000000",
2821 => "00000000",
2822 => "00000000",
2823 => "00000000",
2824 => "00000000",
2825 => "00000000",
2826 => "00000000",
2827 => "00000000",
2828 => "00000000",
2829 => "00000000",
2830 => "00000000",
2831 => "00000000",
2832 => "00000000",
2833 => "00000000",
2834 => "00000000",
2835 => "00000000",
2836 => "00000000",
2837 => "00000000",
2838 => "00000000",
2839 => "00000000",
2840 => "00000000",
2841 => "00000000",
2842 => "00000000",
2843 => "00000000",
2844 => "00000000",
2845 => "00000000",
2846 => "00000000",
2847 => "00000000",
2848 => "00000000",
2849 => "00000000",
2850 => "00000000",
2851 => "00000000",
2852 => "00000000",
2853 => "00000000",
2854 => "00000000",
2855 => "00000000",
2856 => "00000000",
2857 => "00000000",
2858 => "00000000",
2859 => "00000000",
2860 => "00000000",
2861 => "00000000",
2862 => "00000000",
2863 => "00000000",
2864 => "00000000",
2865 => "00000000",
2866 => "00000000",
2867 => "00000000",
2868 => "00000000",
2869 => "00000000",
2870 => "00000000",
2871 => "00000000",
2872 => "00000000",
2873 => "00000000",
2874 => "00000000",
2875 => "00000000",
2876 => "00000000",
2877 => "00000000",
2878 => "00000000",
2879 => "00000000",
2880 => "00000000",
2881 => "00000000",
2882 => "00000000",
2883 => "00000000",
2884 => "00000000",
2885 => "00000000",
2886 => "00000000",
2887 => "00000000",
2888 => "00000000",
2889 => "00000000",
2890 => "00000000",
2891 => "00000000",
2892 => "00000000",
2893 => "00000000",
2894 => "00000000",
2895 => "00000000",
2896 => "00000000",
2897 => "00000000",
2898 => "00000000",
2899 => "00000000",
2900 => "00000000",
2901 => "00000000",
2902 => "00000000",
2903 => "00000000",
2904 => "00000000",
2905 => "00000000",
2906 => "00000000",
2907 => "00000000",
2908 => "00000000",
2909 => "00000000",
2910 => "00000000",
2911 => "00000000",
2912 => "00000000",
2913 => "00000000",
2914 => "00000000",
2915 => "00000000",
2916 => "00000000",
2917 => "00000000",
2918 => "00000000",
2919 => "00000000",
2920 => "00000000",
2921 => "00000000",
2922 => "00000000",
2923 => "00000000",
2924 => "00000000",
2925 => "00000000",
2926 => "00000000",
2927 => "00000000",
2928 => "00000000",
2929 => "00000000",
2930 => "00000000",
2931 => "00000000",
2932 => "00000000",
2944 => "00000000",
2945 => "00000000",
2946 => "00000000",
2947 => "00000000",
2948 => "00000000",
2949 => "00000000",
2950 => "00000000",
2951 => "00000000",
2952 => "00000000",
2953 => "00000000",
2954 => "00000000",
2955 => "00000000",
2956 => "00000000",
2957 => "00000000",
2958 => "00000000",
2959 => "00000000",
2960 => "00000000",
2961 => "00000000",
2962 => "00000000",
2963 => "00000000",
2964 => "00000000",
2965 => "00000000",
2966 => "00000000",
2967 => "00000000",
2968 => "00000000",
2969 => "00000000",
2970 => "00000000",
2971 => "00000000",
2972 => "00000000",
2973 => "00000000",
2974 => "00000000",
2975 => "00000000",
2976 => "00000000",
2977 => "00000000",
2978 => "00000000",
2979 => "00000000",
2980 => "00000000",
2981 => "00000000",
2982 => "00000000",
2983 => "00000000",
2984 => "00000000",
2985 => "00000000",
2986 => "00000000",
2987 => "00000000",
2988 => "00000000",
2989 => "00000000",
2990 => "00000000",
2991 => "00000000",
2992 => "00000000",
2993 => "00000000",
2994 => "00000000",
2995 => "00000000",
2996 => "00000000",
2997 => "00000000",
2998 => "00000000",
2999 => "00000000",
3000 => "00000000",
3001 => "00000000",
3002 => "00000000",
3003 => "00000000",
3004 => "00000000",
3005 => "00000000",
3006 => "00000000",
3007 => "00000000",
3008 => "00000000",
3009 => "00000000",
3010 => "00000000",
3011 => "00000000",
3012 => "00000000",
3013 => "00000000",
3014 => "00000000",
3015 => "00000000",
3016 => "00000000",
3017 => "00000000",
3018 => "00000000",
3019 => "00000000",
3020 => "00000000",
3021 => "00000000",
3022 => "00000000",
3023 => "00000000",
3024 => "00000000",
3025 => "00000000",
3026 => "00000000",
3027 => "00000000",
3028 => "00000000",
3029 => "00000000",
3030 => "00000000",
3031 => "00000000",
3032 => "00000000",
3033 => "00000000",
3034 => "00000000",
3035 => "00000000",
3036 => "00000000",
3037 => "00000000",
3038 => "00000000",
3039 => "00000000",
3040 => "00000000",
3041 => "00000000",
3042 => "00000000",
3043 => "00000000",
3044 => "00000000",
3045 => "00000000",
3046 => "00000000",
3047 => "00000000",
3048 => "00000000",
3049 => "00000000",
3050 => "00000000",
3051 => "00000000",
3052 => "00000000",
3053 => "00000000",
3054 => "00000000",
3055 => "00000000",
3056 => "00000000",
3057 => "00000000",
3058 => "00000000",
3059 => "00000000",
3060 => "00000000",
3072 => "00000000",
3073 => "00000000",
3074 => "00000000",
3075 => "00000000",
3076 => "00000000",
3077 => "00000000",
3078 => "00000000",
3079 => "00000000",
3080 => "00000000",
3081 => "00000000",
3082 => "00000000",
3083 => "00000000",
3084 => "00000000",
3085 => "00000000",
3086 => "00000000",
3087 => "00000000",
3088 => "00000000",
3089 => "00000000",
3090 => "00000000",
3091 => "00000000",
3092 => "00000000",
3093 => "00000000",
3094 => "00000000",
3095 => "00000000",
3096 => "00000000",
3097 => "00000000",
3098 => "00000000",
3099 => "00000000",
3100 => "00000000",
3101 => "00000000",
3102 => "00000000",
3103 => "00000000",
3104 => "00000000",
3105 => "00000000",
3106 => "00000000",
3107 => "00000000",
3108 => "00000000",
3109 => "00000000",
3110 => "00000000",
3111 => "00000000",
3112 => "00000000",
3113 => "00000000",
3114 => "00000000",
3115 => "00000000",
3116 => "00000000",
3117 => "00000000",
3118 => "00000000",
3119 => "00000000",
3120 => "00000000",
3121 => "00000000",
3122 => "00000000",
3123 => "00000000",
3124 => "00000000",
3125 => "00000000",
3126 => "00000000",
3127 => "00000000",
3128 => "00000000",
3129 => "00000000",
3130 => "00000000",
3131 => "00000000",
3132 => "00000000",
3133 => "00000000",
3134 => "00000000",
3135 => "00000000",
3136 => "00000000",
3137 => "00000000",
3138 => "00000000",
3139 => "00000000",
3140 => "00000000",
3141 => "00000000",
3142 => "00000000",
3143 => "00000000",
3144 => "00000000",
3145 => "00000000",
3146 => "00000000",
3147 => "00000000",
3148 => "00000000",
3149 => "00000000",
3150 => "00000000",
3151 => "00000000",
3152 => "00000000",
3153 => "00000000",
3154 => "00000000",
3155 => "00000000",
3156 => "00000000",
3157 => "00000000",
3158 => "00000000",
3159 => "00000000",
3160 => "00000000",
3161 => "00000000",
3162 => "00000000",
3163 => "00000000",
3164 => "00000000",
3165 => "00000000",
3166 => "00000000",
3167 => "00000000",
3168 => "00000000",
3169 => "00000000",
3170 => "00000000",
3171 => "00000000",
3172 => "00000000",
3173 => "00000000",
3174 => "00000000",
3175 => "00000000",
3176 => "00000000",
3177 => "00000000",
3178 => "00000000",
3179 => "00000000",
3180 => "00000000",
3181 => "00000000",
3182 => "00000000",
3183 => "00000000",
3184 => "00000000",
3185 => "00000000",
3186 => "00000000",
3187 => "00000000",
3188 => "00000000",
3200 => "00000000",
3201 => "00000000",
3202 => "00000000",
3203 => "00000000",
3204 => "00000000",
3205 => "00000000",
3206 => "00000000",
3207 => "00000000",
3208 => "00000000",
3209 => "00000000",
3210 => "00000000",
3211 => "00000000",
3212 => "00000000",
3213 => "00000000",
3214 => "00000000",
3215 => "00000000",
3216 => "00000000",
3217 => "00000000",
3218 => "00000000",
3219 => "00000000",
3220 => "00000000",
3221 => "00000000",
3222 => "00000000",
3223 => "00000000",
3224 => "00000000",
3225 => "00000000",
3226 => "00000000",
3227 => "00000000",
3228 => "00000000",
3229 => "00000000",
3230 => "00000000",
3231 => "00000000",
3232 => "00000000",
3233 => "00000000",
3234 => "00000000",
3235 => "00000000",
3236 => "00000000",
3237 => "00000000",
3238 => "00000000",
3239 => "00000000",
3240 => "00000000",
3241 => "00000000",
3242 => "00000000",
3243 => "00000000",
3244 => "00000000",
3245 => "00000000",
3246 => "00000000",
3247 => "00000000",
3248 => "00000000",
3249 => "00000000",
3250 => "00000000",
3251 => "00000000",
3252 => "00000000",
3253 => "00000000",
3254 => "00000000",
3255 => "00000000",
3256 => "00000000",
3257 => "00000000",
3258 => "00000000",
3259 => "00000000",
3260 => "00000000",
3261 => "00000000",
3262 => "00000000",
3263 => "00000000",
3264 => "00000000",
3265 => "00000000",
3266 => "00000000",
3267 => "00000000",
3268 => "00000000",
3269 => "00000000",
3270 => "00000000",
3271 => "00000000",
3272 => "00000000",
3273 => "00000000",
3274 => "00000000",
3275 => "00000000",
3276 => "00000000",
3277 => "00000000",
3278 => "00000000",
3279 => "00000000",
3280 => "00000000",
3281 => "00000000",
3282 => "00000000",
3283 => "00000000",
3284 => "00000000",
3285 => "00000000",
3286 => "00000000",
3287 => "00000000",
3288 => "00000000",
3289 => "00000000",
3290 => "00000000",
3291 => "00000000",
3292 => "00000000",
3293 => "00000000",
3294 => "00000000",
3295 => "00000000",
3296 => "00000000",
3297 => "00000000",
3298 => "00000000",
3299 => "00000000",
3300 => "00000000",
3301 => "00000000",
3302 => "00000000",
3303 => "00000000",
3304 => "00000000",
3305 => "00000000",
3306 => "00000000",
3307 => "00000000",
3308 => "00000000",
3309 => "00000000",
3310 => "00000000",
3311 => "00000000",
3312 => "00000000",
3313 => "00000000",
3314 => "00000000",
3315 => "00000000",
3316 => "00000000",
3328 => "00000000",
3329 => "00000000",
3330 => "00000000",
3331 => "00000000",
3332 => "00000000",
3333 => "00000000",
3334 => "00000000",
3335 => "00000000",
3336 => "00000000",
3337 => "00000000",
3338 => "00000000",
3339 => "00000000",
3340 => "00000000",
3341 => "00000000",
3342 => "00000000",
3343 => "00000000",
3344 => "00000000",
3345 => "00000000",
3346 => "00000000",
3347 => "00000000",
3348 => "00000000",
3349 => "00000000",
3350 => "00000000",
3351 => "00000000",
3352 => "00000000",
3353 => "00000000",
3354 => "00000000",
3355 => "00000000",
3356 => "00000000",
3357 => "00000000",
3358 => "00000000",
3359 => "00000000",
3360 => "00000000",
3361 => "00000000",
3362 => "00000000",
3363 => "00000000",
3364 => "00000000",
3365 => "00000000",
3366 => "00000000",
3367 => "00000000",
3368 => "00000000",
3369 => "00000000",
3370 => "00000000",
3371 => "00000000",
3372 => "00000000",
3373 => "00000000",
3374 => "00000000",
3375 => "00000000",
3376 => "00000000",
3377 => "00000000",
3378 => "00000000",
3379 => "00000000",
3380 => "00000000",
3381 => "00000000",
3382 => "00000000",
3383 => "00000000",
3384 => "00000000",
3385 => "00000000",
3386 => "00000000",
3387 => "00000000",
3388 => "00000000",
3389 => "00000000",
3390 => "00000000",
3391 => "00000000",
3392 => "00000000",
3393 => "00000000",
3394 => "00000000",
3395 => "00000000",
3396 => "00000000",
3397 => "00000000",
3398 => "00000000",
3399 => "00000000",
3400 => "00000000",
3401 => "00000000",
3402 => "00000000",
3403 => "00000000",
3404 => "00000000",
3405 => "00000000",
3406 => "00000000",
3407 => "00000000",
3408 => "00000000",
3409 => "00000000",
3410 => "00000000",
3411 => "00000000",
3412 => "00000000",
3413 => "00000000",
3414 => "00000000",
3415 => "00000000",
3416 => "00000000",
3417 => "00000000",
3418 => "00000000",
3419 => "00000000",
3420 => "00000000",
3421 => "00000000",
3422 => "00000000",
3423 => "00000000",
3424 => "00000000",
3425 => "00000000",
3426 => "00000000",
3427 => "00000000",
3428 => "00000000",
3429 => "00000000",
3430 => "00000000",
3431 => "00000000",
3432 => "00000000",
3433 => "00000000",
3434 => "00000000",
3435 => "00000000",
3436 => "00000000",
3437 => "00000000",
3438 => "00000000",
3439 => "00000000",
3440 => "00000000",
3441 => "00000000",
3442 => "00000000",
3443 => "00000000",
3444 => "00000000",
3456 => "00000000",
3457 => "00000000",
3458 => "00000000",
3459 => "00000000",
3460 => "00000000",
3461 => "00000000",
3462 => "00000000",
3463 => "00000000",
3464 => "00000000",
3465 => "00000000",
3466 => "00000000",
3467 => "00000000",
3468 => "00000000",
3469 => "00000000",
3470 => "00000000",
3471 => "00000000",
3472 => "00000000",
3473 => "00000000",
3474 => "00000000",
3475 => "00000000",
3476 => "00000000",
3477 => "00000000",
3478 => "00000000",
3479 => "00000000",
3480 => "00000000",
3481 => "00000000",
3482 => "00000000",
3483 => "00000000",
3484 => "00000000",
3485 => "00000000",
3486 => "00000000",
3487 => "00000000",
3488 => "00000000",
3489 => "00000000",
3490 => "00000000",
3491 => "00000000",
3492 => "00000000",
3493 => "00000000",
3494 => "00000000",
3495 => "00000000",
3496 => "00000000",
3497 => "00000000",
3498 => "00000000",
3499 => "00000000",
3500 => "00000000",
3501 => "00000000",
3502 => "00000000",
3503 => "00000000",
3504 => "00000000",
3505 => "00000000",
3506 => "00000000",
3507 => "00000000",
3508 => "00000000",
3509 => "00000000",
3510 => "00000000",
3511 => "00000000",
3512 => "00000000",
3513 => "00000000",
3514 => "00000000",
3515 => "00000000",
3516 => "00000000",
3517 => "00000000",
3518 => "00000000",
3519 => "00000000",
3520 => "00000000",
3521 => "00000000",
3522 => "00000000",
3523 => "00000000",
3524 => "00000000",
3525 => "00000000",
3526 => "00000000",
3527 => "00000000",
3528 => "00000000",
3529 => "00000000",
3530 => "00000000",
3531 => "00000000",
3532 => "00000000",
3533 => "00000000",
3534 => "00000000",
3535 => "00000000",
3536 => "00000000",
3537 => "00000000",
3538 => "00000000",
3539 => "00000000",
3540 => "00000000",
3541 => "00000000",
3542 => "00000000",
3543 => "00000000",
3544 => "00000000",
3545 => "00000000",
3546 => "00000000",
3547 => "00000000",
3548 => "00000000",
3549 => "00000000",
3550 => "00000000",
3551 => "00000000",
3552 => "00000000",
3553 => "00000000",
3554 => "00000000",
3555 => "00000000",
3556 => "00000000",
3557 => "00000000",
3558 => "00000000",
3559 => "00000000",
3560 => "00000000",
3561 => "00000000",
3562 => "00000000",
3563 => "00000000",
3564 => "00000000",
3565 => "00000000",
3566 => "00000000",
3567 => "00000000",
3568 => "00000000",
3569 => "00000000",
3570 => "00000000",
3571 => "00000000",
3572 => "00000000",
3584 => "00000000",
3585 => "00000000",
3586 => "00000000",
3587 => "00000000",
3588 => "00000000",
3589 => "00000000",
3590 => "00000000",
3591 => "00000000",
3592 => "00000000",
3593 => "00000000",
3594 => "00000000",
3595 => "00000000",
3596 => "00000000",
3597 => "00000000",
3598 => "00000000",
3599 => "00000000",
3600 => "00000000",
3601 => "00000000",
3602 => "00000000",
3603 => "00000000",
3604 => "00000000",
3605 => "00000000",
3606 => "00000000",
3607 => "00000000",
3608 => "00000000",
3609 => "00000000",
3610 => "00000000",
3611 => "00000000",
3612 => "00000000",
3613 => "00000000",
3614 => "00000000",
3615 => "00000000",
3616 => "00000000",
3617 => "00000000",
3618 => "00000000",
3619 => "00000000",
3620 => "00000000",
3621 => "00000000",
3622 => "00000000",
3623 => "00000000",
3624 => "00000000",
3625 => "00000000",
3626 => "00000000",
3627 => "00000000",
3628 => "00000000",
3629 => "00000000",
3630 => "00000000",
3631 => "00000000",
3632 => "00000000",
3633 => "00000000",
3634 => "00000000",
3635 => "00000000",
3636 => "00000000",
3637 => "00000000",
3638 => "00000000",
3639 => "00000000",
3640 => "00000000",
3641 => "00000000",
3642 => "00000000",
3643 => "00000000",
3644 => "00000000",
3645 => "00000000",
3646 => "00000000",
3647 => "00000000",
3648 => "00000000",
3649 => "00000000",
3650 => "00000000",
3651 => "00000000",
3652 => "00000000",
3653 => "00000000",
3654 => "00000000",
3655 => "00000000",
3656 => "00000000",
3657 => "00000000",
3658 => "00000000",
3659 => "00000000",
3660 => "00000000",
3661 => "00000000",
3662 => "00000000",
3663 => "00000000",
3664 => "00000000",
3665 => "00000000",
3666 => "00000000",
3667 => "00000000",
3668 => "00000000",
3669 => "00000000",
3670 => "00000000",
3671 => "00000000",
3672 => "00000000",
3673 => "00000000",
3674 => "00000000",
3675 => "00000000",
3676 => "00000000",
3677 => "00000000",
3678 => "00000000",
3679 => "00000000",
3680 => "00000000",
3681 => "00000000",
3682 => "00000000",
3683 => "00000000",
3684 => "00000000",
3685 => "00000000",
3686 => "00000000",
3687 => "00000000",
3688 => "00000000",
3689 => "00000000",
3690 => "00000000",
3691 => "00000000",
3692 => "00000000",
3693 => "00000000",
3694 => "00000000",
3695 => "00000000",
3696 => "00000000",
3697 => "00000000",
3698 => "00000000",
3699 => "00000000",
3700 => "00000000",
3712 => "00000000",
3713 => "00000000",
3714 => "00000000",
3715 => "00000000",
3716 => "00000000",
3717 => "00000000",
3718 => "00000000",
3719 => "00000000",
3720 => "00000000",
3721 => "00000000",
3722 => "00000000",
3723 => "00000000",
3724 => "00000000",
3725 => "00000000",
3726 => "00000000",
3727 => "00000000",
3728 => "00000000",
3729 => "00000000",
3730 => "00000000",
3731 => "00000000",
3732 => "00000000",
3733 => "00000000",
3734 => "00000000",
3735 => "00000000",
3736 => "00000000",
3737 => "00000000",
3738 => "00000000",
3739 => "00000000",
3740 => "00000000",
3741 => "00000000",
3742 => "00000000",
3743 => "00000000",
3744 => "00000000",
3745 => "00000000",
3746 => "00000000",
3747 => "00000000",
3748 => "00000000",
3749 => "00000000",
3750 => "00000000",
3751 => "00000000",
3752 => "00000000",
3753 => "00000000",
3754 => "00000000",
3755 => "00000000",
3756 => "00000000",
3757 => "00000000",
3758 => "00000000",
3759 => "00000000",
3760 => "00000000",
3761 => "00000000",
3762 => "00000000",
3763 => "00000000",
3764 => "00000000",
3765 => "00000000",
3766 => "00000000",
3767 => "00000000",
3768 => "00000000",
3769 => "00000000",
3770 => "00000000",
3771 => "00000000",
3772 => "00000000",
3773 => "00000000",
3774 => "00000000",
3775 => "00000000",
3776 => "00000000",
3777 => "00000000",
3778 => "00000000",
3779 => "00000000",
3780 => "00000000",
3781 => "00000000",
3782 => "00000000",
3783 => "00000000",
3784 => "00000000",
3785 => "00000000",
3786 => "00000000",
3787 => "00000000",
3788 => "00000000",
3789 => "00000000",
3790 => "00000000",
3791 => "00000000",
3792 => "00000000",
3793 => "00000000",
3794 => "00000000",
3795 => "00000000",
3796 => "00000000",
3797 => "00000000",
3798 => "00000000",
3799 => "00000000",
3800 => "00000000",
3801 => "00000000",
3802 => "00000000",
3803 => "00000000",
3804 => "00000000",
3805 => "00000000",
3806 => "00000000",
3807 => "00000000",
3808 => "00000000",
3809 => "00000000",
3810 => "00000000",
3811 => "00000000",
3812 => "00000000",
3813 => "00000000",
3814 => "00000000",
3815 => "00000000",
3816 => "00000000",
3817 => "00000000",
3818 => "00000000",
3819 => "00000000",
3820 => "00000000",
3821 => "00000000",
3822 => "00000000",
3823 => "00000000",
3824 => "00000000",
3825 => "00000000",
3826 => "00000000",
3827 => "00000000",
3828 => "00000000",
3840 => "00000000",
3841 => "00000000",
3842 => "00000000",
3843 => "00000000",
3844 => "00000000",
3845 => "00000000",
3846 => "00000000",
3847 => "00000000",
3848 => "00000000",
3849 => "00000000",
3850 => "00000000",
3851 => "00000000",
3852 => "00000000",
3853 => "00000000",
3854 => "00000000",
3855 => "00000000",
3856 => "00000000",
3857 => "00000000",
3858 => "00000000",
3859 => "00000000",
3860 => "00000000",
3861 => "00000000",
3862 => "00000000",
3863 => "00000000",
3864 => "00000000",
3865 => "00000000",
3866 => "00000000",
3867 => "00000000",
3868 => "00000000",
3869 => "00000000",
3870 => "00000000",
3871 => "00000000",
3872 => "00000000",
3873 => "00000000",
3874 => "00000000",
3875 => "00000000",
3876 => "00000000",
3877 => "00000000",
3878 => "00000000",
3879 => "00000000",
3880 => "00000000",
3881 => "00000000",
3882 => "00000000",
3883 => "00000000",
3884 => "00000000",
3885 => "00000000",
3886 => "00000000",
3887 => "00000000",
3888 => "00000000",
3889 => "00000000",
3890 => "00000000",
3891 => "00000000",
3892 => "00000000",
3893 => "00000000",
3894 => "00000000",
3895 => "00000000",
3896 => "00000000",
3897 => "00000000",
3898 => "00000000",
3899 => "00000000",
3900 => "00000000",
3901 => "00000000",
3902 => "00000000",
3903 => "00000000",
3904 => "00000000",
3905 => "00000000",
3906 => "00000000",
3907 => "00000000",
3908 => "00000000",
3909 => "00000000",
3910 => "00000000",
3911 => "00000000",
3912 => "00000000",
3913 => "00000000",
3914 => "00000000",
3915 => "00000000",
3916 => "00000000",
3917 => "00000000",
3918 => "00000000",
3919 => "00000000",
3920 => "00000000",
3921 => "00000000",
3922 => "00000000",
3923 => "00000000",
3924 => "00000000",
3925 => "00000000",
3926 => "00000000",
3927 => "00000000",
3928 => "00000000",
3929 => "00000000",
3930 => "00000000",
3931 => "00000000",
3932 => "00000000",
3933 => "00000000",
3934 => "00000000",
3935 => "00000000",
3936 => "00000000",
3937 => "00000000",
3938 => "00000000",
3939 => "00000000",
3940 => "00000000",
3941 => "00000000",
3942 => "00000000",
3943 => "00000000",
3944 => "00000000",
3945 => "00000000",
3946 => "00000000",
3947 => "00000000",
3948 => "00000000",
3949 => "00000000",
3950 => "00000000",
3951 => "00000000",
3952 => "00000000",
3953 => "00000000",
3954 => "00000000",
3955 => "00000000",
3956 => "00000000",
3968 => "00000000",
3969 => "00000000",
3970 => "00000000",
3971 => "00000000",
3972 => "00000000",
3973 => "00000000",
3974 => "00000000",
3975 => "00000000",
3976 => "00000000",
3977 => "00000000",
3978 => "00000000",
3979 => "00000000",
3980 => "00000000",
3981 => "00000000",
3982 => "00000000",
3983 => "00000000",
3984 => "00000000",
3985 => "00000000",
3986 => "00000000",
3987 => "00000000",
3988 => "00000000",
3989 => "00000000",
3990 => "00000000",
3991 => "00000000",
3992 => "00000000",
3993 => "00000000",
3994 => "00000000",
3995 => "00000000",
3996 => "00000000",
3997 => "00000000",
3998 => "00000000",
3999 => "00000000",
4000 => "00000000",
4001 => "00000000",
4002 => "00000000",
4003 => "00000000",
4004 => "00000000",
4005 => "00000000",
4006 => "00000000",
4007 => "00000000",
4008 => "00000000",
4009 => "00000000",
4010 => "00000000",
4011 => "00000000",
4012 => "00000000",
4013 => "00000000",
4014 => "00000000",
4015 => "00000000",
4016 => "00000000",
4017 => "00000000",
4018 => "00000000",
4019 => "00000000",
4020 => "00000000",
4021 => "00000000",
4022 => "00000000",
4023 => "00000000",
4024 => "00000000",
4025 => "00000000",
4026 => "00000000",
4027 => "00000000",
4028 => "00000000",
4029 => "00000000",
4030 => "00000000",
4031 => "00000000",
4032 => "00000000",
4033 => "00000000",
4034 => "00000000",
4035 => "00000000",
4036 => "00000000",
4037 => "00000000",
4038 => "00000000",
4039 => "00000000",
4040 => "00000000",
4041 => "00000000",
4042 => "00000000",
4043 => "00000000",
4044 => "00000000",
4045 => "00000000",
4046 => "00000000",
4047 => "00000000",
4048 => "00000000",
4049 => "00000000",
4050 => "00000000",
4051 => "00000000",
4052 => "00000000",
4053 => "00000000",
4054 => "00000000",
4055 => "00000000",
4056 => "00000000",
4057 => "00000000",
4058 => "00000000",
4059 => "00000000",
4060 => "00000000",
4061 => "00000000",
4062 => "00000000",
4063 => "00000000",
4064 => "00000000",
4065 => "00000000",
4066 => "00000000",
4067 => "00000000",
4068 => "00000000",
4069 => "00000000",
4070 => "00000000",
4071 => "00000000",
4072 => "00000000",
4073 => "00000000",
4074 => "00000000",
4075 => "00000000",
4076 => "00000000",
4077 => "00000000",
4078 => "00000000",
4079 => "00000000",
4080 => "00000000",
4081 => "00000000",
4082 => "00000000",
4083 => "00000000",
4084 => "00000000",
4096 => "00000000",
4097 => "00000000",
4098 => "00000000",
4099 => "00000000",
4100 => "00000000",
4101 => "00000000",
4102 => "00000000",
4103 => "00000000",
4104 => "00000000",
4105 => "00000000",
4106 => "00000000",
4107 => "00000000",
4108 => "00000000",
4109 => "00000000",
4110 => "00000000",
4111 => "00000000",
4112 => "00000000",
4113 => "00000000",
4114 => "00000000",
4115 => "00000000",
4116 => "00000000",
4117 => "00000000",
4118 => "00000000",
4119 => "00000000",
4120 => "00000000",
4121 => "00000000",
4122 => "00000000",
4123 => "00000000",
4124 => "00000000",
4125 => "00000000",
4126 => "00000000",
4127 => "00000000",
4128 => "00000000",
4129 => "00000000",
4130 => "00000000",
4131 => "00000000",
4132 => "00000000",
4133 => "00000000",
4134 => "00000000",
4135 => "00000000",
4136 => "00000000",
4137 => "00000000",
4138 => "00000000",
4139 => "00000000",
4140 => "00000000",
4141 => "00000000",
4142 => "00000000",
4143 => "00000000",
4144 => "00000000",
4145 => "00000000",
4146 => "00000000",
4147 => "00000000",
4148 => "00000000",
4149 => "00000000",
4150 => "00000000",
4151 => "00000000",
4152 => "00000000",
4153 => "00000000",
4154 => "00000000",
4155 => "00000000",
4156 => "00000000",
4157 => "00000000",
4158 => "00000000",
4159 => "00000000",
4160 => "00000000",
4161 => "00000000",
4162 => "00000000",
4163 => "00000000",
4164 => "00000000",
4165 => "00000000",
4166 => "00000000",
4167 => "00000000",
4168 => "00000000",
4169 => "00000000",
4170 => "00000000",
4171 => "00000000",
4172 => "00000000",
4173 => "00000000",
4174 => "00000000",
4175 => "00000000",
4176 => "00000000",
4177 => "00000000",
4178 => "00000000",
4179 => "00000000",
4180 => "00000000",
4181 => "00000000",
4182 => "00000000",
4183 => "00000000",
4184 => "00000000",
4185 => "00000000",
4186 => "00000000",
4187 => "00000000",
4188 => "00000000",
4189 => "00000000",
4190 => "00000000",
4191 => "00000000",
4192 => "00000000",
4193 => "00000000",
4194 => "00000000",
4195 => "00000000",
4196 => "00000000",
4197 => "00000000",
4198 => "00000000",
4199 => "00000000",
4200 => "00000000",
4201 => "00000000",
4202 => "00000000",
4203 => "00000000",
4204 => "00000000",
4205 => "00000000",
4206 => "00000000",
4207 => "00000000",
4208 => "00000000",
4209 => "00000000",
4210 => "00000000",
4211 => "00000000",
4212 => "00000000",
4224 => "00000000",
4225 => "00000000",
4226 => "00000000",
4227 => "00000000",
4228 => "00000000",
4229 => "00000000",
4230 => "00000000",
4231 => "00000000",
4232 => "00000000",
4233 => "00000000",
4234 => "00000000",
4235 => "00000000",
4236 => "00000000",
4237 => "00000000",
4238 => "00000000",
4239 => "00000000",
4240 => "00000000",
4241 => "00000000",
4242 => "00000000",
4243 => "00000000",
4244 => "00000000",
4245 => "00000000",
4246 => "00000000",
4247 => "00000000",
4248 => "00000000",
4249 => "00000000",
4250 => "00000000",
4251 => "00000000",
4252 => "00000000",
4253 => "00000000",
4254 => "00000000",
4255 => "00000000",
4256 => "00000000",
4257 => "00000000",
4258 => "00000000",
4259 => "00000000",
4260 => "00000000",
4261 => "00000000",
4262 => "00000000",
4263 => "00000000",
4264 => "00000000",
4265 => "00000000",
4266 => "00000000",
4267 => "00000000",
4268 => "00000000",
4269 => "00000000",
4270 => "00000000",
4271 => "00000000",
4272 => "00000000",
4273 => "00000000",
4274 => "00000000",
4275 => "00000000",
4276 => "00000000",
4277 => "00000000",
4278 => "00000000",
4279 => "00000000",
4280 => "00000000",
4281 => "00000000",
4282 => "00000000",
4283 => "00000000",
4284 => "00000000",
4285 => "00000000",
4286 => "00000000",
4287 => "00000000",
4288 => "00000000",
4289 => "00000000",
4290 => "00000000",
4291 => "00000000",
4292 => "00000000",
4293 => "00000000",
4294 => "00000000",
4295 => "00000000",
4296 => "00000000",
4297 => "00000000",
4298 => "00000000",
4299 => "00000000",
4300 => "00000000",
4301 => "00000000",
4302 => "00000000",
4303 => "00000000",
4304 => "00000000",
4305 => "00000000",
4306 => "00000000",
4307 => "00000000",
4308 => "00000000",
4309 => "00000000",
4310 => "00000000",
4311 => "00000000",
4312 => "00000000",
4313 => "00000000",
4314 => "00000000",
4315 => "00000000",
4316 => "00000000",
4317 => "00000000",
4318 => "00000000",
4319 => "00000000",
4320 => "00000000",
4321 => "00000000",
4322 => "00000000",
4323 => "00000000",
4324 => "00000000",
4325 => "00000000",
4326 => "00000000",
4327 => "00000000",
4328 => "00000000",
4329 => "00000000",
4330 => "00000000",
4331 => "00000000",
4332 => "00000000",
4333 => "00000000",
4334 => "00000000",
4335 => "00000000",
4336 => "00000000",
4337 => "00000000",
4338 => "00000000",
4339 => "00000000",
4340 => "00000000",
4352 => "00000000",
4353 => "00000000",
4354 => "00000000",
4355 => "00000000",
4356 => "00000000",
4357 => "00000000",
4358 => "00000000",
4359 => "00000000",
4360 => "00000000",
4361 => "00000000",
4362 => "00000000",
4363 => "00000000",
4364 => "00000000",
4365 => "00000000",
4366 => "00000000",
4367 => "00000000",
4368 => "00000000",
4369 => "00000000",
4370 => "00000000",
4371 => "01001001",
4372 => "00000000",
4373 => "01010010",
4374 => "01100011",
4375 => "00001001",
4376 => "00000000",
4377 => "00000000",
4378 => "00000000",
4379 => "00000000",
4380 => "00000000",
4381 => "00000000",
4382 => "00000000",
4383 => "00000000",
4384 => "00000000",
4385 => "00000000",
4386 => "00000000",
4387 => "00000000",
4388 => "00000000",
4389 => "00000000",
4390 => "00000000",
4391 => "00000000",
4392 => "00000000",
4393 => "00000000",
4394 => "00000000",
4395 => "00000000",
4396 => "00000000",
4397 => "00000000",
4398 => "00000000",
4399 => "00000000",
4400 => "00000000",
4401 => "00000000",
4402 => "00000000",
4403 => "00000000",
4404 => "00000000",
4405 => "00000000",
4406 => "00000000",
4407 => "00010001",
4408 => "01100010",
4409 => "00001000",
4410 => "00000000",
4411 => "00000000",
4412 => "00000000",
4413 => "00000000",
4414 => "00000000",
4415 => "00000000",
4416 => "00000000",
4417 => "00000000",
4418 => "00000000",
4419 => "00000000",
4420 => "00000000",
4421 => "00000000",
4422 => "00000000",
4423 => "00000000",
4424 => "00000000",
4425 => "00000000",
4426 => "00000000",
4427 => "00000000",
4428 => "00000000",
4429 => "00000000",
4430 => "00000000",
4431 => "00000000",
4432 => "00000000",
4433 => "00000000",
4434 => "00000000",
4435 => "00000000",
4436 => "00000000",
4437 => "00000000",
4438 => "00000000",
4439 => "00000000",
4440 => "00000000",
4441 => "00000000",
4442 => "00000000",
4443 => "00000000",
4444 => "00000000",
4445 => "00000000",
4446 => "00000000",
4447 => "00000000",
4448 => "00000000",
4449 => "00001001",
4450 => "01010010",
4451 => "01010010",
4452 => "01010010",
4453 => "01010010",
4454 => "01010010",
4455 => "01001001",
4456 => "00001001",
4457 => "00000000",
4458 => "00000000",
4459 => "00000000",
4460 => "00000000",
4461 => "00000000",
4462 => "00000000",
4463 => "00000000",
4464 => "00000000",
4465 => "00000000",
4466 => "00000000",
4467 => "00000000",
4468 => "00000000",
4480 => "00000000",
4481 => "00000000",
4482 => "00000000",
4483 => "00000000",
4484 => "00000000",
4485 => "00000000",
4486 => "00000000",
4487 => "00000000",
4488 => "00000000",
4489 => "00000000",
4490 => "00000000",
4491 => "00000000",
4492 => "00000000",
4493 => "00000000",
4494 => "01010010",
4495 => "00001000",
4496 => "01010010",
4497 => "10100100",
4498 => "01001001",
4499 => "11110110",
4500 => "01011011",
4501 => "10101101",
4502 => "11111111",
4503 => "01010010",
4504 => "00000000",
4505 => "00000000",
4506 => "00000000",
4507 => "00000000",
4508 => "00000000",
4509 => "00000000",
4510 => "00000000",
4511 => "00000000",
4512 => "00000000",
4513 => "00000000",
4514 => "00000000",
4515 => "00000000",
4516 => "00000000",
4517 => "00000000",
4518 => "00000000",
4519 => "00000000",
4520 => "00000000",
4521 => "00000000",
4522 => "00000000",
4523 => "00000000",
4524 => "00000000",
4525 => "00000000",
4526 => "00000000",
4527 => "00000000",
4528 => "00000000",
4529 => "00000000",
4530 => "00000000",
4531 => "00000000",
4532 => "00000000",
4533 => "00011001",
4534 => "01101010",
4535 => "01101011",
4536 => "01110011",
4537 => "01101010",
4538 => "00011001",
4539 => "00000000",
4540 => "00000000",
4541 => "00000000",
4542 => "00000000",
4543 => "00000000",
4544 => "00000000",
4545 => "00000000",
4546 => "00000000",
4547 => "00000000",
4548 => "00000000",
4549 => "00000000",
4550 => "00000000",
4551 => "00000000",
4552 => "00000000",
4553 => "00000000",
4554 => "00000000",
4555 => "00000000",
4556 => "00000000",
4557 => "00000000",
4558 => "00000000",
4559 => "00000000",
4560 => "00000000",
4561 => "00000000",
4562 => "00000000",
4563 => "00000000",
4564 => "00000000",
4565 => "00000000",
4566 => "00000000",
4567 => "00000000",
4568 => "00000000",
4569 => "00000000",
4570 => "00000000",
4571 => "00000000",
4572 => "00000000",
4573 => "00000000",
4574 => "01010010",
4575 => "10100100",
4576 => "10110110",
4577 => "11110110",
4578 => "11110110",
4579 => "10110110",
4580 => "10110110",
4581 => "10110110",
4582 => "11110110",
4583 => "11110110",
4584 => "11110110",
4585 => "10101101",
4586 => "10100100",
4587 => "01001001",
4588 => "00000000",
4589 => "00000000",
4590 => "00000000",
4591 => "00000000",
4592 => "00000000",
4593 => "00000000",
4594 => "00000000",
4595 => "00000000",
4596 => "00000000",
4608 => "00000000",
4609 => "00000000",
4610 => "00000000",
4611 => "00000000",
4612 => "00000000",
4613 => "00000000",
4614 => "00000000",
4615 => "00001001",
4616 => "00000000",
4617 => "01010010",
4618 => "00001001",
4619 => "01010010",
4620 => "10101101",
4621 => "01001001",
4622 => "11111111",
4623 => "10101101",
4624 => "10101101",
4625 => "11111111",
4626 => "11110110",
4627 => "11111111",
4628 => "11111111",
4629 => "11111111",
4630 => "11111111",
4631 => "01010010",
4632 => "00000000",
4633 => "00000000",
4634 => "00000000",
4635 => "00000000",
4636 => "00000000",
4637 => "00000000",
4638 => "00000000",
4639 => "00000000",
4640 => "00000000",
4641 => "00000000",
4642 => "00000000",
4643 => "00000000",
4644 => "00000000",
4645 => "00000000",
4646 => "00000000",
4647 => "00000000",
4648 => "00000000",
4649 => "00000000",
4650 => "00000000",
4651 => "00000000",
4652 => "00000000",
4653 => "00000000",
4654 => "00000000",
4655 => "00000000",
4656 => "00000000",
4657 => "00000000",
4658 => "00000000",
4659 => "00001000",
4660 => "00010001",
4661 => "01110011",
4662 => "01110011",
4663 => "01101011",
4664 => "01101011",
4665 => "01110011",
4666 => "01101011",
4667 => "00010001",
4668 => "00000000",
4669 => "00000000",
4670 => "00000000",
4671 => "00000000",
4672 => "00000000",
4673 => "00000000",
4674 => "00000000",
4675 => "00000000",
4676 => "00000000",
4677 => "00000000",
4678 => "00000000",
4679 => "00000000",
4680 => "00000000",
4681 => "00000000",
4682 => "00000000",
4683 => "00000000",
4684 => "00000000",
4685 => "00000000",
4686 => "00000000",
4687 => "00000000",
4688 => "00000000",
4689 => "00000000",
4690 => "00000000",
4691 => "00000000",
4692 => "00000000",
4693 => "00000000",
4694 => "00000000",
4695 => "00000000",
4696 => "00000000",
4697 => "00000000",
4698 => "00000000",
4699 => "00001000",
4700 => "01011011",
4701 => "11110110",
4702 => "11110110",
4703 => "10101101",
4704 => "01011011",
4705 => "01010001",
4706 => "01001001",
4707 => "01001001",
4708 => "00001000",
4709 => "01001000",
4710 => "01001001",
4711 => "01001001",
4712 => "01010010",
4713 => "10011011",
4714 => "10101101",
4715 => "11110110",
4716 => "10101101",
4717 => "01010010",
4718 => "00000000",
4719 => "00000000",
4720 => "00000000",
4721 => "00000000",
4722 => "00000000",
4723 => "00000000",
4724 => "00000000",
4736 => "00000000",
4737 => "00000000",
4738 => "01010010",
4739 => "00000000",
4740 => "01011011",
4741 => "01010010",
4742 => "01010010",
4743 => "11110110",
4744 => "01010010",
4745 => "11110110",
4746 => "10110110",
4747 => "10110110",
4748 => "11111111",
4749 => "11111111",
4750 => "11111111",
4751 => "11111111",
4752 => "11111111",
4753 => "11111111",
4754 => "11111111",
4755 => "11110110",
4756 => "11110110",
4757 => "11111111",
4758 => "11111111",
4759 => "11111111",
4760 => "01010010",
4761 => "00000000",
4762 => "00000000",
4763 => "00000000",
4764 => "00000000",
4765 => "00000000",
4766 => "00000000",
4767 => "00000000",
4768 => "00000000",
4769 => "00000000",
4770 => "00000000",
4771 => "00000000",
4772 => "00000000",
4773 => "00000000",
4774 => "00000000",
4775 => "00000000",
4776 => "00000000",
4777 => "00000000",
4778 => "00000000",
4779 => "00000000",
4780 => "00000000",
4781 => "00000000",
4782 => "00000000",
4783 => "00000000",
4784 => "00000000",
4785 => "00000000",
4786 => "00000000",
4787 => "00011001",
4788 => "01110011",
4789 => "01101011",
4790 => "01101011",
4791 => "01101011",
4792 => "01101011",
4793 => "01101011",
4794 => "01101011",
4795 => "01101010",
4796 => "00001000",
4797 => "00000000",
4798 => "00000000",
4799 => "00000000",
4800 => "00000000",
4801 => "00000000",
4802 => "00000000",
4803 => "00000000",
4804 => "00000000",
4805 => "00000000",
4806 => "00000000",
4807 => "00000000",
4808 => "00000000",
4809 => "00000000",
4810 => "00000000",
4811 => "00000000",
4812 => "00000000",
4813 => "00000000",
4814 => "00000000",
4815 => "00000000",
4816 => "00000000",
4817 => "00000000",
4818 => "00000000",
4819 => "00000000",
4820 => "00000000",
4821 => "00000000",
4822 => "00000000",
4823 => "00000000",
4824 => "00000000",
4825 => "00000000",
4826 => "01011011",
4827 => "11110110",
4828 => "10110110",
4829 => "01011011",
4830 => "01001001",
4831 => "01001000",
4832 => "01010001",
4833 => "10011011",
4834 => "10100011",
4835 => "10101100",
4836 => "10101100",
4837 => "10101100",
4838 => "10101100",
4839 => "10100011",
4840 => "10011010",
4841 => "01010001",
4842 => "01001000",
4843 => "01001001",
4844 => "10100100",
4845 => "11110110",
4846 => "10101101",
4847 => "01001001",
4848 => "00000000",
4849 => "00000000",
4850 => "00000000",
4851 => "00000000",
4852 => "00000000",
4864 => "01011011",
4865 => "01010010",
4866 => "11111111",
4867 => "01011011",
4868 => "11110110",
4869 => "11110110",
4870 => "10110110",
4871 => "11111111",
4872 => "11111111",
4873 => "11111111",
4874 => "11111111",
4875 => "11111111",
4876 => "11111111",
4877 => "11111110",
4878 => "11110110",
4879 => "11110101",
4880 => "11110101",
4881 => "11101101",
4882 => "11101100",
4883 => "11101100",
4884 => "11101101",
4885 => "11111111",
4886 => "11111111",
4887 => "10110110",
4888 => "00001001",
4889 => "00000000",
4890 => "00000000",
4891 => "00000000",
4892 => "00000000",
4893 => "00000000",
4894 => "00000000",
4895 => "00000000",
4896 => "00000000",
4897 => "00000000",
4898 => "00000000",
4899 => "00000000",
4900 => "00000000",
4901 => "00000000",
4902 => "00000000",
4903 => "00000000",
4904 => "00000000",
4905 => "00000000",
4906 => "00000000",
4907 => "00000000",
4908 => "00000000",
4909 => "00000000",
4910 => "00000000",
4911 => "00000000",
4912 => "00000000",
4913 => "00000000",
4914 => "00001000",
4915 => "01101010",
4916 => "01101011",
4917 => "01101011",
4918 => "01101011",
4919 => "01101011",
4920 => "01101011",
4921 => "01101011",
4922 => "01101011",
4923 => "01101011",
4924 => "01100010",
4925 => "00001000",
4926 => "00000000",
4927 => "00000000",
4928 => "00000000",
4929 => "00000000",
4930 => "00000000",
4931 => "00000000",
4932 => "00000000",
4933 => "00000000",
4934 => "00000000",
4935 => "00000000",
4936 => "00000000",
4937 => "00000000",
4938 => "00000000",
4939 => "00000000",
4940 => "00000000",
4941 => "00000000",
4942 => "00000000",
4943 => "00000000",
4944 => "00000000",
4945 => "00000000",
4946 => "00000000",
4947 => "00000000",
4948 => "00000000",
4949 => "00000000",
4950 => "00000000",
4951 => "00000000",
4952 => "00001001",
4953 => "10101101",
4954 => "11110110",
4955 => "01011011",
4956 => "00001000",
4957 => "01010001",
4958 => "10100011",
4959 => "11110101",
4960 => "11110101",
4961 => "11110101",
4962 => "11110101",
4963 => "11101100",
4964 => "11101100",
4965 => "11101100",
4966 => "11101101",
4967 => "11110101",
4968 => "11110101",
4969 => "11110101",
4970 => "11101100",
4971 => "10100011",
4972 => "01001001",
4973 => "01001001",
4974 => "10100100",
4975 => "11111111",
4976 => "01011011",
4977 => "00000000",
4978 => "00000000",
4979 => "00000000",
4980 => "00000000",
4992 => "11111111",
4993 => "11110110",
4994 => "11111111",
4995 => "11111111",
4996 => "11111111",
4997 => "11111111",
4998 => "11111111",
4999 => "11111110",
5000 => "11110110",
5001 => "11110110",
5002 => "11110101",
5003 => "11101101",
5004 => "11101100",
5005 => "11101100",
5006 => "11101100",
5007 => "11101100",
5008 => "11101100",
5009 => "11101100",
5010 => "11101100",
5011 => "11101100",
5012 => "11101100",
5013 => "11111111",
5014 => "11111111",
5015 => "10101101",
5016 => "00001000",
5017 => "00000000",
5018 => "00000000",
5019 => "00000000",
5020 => "00000000",
5021 => "00000000",
5022 => "00000000",
5023 => "00000000",
5024 => "00000000",
5025 => "00000000",
5026 => "00000000",
5027 => "00000000",
5028 => "00000000",
5029 => "00000000",
5030 => "00000000",
5031 => "00000000",
5032 => "00000000",
5033 => "00000000",
5034 => "00000000",
5035 => "00000000",
5036 => "00000000",
5037 => "00000000",
5038 => "00000000",
5039 => "00000000",
5040 => "00000000",
5041 => "00011001",
5042 => "01101010",
5043 => "01101011",
5044 => "01101011",
5045 => "01101011",
5046 => "01101011",
5047 => "01101011",
5048 => "01101011",
5049 => "01101011",
5050 => "01101011",
5051 => "01101011",
5052 => "01110011",
5053 => "01100010",
5054 => "00001000",
5055 => "00000000",
5056 => "00000000",
5057 => "00000000",
5058 => "00000000",
5059 => "00000000",
5060 => "00000000",
5061 => "00000000",
5062 => "00000000",
5063 => "00000000",
5064 => "00000000",
5065 => "00000000",
5066 => "00000000",
5067 => "00000000",
5068 => "00000000",
5069 => "00000000",
5070 => "00000000",
5071 => "00000000",
5072 => "00000000",
5073 => "00000000",
5074 => "00000000",
5075 => "00000000",
5076 => "00000000",
5077 => "00000000",
5078 => "00000000",
5079 => "01001001",
5080 => "11110110",
5081 => "10101101",
5082 => "01001001",
5083 => "01001001",
5084 => "10100011",
5085 => "11110101",
5086 => "11101100",
5087 => "10101100",
5088 => "10101100",
5089 => "10101100",
5090 => "10101100",
5091 => "10101100",
5092 => "10101100",
5093 => "10101100",
5094 => "10101100",
5095 => "10101100",
5096 => "10101100",
5097 => "10101100",
5098 => "10101100",
5099 => "11110101",
5100 => "11110101",
5101 => "10100011",
5102 => "00001000",
5103 => "01010010",
5104 => "11110110",
5105 => "10100100",
5106 => "00000000",
5107 => "00000000",
5108 => "00000000",
5120 => "11111111",
5121 => "11111111",
5122 => "11110110",
5123 => "11110110",
5124 => "11110101",
5125 => "11110101",
5126 => "11101100",
5127 => "11101100",
5128 => "11101100",
5129 => "11101100",
5130 => "11101100",
5131 => "11101100",
5132 => "11101100",
5133 => "11101100",
5134 => "11101100",
5135 => "11101100",
5136 => "11101100",
5137 => "11101100",
5138 => "11101100",
5139 => "11101100",
5140 => "11101100",
5141 => "11111110",
5142 => "11111111",
5143 => "11111111",
5144 => "10101101",
5145 => "00000000",
5146 => "00000000",
5147 => "00000000",
5148 => "00000000",
5149 => "00000000",
5150 => "00000000",
5151 => "00000000",
5152 => "00000000",
5153 => "00000000",
5154 => "00000000",
5155 => "00000000",
5156 => "00000000",
5157 => "00000000",
5158 => "00000000",
5159 => "00000000",
5160 => "00000000",
5161 => "00000000",
5162 => "00000000",
5163 => "00000000",
5164 => "00000000",
5165 => "00000000",
5166 => "00000000",
5167 => "00000000",
5168 => "01011001",
5169 => "01110011",
5170 => "01101011",
5171 => "01101011",
5172 => "01101011",
5173 => "01101010",
5174 => "01101010",
5175 => "01101011",
5176 => "01101011",
5177 => "01101010",
5178 => "01101010",
5179 => "01101011",
5180 => "01101011",
5181 => "01110011",
5182 => "01100010",
5183 => "00001000",
5184 => "00000000",
5185 => "00000000",
5186 => "00000000",
5187 => "00000000",
5188 => "00000000",
5189 => "00000000",
5190 => "00000000",
5191 => "00000000",
5192 => "00000000",
5193 => "00000000",
5194 => "00000000",
5195 => "00000000",
5196 => "00000000",
5197 => "00000000",
5198 => "00000000",
5199 => "00000000",
5200 => "00000000",
5201 => "00000000",
5202 => "00000000",
5203 => "00000000",
5204 => "00000000",
5205 => "00000000",
5206 => "01001001",
5207 => "11110110",
5208 => "10100100",
5209 => "00000000",
5210 => "01010001",
5211 => "11101100",
5212 => "11101100",
5213 => "10101100",
5214 => "10101011",
5215 => "10101100",
5216 => "10101100",
5217 => "10101100",
5218 => "10101100",
5219 => "10101100",
5220 => "11101100",
5221 => "10101100",
5222 => "10101100",
5223 => "10101100",
5224 => "10101100",
5225 => "10101100",
5226 => "10101100",
5227 => "10101100",
5228 => "10101100",
5229 => "11110101",
5230 => "10101100",
5231 => "01001000",
5232 => "01001001",
5233 => "11110110",
5234 => "10101101",
5235 => "00000000",
5236 => "00000000",
5248 => "11101101",
5249 => "11101100",
5250 => "11101100",
5251 => "11101100",
5252 => "11101100",
5253 => "10100011",
5254 => "10101100",
5255 => "11101100",
5256 => "11101101",
5257 => "11101100",
5258 => "11101100",
5259 => "11101100",
5260 => "11101100",
5261 => "11101100",
5262 => "11101100",
5263 => "11101100",
5264 => "11101100",
5265 => "11101100",
5266 => "11101100",
5267 => "11101100",
5268 => "11101100",
5269 => "11110110",
5270 => "11111111",
5271 => "11111111",
5272 => "01010010",
5273 => "00000000",
5274 => "00000000",
5275 => "00000000",
5276 => "00000000",
5277 => "00000000",
5278 => "00000000",
5279 => "00000000",
5280 => "00000000",
5281 => "00000000",
5282 => "00000000",
5283 => "00000000",
5284 => "00000000",
5285 => "00000000",
5286 => "00000000",
5287 => "00000000",
5288 => "00000000",
5289 => "00000000",
5290 => "00000000",
5291 => "00000000",
5292 => "00000000",
5293 => "00010001",
5294 => "00010001",
5295 => "01100001",
5296 => "01110011",
5297 => "01101010",
5298 => "01100010",
5299 => "01101010",
5300 => "01101010",
5301 => "01101010",
5302 => "01101010",
5303 => "01101010",
5304 => "01101010",
5305 => "01101010",
5306 => "01101010",
5307 => "01101010",
5308 => "01101010",
5309 => "01101010",
5310 => "01101011",
5311 => "01100010",
5312 => "00010001",
5313 => "01011001",
5314 => "00001000",
5315 => "00000000",
5316 => "00000000",
5317 => "00000000",
5318 => "00000000",
5319 => "00000000",
5320 => "00000000",
5321 => "00000000",
5322 => "00000000",
5323 => "00000000",
5324 => "00000000",
5325 => "00000000",
5326 => "00000000",
5327 => "00000000",
5328 => "00000000",
5329 => "00000000",
5330 => "00000000",
5331 => "00000000",
5332 => "00000000",
5333 => "00001001",
5334 => "11110110",
5335 => "10100100",
5336 => "00000000",
5337 => "10011010",
5338 => "11101100",
5339 => "10101011",
5340 => "10100011",
5341 => "10101011",
5342 => "10101011",
5343 => "10101011",
5344 => "10101011",
5345 => "11101011",
5346 => "11101011",
5347 => "11101011",
5348 => "11101011",
5349 => "11101100",
5350 => "11101100",
5351 => "11101100",
5352 => "11101100",
5353 => "11101011",
5354 => "11101011",
5355 => "10101011",
5356 => "10101011",
5357 => "10100011",
5358 => "10101100",
5359 => "11101100",
5360 => "01010000",
5361 => "01001001",
5362 => "10110110",
5363 => "10100100",
5364 => "00000000",
5376 => "11101100",
5377 => "11101100",
5378 => "11101100",
5379 => "10100100",
5380 => "10100011",
5381 => "10100100",
5382 => "10011011",
5383 => "10100100",
5384 => "11101100",
5385 => "11101100",
5386 => "11101100",
5387 => "11101100",
5388 => "11101100",
5389 => "11101100",
5390 => "11101100",
5391 => "11101100",
5392 => "11101100",
5393 => "11101100",
5394 => "11101100",
5395 => "11101100",
5396 => "11101100",
5397 => "11110101",
5398 => "11111111",
5399 => "11111111",
5400 => "01011011",
5401 => "00000000",
5402 => "00000000",
5403 => "00000000",
5404 => "00000000",
5405 => "00000000",
5406 => "00000000",
5407 => "00000000",
5408 => "00000000",
5409 => "00000000",
5410 => "00000000",
5411 => "00000000",
5412 => "00000000",
5413 => "00000000",
5414 => "00000000",
5415 => "00000000",
5416 => "00000000",
5417 => "00000000",
5418 => "00000000",
5419 => "00000000",
5420 => "00000000",
5421 => "00011001",
5422 => "01110011",
5423 => "01101010",
5424 => "01101010",
5425 => "01100010",
5426 => "01101010",
5427 => "01101010",
5428 => "01101010",
5429 => "01101010",
5430 => "01101010",
5431 => "01101010",
5432 => "01101010",
5433 => "01101010",
5434 => "01101010",
5435 => "01101010",
5436 => "01101010",
5437 => "01100010",
5438 => "01100010",
5439 => "01101010",
5440 => "01110010",
5441 => "01110010",
5442 => "00010001",
5443 => "00000000",
5444 => "00000000",
5445 => "00000000",
5446 => "00000000",
5447 => "00000000",
5448 => "00000000",
5449 => "00000000",
5450 => "00000000",
5451 => "00000000",
5452 => "00000000",
5453 => "00000000",
5454 => "00000000",
5455 => "00000000",
5456 => "00000000",
5457 => "00000000",
5458 => "00000000",
5459 => "00000000",
5460 => "00000000",
5461 => "10101101",
5462 => "10101101",
5463 => "00000000",
5464 => "01010001",
5465 => "10101100",
5466 => "10100011",
5467 => "10100011",
5468 => "10101011",
5469 => "10101011",
5470 => "10101011",
5471 => "10101011",
5472 => "10101011",
5473 => "11101011",
5474 => "11101011",
5475 => "11101011",
5476 => "11101011",
5477 => "11101010",
5478 => "10100010",
5479 => "10100010",
5480 => "10100010",
5481 => "10100010",
5482 => "10100010",
5483 => "10100010",
5484 => "10100010",
5485 => "10100011",
5486 => "10100011",
5487 => "10101011",
5488 => "10101011",
5489 => "01001000",
5490 => "01001001",
5491 => "11110110",
5492 => "01011011",
5504 => "11101100",
5505 => "11101100",
5506 => "11101100",
5507 => "10100100",
5508 => "10100100",
5509 => "10100100",
5510 => "10101100",
5511 => "10101100",
5512 => "10100100",
5513 => "11101100",
5514 => "11101100",
5515 => "11101100",
5516 => "11101100",
5517 => "11101100",
5518 => "11101100",
5519 => "11101100",
5520 => "11101100",
5521 => "11101100",
5522 => "11101100",
5523 => "11101100",
5524 => "11101100",
5525 => "11110101",
5526 => "11111111",
5527 => "11111111",
5528 => "11111111",
5529 => "01010010",
5530 => "00000000",
5531 => "00000000",
5532 => "00000000",
5533 => "00000000",
5534 => "00000000",
5535 => "00000000",
5536 => "00000000",
5537 => "00000000",
5538 => "00000000",
5539 => "00000000",
5540 => "00000000",
5541 => "00000000",
5542 => "00000000",
5543 => "00000000",
5544 => "00000000",
5545 => "00000000",
5546 => "00000000",
5547 => "00000000",
5548 => "00001000",
5549 => "00011001",
5550 => "01101010",
5551 => "01100010",
5552 => "01100010",
5553 => "01100010",
5554 => "01101010",
5555 => "01101010",
5556 => "01101010",
5557 => "01101010",
5558 => "01101010",
5559 => "01101010",
5560 => "01101010",
5561 => "01101010",
5562 => "01101010",
5563 => "01101010",
5564 => "01101010",
5565 => "01100010",
5566 => "01100010",
5567 => "01100010",
5568 => "01100010",
5569 => "01101010",
5570 => "00010001",
5571 => "00000000",
5572 => "00000000",
5573 => "00000000",
5574 => "00000000",
5575 => "00000000",
5576 => "00000000",
5577 => "00000000",
5578 => "00000000",
5579 => "00000000",
5580 => "00000000",
5581 => "00000000",
5582 => "00000000",
5583 => "00000000",
5584 => "00000000",
5585 => "00000000",
5586 => "00000000",
5587 => "00000000",
5588 => "10100100",
5589 => "11110110",
5590 => "01001001",
5591 => "01010000",
5592 => "10100011",
5593 => "10100011",
5594 => "10100011",
5595 => "10100011",
5596 => "10100011",
5597 => "10101011",
5598 => "10101011",
5599 => "11101011",
5600 => "11101011",
5601 => "10101010",
5602 => "10100010",
5603 => "10100010",
5604 => "10100010",
5605 => "10100011",
5606 => "10101011",
5607 => "10101100",
5608 => "10101101",
5609 => "10110101",
5610 => "11110110",
5611 => "11110110",
5612 => "11110110",
5613 => "10100010",
5614 => "10100011",
5615 => "10100011",
5616 => "10100011",
5617 => "10100010",
5618 => "01001000",
5619 => "01010010",
5620 => "11111110",
5632 => "11101100",
5633 => "11101100",
5634 => "11101100",
5635 => "11101100",
5636 => "10101100",
5637 => "10101101",
5638 => "10101101",
5639 => "10101101",
5640 => "10101101",
5641 => "11101100",
5642 => "11101100",
5643 => "11101100",
5644 => "11101100",
5645 => "11101100",
5646 => "11101100",
5647 => "11101100",
5648 => "11101100",
5649 => "11101100",
5650 => "11101100",
5651 => "11101100",
5652 => "11101100",
5653 => "11101100",
5654 => "11111111",
5655 => "11111111",
5656 => "10101101",
5657 => "00000000",
5658 => "00000000",
5659 => "00000000",
5660 => "00000000",
5661 => "00000000",
5662 => "00000000",
5663 => "00000000",
5664 => "00000000",
5665 => "00000000",
5666 => "00000000",
5667 => "00000000",
5668 => "00000000",
5669 => "00000000",
5670 => "00000000",
5671 => "00000000",
5672 => "00000000",
5673 => "00000000",
5674 => "00000000",
5675 => "00000000",
5676 => "00000000",
5677 => "00010001",
5678 => "01101010",
5679 => "01100010",
5680 => "01100010",
5681 => "01100010",
5682 => "01101010",
5683 => "01101010",
5684 => "01101010",
5685 => "01101010",
5686 => "01101010",
5687 => "01101010",
5688 => "01101010",
5689 => "01101010",
5690 => "01101010",
5691 => "01101010",
5692 => "01101010",
5693 => "01101010",
5694 => "01100010",
5695 => "01100010",
5696 => "01100010",
5697 => "01101010",
5698 => "01100010",
5699 => "00001000",
5700 => "00000000",
5701 => "00000000",
5702 => "00000000",
5703 => "00000000",
5704 => "00000000",
5705 => "00000000",
5706 => "00000000",
5707 => "00000000",
5708 => "00000000",
5709 => "00000000",
5710 => "00000000",
5711 => "00000000",
5712 => "00000000",
5713 => "00000000",
5714 => "00000000",
5715 => "01001001",
5716 => "11110110",
5717 => "01010010",
5718 => "01001000",
5719 => "10011001",
5720 => "10100011",
5721 => "10100010",
5722 => "10100011",
5723 => "10100011",
5724 => "10100011",
5725 => "10101011",
5726 => "10101011",
5727 => "10100010",
5728 => "10100001",
5729 => "10100010",
5730 => "10101100",
5731 => "10101101",
5732 => "11110110",
5733 => "11111111",
5734 => "11111111",
5735 => "11111111",
5736 => "11111111",
5737 => "11111111",
5738 => "11111111",
5739 => "11111111",
5740 => "11110110",
5741 => "10011010",
5742 => "10100010",
5743 => "10100011",
5744 => "10100011",
5745 => "10100011",
5746 => "10010000",
5747 => "01001000",
5748 => "10100100",
5760 => "11101100",
5761 => "11101100",
5762 => "11101100",
5763 => "10011011",
5764 => "10100100",
5765 => "10101101",
5766 => "10101101",
5767 => "10101101",
5768 => "10100100",
5769 => "10100011",
5770 => "11101100",
5771 => "11101100",
5772 => "11101100",
5773 => "11101100",
5774 => "11101100",
5775 => "11101100",
5776 => "11101100",
5777 => "11101100",
5778 => "11101100",
5779 => "11101100",
5780 => "11101100",
5781 => "11101100",
5782 => "11111110",
5783 => "11111111",
5784 => "10101101",
5785 => "01001001",
5786 => "00000000",
5787 => "00000000",
5788 => "00000000",
5789 => "00000000",
5790 => "00000000",
5791 => "00000000",
5792 => "00000000",
5793 => "00000000",
5794 => "00000000",
5795 => "00000000",
5796 => "00000000",
5797 => "00000000",
5798 => "00000000",
5799 => "00000000",
5800 => "00000000",
5801 => "00000000",
5802 => "00000000",
5803 => "00000000",
5804 => "00011001",
5805 => "00011001",
5806 => "01101010",
5807 => "01100010",
5808 => "01100010",
5809 => "01100010",
5810 => "01101010",
5811 => "01101010",
5812 => "01101010",
5813 => "01101010",
5814 => "01101010",
5815 => "01101010",
5816 => "01101010",
5817 => "01101010",
5818 => "01101010",
5819 => "01101010",
5820 => "01101010",
5821 => "01101010",
5822 => "01100010",
5823 => "01100010",
5824 => "01100010",
5825 => "01101010",
5826 => "00011001",
5827 => "00000000",
5828 => "00000000",
5829 => "00000000",
5830 => "00000000",
5831 => "00000000",
5832 => "00000000",
5833 => "00000000",
5834 => "00000000",
5835 => "00000000",
5836 => "00000000",
5837 => "00000000",
5838 => "00000000",
5839 => "00000000",
5840 => "00000000",
5841 => "00000000",
5842 => "00000000",
5843 => "10101101",
5844 => "10101101",
5845 => "01001000",
5846 => "01010000",
5847 => "10100010",
5848 => "10100010",
5849 => "10100010",
5850 => "10100010",
5851 => "10100010",
5852 => "10100010",
5853 => "10101010",
5854 => "10100010",
5855 => "10100010",
5856 => "10110110",
5857 => "11110111",
5858 => "11111111",
5859 => "11111111",
5860 => "11111111",
5861 => "11110110",
5862 => "11110110",
5863 => "11110110",
5864 => "11111111",
5865 => "11111110",
5866 => "11111111",
5867 => "11111111",
5868 => "11110110",
5869 => "10011010",
5870 => "10100010",
5871 => "10100010",
5872 => "10100010",
5873 => "10100010",
5874 => "10011001",
5875 => "01001000",
5876 => "01001001",
5888 => "11101100",
5889 => "11101100",
5890 => "11101100",
5891 => "10100100",
5892 => "10100100",
5893 => "10101100",
5894 => "10101101",
5895 => "10100100",
5896 => "10100100",
5897 => "01011011",
5898 => "11101100",
5899 => "11101100",
5900 => "11101100",
5901 => "11101100",
5902 => "11101100",
5903 => "11101100",
5904 => "11101100",
5905 => "11101100",
5906 => "11101100",
5907 => "11101100",
5908 => "11101100",
5909 => "11101100",
5910 => "11110110",
5911 => "11111111",
5912 => "11111111",
5913 => "10101101",
5914 => "00000000",
5915 => "00000000",
5916 => "00000000",
5917 => "00000000",
5918 => "00000000",
5919 => "00000000",
5920 => "00000000",
5921 => "00000000",
5922 => "00000000",
5923 => "00000000",
5924 => "00000000",
5925 => "00000000",
5926 => "00000000",
5927 => "00000000",
5928 => "00000000",
5929 => "00000000",
5930 => "00000000",
5931 => "00000000",
5932 => "00011001",
5933 => "01110010",
5934 => "01100010",
5935 => "01100010",
5936 => "01100010",
5937 => "01100010",
5938 => "01101010",
5939 => "01101010",
5940 => "01100010",
5941 => "01100010",
5942 => "01101010",
5943 => "01101010",
5944 => "01101010",
5945 => "01100010",
5946 => "01100010",
5947 => "01101010",
5948 => "01101010",
5949 => "01100010",
5950 => "01100010",
5951 => "01100010",
5952 => "01100010",
5953 => "01100010",
5954 => "01100001",
5955 => "00011001",
5956 => "00000000",
5957 => "00000000",
5958 => "00000000",
5959 => "00000000",
5960 => "00000000",
5961 => "00000000",
5962 => "00000000",
5963 => "00000000",
5964 => "00000000",
5965 => "00000000",
5966 => "00000000",
5967 => "00000000",
5968 => "00000000",
5969 => "00000000",
5970 => "01010001",
5971 => "11110110",
5972 => "01010010",
5973 => "01001000",
5974 => "10010000",
5975 => "10100010",
5976 => "10100010",
5977 => "10100010",
5978 => "10100010",
5979 => "10100010",
5980 => "10100010",
5981 => "10101010",
5982 => "10100001",
5983 => "10100011",
5984 => "11111111",
5985 => "11110110",
5986 => "11110110",
5987 => "11110110",
5988 => "11110110",
5989 => "11110110",
5990 => "11110110",
5991 => "11110110",
5992 => "11110110",
5993 => "11111110",
5994 => "11110110",
5995 => "11111111",
5996 => "11110110",
5997 => "10011010",
5998 => "10100010",
5999 => "10100010",
6000 => "10100010",
6001 => "10100010",
6002 => "10011010",
6003 => "10010000",
6004 => "01001000",
6016 => "11101100",
6017 => "11101100",
6018 => "11101100",
6019 => "11101100",
6020 => "10100100",
6021 => "10100100",
6022 => "10100100",
6023 => "10100100",
6024 => "10101101",
6025 => "10101101",
6026 => "10100100",
6027 => "11101100",
6028 => "11101100",
6029 => "11101100",
6030 => "11101100",
6031 => "11101100",
6032 => "11101100",
6033 => "11101100",
6034 => "11101100",
6035 => "11101100",
6036 => "11101100",
6037 => "11101100",
6038 => "11110110",
6039 => "11111111",
6040 => "11111111",
6041 => "01010010",
6042 => "00000000",
6043 => "00000000",
6044 => "00000000",
6045 => "00000000",
6046 => "00000000",
6047 => "00000000",
6048 => "00000000",
6049 => "00000000",
6050 => "00000000",
6051 => "00000000",
6052 => "00000000",
6053 => "00000000",
6054 => "00000000",
6055 => "00000000",
6056 => "00000000",
6057 => "00000000",
6058 => "00000000",
6059 => "00000000",
6060 => "00000000",
6061 => "01100010",
6062 => "01100010",
6063 => "01100010",
6064 => "01100010",
6065 => "01100010",
6066 => "01101010",
6067 => "01101010",
6068 => "01100010",
6069 => "01100010",
6070 => "01100010",
6071 => "01100010",
6072 => "01101010",
6073 => "01100010",
6074 => "01100010",
6075 => "01100010",
6076 => "01101010",
6077 => "01100010",
6078 => "01100010",
6079 => "01100010",
6080 => "01100010",
6081 => "01100010",
6082 => "01011001",
6083 => "00001000",
6084 => "00000000",
6085 => "00000000",
6086 => "00000000",
6087 => "00000000",
6088 => "00000000",
6089 => "00000000",
6090 => "00000000",
6091 => "00000000",
6092 => "00000000",
6093 => "00000000",
6094 => "00000000",
6095 => "00000000",
6096 => "00000000",
6097 => "00000000",
6098 => "10100100",
6099 => "10101101",
6100 => "01001000",
6101 => "01010000",
6102 => "10011000",
6103 => "10100010",
6104 => "10100010",
6105 => "10100010",
6106 => "10100010",
6107 => "10100010",
6108 => "10100010",
6109 => "11101010",
6110 => "10100000",
6111 => "10100011",
6112 => "11111111",
6113 => "11110110",
6114 => "11110110",
6115 => "11110110",
6116 => "11110110",
6117 => "11110110",
6118 => "11110110",
6119 => "11110110",
6120 => "11110110",
6121 => "11110110",
6122 => "11110110",
6123 => "11111111",
6124 => "11110110",
6125 => "10011010",
6126 => "10100001",
6127 => "10100010",
6128 => "10100010",
6129 => "10100010",
6130 => "10011010",
6131 => "10010000",
6132 => "01001000",
6144 => "11101100",
6145 => "11101100",
6146 => "11101100",
6147 => "11101100",
6148 => "01011011",
6149 => "10100100",
6150 => "10100100",
6151 => "10100100",
6152 => "01100100",
6153 => "10100101",
6154 => "10101101",
6155 => "11101100",
6156 => "11101100",
6157 => "11101100",
6158 => "11101100",
6159 => "11101100",
6160 => "11101100",
6161 => "11101100",
6162 => "11101100",
6163 => "11101100",
6164 => "11101100",
6165 => "11101100",
6166 => "11110101",
6167 => "11111111",
6168 => "11111111",
6169 => "01011011",
6170 => "00001001",
6171 => "00000000",
6172 => "00000000",
6173 => "00000000",
6174 => "00000000",
6175 => "00000000",
6176 => "00000000",
6177 => "00000000",
6178 => "00000000",
6179 => "00000000",
6180 => "00000000",
6181 => "00000000",
6182 => "00000000",
6183 => "00000000",
6184 => "00000000",
6185 => "00000000",
6186 => "00000000",
6187 => "00000000",
6188 => "00000000",
6189 => "00010001",
6190 => "01100010",
6191 => "01100010",
6192 => "01100010",
6193 => "01100010",
6194 => "01100010",
6195 => "01101010",
6196 => "01100010",
6197 => "01100010",
6198 => "01101010",
6199 => "01100010",
6200 => "01101010",
6201 => "01100010",
6202 => "01100010",
6203 => "01101010",
6204 => "01100010",
6205 => "01100010",
6206 => "01100010",
6207 => "01100010",
6208 => "01100010",
6209 => "01101010",
6210 => "00001000",
6211 => "00000000",
6212 => "00000000",
6213 => "00000000",
6214 => "00000000",
6215 => "00000000",
6216 => "00000000",
6217 => "00000000",
6218 => "00000000",
6219 => "00000000",
6220 => "00000000",
6221 => "00000000",
6222 => "00000000",
6223 => "00000000",
6224 => "00000000",
6225 => "00000000",
6226 => "10110110",
6227 => "01011011",
6228 => "01001000",
6229 => "10010000",
6230 => "10011000",
6231 => "10100001",
6232 => "10100001",
6233 => "10100001",
6234 => "10100001",
6235 => "10100001",
6236 => "10100001",
6237 => "11101001",
6238 => "10100000",
6239 => "10100011",
6240 => "11110111",
6241 => "11110110",
6242 => "11110110",
6243 => "11110110",
6244 => "11110110",
6245 => "11110110",
6246 => "11111111",
6247 => "11111111",
6248 => "11111111",
6249 => "11110111",
6250 => "11110110",
6251 => "11111111",
6252 => "11110110",
6253 => "10011001",
6254 => "10100001",
6255 => "10100001",
6256 => "10100001",
6257 => "10100001",
6258 => "10011001",
6259 => "10010000",
6260 => "10010000",
6272 => "11101100",
6273 => "11101100",
6274 => "11101100",
6275 => "11101100",
6276 => "01011011",
6277 => "10100100",
6278 => "10100100",
6279 => "10100100",
6280 => "10100100",
6281 => "01100100",
6282 => "01011011",
6283 => "11101100",
6284 => "11101100",
6285 => "11101100",
6286 => "11101100",
6287 => "11101100",
6288 => "11101100",
6289 => "11101100",
6290 => "11101100",
6291 => "11101100",
6292 => "11101100",
6293 => "11101100",
6294 => "11101100",
6295 => "11111111",
6296 => "11111111",
6297 => "11111111",
6298 => "01010010",
6299 => "00000000",
6300 => "00000000",
6301 => "00000000",
6302 => "00000000",
6303 => "00000000",
6304 => "00000000",
6305 => "00000000",
6306 => "00000000",
6307 => "00000000",
6308 => "00000000",
6309 => "00000000",
6310 => "00000000",
6311 => "00000000",
6312 => "00000000",
6313 => "00000000",
6314 => "00000000",
6315 => "00000000",
6316 => "00000000",
6317 => "00010001",
6318 => "01101010",
6319 => "01100010",
6320 => "01100010",
6321 => "01100010",
6322 => "01100010",
6323 => "01100010",
6324 => "01101010",
6325 => "01101010",
6326 => "01100010",
6327 => "01100010",
6328 => "01100010",
6329 => "01101010",
6330 => "01101010",
6331 => "01101010",
6332 => "01100010",
6333 => "01100010",
6334 => "01100010",
6335 => "01100010",
6336 => "01100010",
6337 => "01100010",
6338 => "01101010",
6339 => "00011001",
6340 => "00000000",
6341 => "00000000",
6342 => "00000000",
6343 => "00000000",
6344 => "00000000",
6345 => "00000000",
6346 => "00000000",
6347 => "00000000",
6348 => "00000000",
6349 => "00000000",
6350 => "00000000",
6351 => "00000000",
6352 => "00000000",
6353 => "01010010",
6354 => "11110110",
6355 => "01010001",
6356 => "01010000",
6357 => "10010000",
6358 => "10011000",
6359 => "10011001",
6360 => "10100001",
6361 => "10100001",
6362 => "10100001",
6363 => "10100000",
6364 => "10100000",
6365 => "11101001",
6366 => "10100000",
6367 => "10100011",
6368 => "11110111",
6369 => "11110110",
6370 => "11110111",
6371 => "11110110",
6372 => "10110110",
6373 => "10101101",
6374 => "10101100",
6375 => "10100011",
6376 => "10100011",
6377 => "10011010",
6378 => "10011010",
6379 => "11110110",
6380 => "11110110",
6381 => "10011001",
6382 => "10100000",
6383 => "10100001",
6384 => "10100001",
6385 => "10100001",
6386 => "10011001",
6387 => "10010000",
6388 => "10010000",
6400 => "11101100",
6401 => "11101100",
6402 => "11101100",
6403 => "11101100",
6404 => "10100011",
6405 => "01011011",
6406 => "10100100",
6407 => "10100011",
6408 => "10100100",
6409 => "01011100",
6410 => "00000001",
6411 => "10100011",
6412 => "11101100",
6413 => "11101100",
6414 => "11101100",
6415 => "11101100",
6416 => "11101100",
6417 => "11101100",
6418 => "11101100",
6419 => "11101100",
6420 => "11101100",
6421 => "11101100",
6422 => "11101100",
6423 => "11111111",
6424 => "11111111",
6425 => "10101101",
6426 => "00000000",
6427 => "00000000",
6428 => "00000000",
6429 => "00000000",
6430 => "00000000",
6431 => "00000000",
6432 => "00000000",
6433 => "00000000",
6434 => "00000000",
6435 => "00000000",
6436 => "00000000",
6437 => "00000000",
6438 => "00000000",
6439 => "00000000",
6440 => "00000000",
6441 => "00000000",
6442 => "00000000",
6443 => "00000000",
6444 => "00000000",
6445 => "00011001",
6446 => "01101010",
6447 => "01100010",
6448 => "01100010",
6449 => "01100010",
6450 => "01100010",
6451 => "01100010",
6452 => "01100010",
6453 => "01100010",
6454 => "01100010",
6455 => "01100010",
6456 => "01100010",
6457 => "01100010",
6458 => "01100010",
6459 => "01100010",
6460 => "01100010",
6461 => "01100010",
6462 => "01100010",
6463 => "01100010",
6464 => "01100010",
6465 => "01100010",
6466 => "00010001",
6467 => "00001000",
6468 => "00000000",
6469 => "00000000",
6470 => "00000000",
6471 => "00000000",
6472 => "00000000",
6473 => "00000000",
6474 => "00000000",
6475 => "00000000",
6476 => "00000000",
6477 => "00000000",
6478 => "00000000",
6479 => "00000000",
6480 => "00000000",
6481 => "01011011",
6482 => "10110110",
6483 => "01001000",
6484 => "01010000",
6485 => "10010000",
6486 => "10010000",
6487 => "10011000",
6488 => "10011000",
6489 => "10100000",
6490 => "10100000",
6491 => "10100000",
6492 => "10100000",
6493 => "11101000",
6494 => "11100000",
6495 => "10100011",
6496 => "11110111",
6497 => "11110110",
6498 => "10100100",
6499 => "10100010",
6500 => "10100000",
6501 => "10100000",
6502 => "10100000",
6503 => "11100000",
6504 => "11101000",
6505 => "11101000",
6506 => "10011000",
6507 => "11110110",
6508 => "11110110",
6509 => "10011001",
6510 => "10100000",
6511 => "10100000",
6512 => "10100000",
6513 => "10011000",
6514 => "10011000",
6515 => "10010000",
6516 => "10010000",
6528 => "11101100",
6529 => "11101100",
6530 => "11101100",
6531 => "11101100",
6532 => "10100100",
6533 => "01010010",
6534 => "10100011",
6535 => "10100100",
6536 => "01100100",
6537 => "10100101",
6538 => "00001010",
6539 => "10011010",
6540 => "11101100",
6541 => "11101100",
6542 => "11101100",
6543 => "11101100",
6544 => "11101100",
6545 => "11101100",
6546 => "11101100",
6547 => "11101100",
6548 => "11101100",
6549 => "11101100",
6550 => "11101011",
6551 => "11110110",
6552 => "11111111",
6553 => "10110110",
6554 => "01010010",
6555 => "00000000",
6556 => "00000000",
6557 => "00000000",
6558 => "00000000",
6559 => "00000000",
6560 => "00000000",
6561 => "00000000",
6562 => "00000000",
6563 => "00000000",
6564 => "00000000",
6565 => "00000000",
6566 => "00000000",
6567 => "00000000",
6568 => "00000000",
6569 => "00000000",
6570 => "00000000",
6571 => "00000000",
6572 => "00000000",
6573 => "00010001",
6574 => "01101010",
6575 => "01100010",
6576 => "01100011",
6577 => "01100010",
6578 => "01100010",
6579 => "01100010",
6580 => "01100010",
6581 => "01100010",
6582 => "01100100",
6583 => "01101101",
6584 => "01101101",
6585 => "01100100",
6586 => "01100010",
6587 => "01100010",
6588 => "01100010",
6589 => "01100010",
6590 => "01100010",
6591 => "01100011",
6592 => "01100010",
6593 => "01100010",
6594 => "00000000",
6595 => "00000000",
6596 => "00000000",
6597 => "00000000",
6598 => "00000000",
6599 => "00000000",
6600 => "00000000",
6601 => "00000000",
6602 => "00000000",
6603 => "00000000",
6604 => "00000000",
6605 => "00000000",
6606 => "00000000",
6607 => "00000000",
6608 => "00000000",
6609 => "10100100",
6610 => "10101101",
6611 => "01001000",
6612 => "10010000",
6613 => "10010000",
6614 => "10010000",
6615 => "10011000",
6616 => "10011000",
6617 => "10100000",
6618 => "10100000",
6619 => "10100000",
6620 => "10100000",
6621 => "11101000",
6622 => "11100000",
6623 => "10100010",
6624 => "11111111",
6625 => "10101101",
6626 => "10011000",
6627 => "11101000",
6628 => "11101000",
6629 => "11110000",
6630 => "11110000",
6631 => "11101000",
6632 => "11101000",
6633 => "11101000",
6634 => "10100001",
6635 => "11110110",
6636 => "11110110",
6637 => "10011001",
6638 => "10100000",
6639 => "10100000",
6640 => "10100000",
6641 => "10011000",
6642 => "10011000",
6643 => "10010000",
6644 => "10010000",
6656 => "11101011",
6657 => "11101011",
6658 => "11101011",
6659 => "11101011",
6660 => "11101100",
6661 => "01010010",
6662 => "01011011",
6663 => "10100100",
6664 => "01100100",
6665 => "01100100",
6666 => "01011100",
6667 => "01010010",
6668 => "11101100",
6669 => "11101100",
6670 => "11101100",
6671 => "11101100",
6672 => "11101100",
6673 => "11101100",
6674 => "11101100",
6675 => "11101100",
6676 => "11101100",
6677 => "11101100",
6678 => "11101011",
6679 => "11110110",
6680 => "11111111",
6681 => "11111111",
6682 => "10110101",
6683 => "01011011",
6684 => "01011011",
6685 => "01011011",
6686 => "01011011",
6687 => "01011011",
6688 => "01011011",
6689 => "01011011",
6690 => "01011011",
6691 => "01011011",
6692 => "01011011",
6693 => "01011011",
6694 => "01011011",
6695 => "01011011",
6696 => "01011011",
6697 => "01011011",
6698 => "01011011",
6699 => "01011011",
6700 => "01011011",
6701 => "01011011",
6702 => "01011010",
6703 => "01101101",
6704 => "01100111",
6705 => "01100110",
6706 => "01100101",
6707 => "01100101",
6708 => "01101110",
6709 => "01101110",
6710 => "01101111",
6711 => "10101111",
6712 => "10101111",
6713 => "01101111",
6714 => "01101110",
6715 => "01100101",
6716 => "01100101",
6717 => "01100101",
6718 => "01100110",
6719 => "01101111",
6720 => "01100101",
6721 => "01011001",
6722 => "01011010",
6723 => "01011011",
6724 => "01011011",
6725 => "01011011",
6726 => "01011011",
6727 => "01011011",
6728 => "01011011",
6729 => "01011011",
6730 => "01011011",
6731 => "01011011",
6732 => "01011011",
6733 => "01011011",
6734 => "01011011",
6735 => "01011011",
6736 => "01011011",
6737 => "10101101",
6738 => "10100100",
6739 => "01001000",
6740 => "10010000",
6741 => "10010000",
6742 => "10010000",
6743 => "10011000",
6744 => "10011000",
6745 => "10100000",
6746 => "10100000",
6747 => "10100000",
6748 => "10100000",
6749 => "11101000",
6750 => "11100000",
6751 => "10100010",
6752 => "11111111",
6753 => "10101101",
6754 => "10100000",
6755 => "11110000",
6756 => "11101000",
6757 => "11101000",
6758 => "11101000",
6759 => "11101000",
6760 => "11101000",
6761 => "11101000",
6762 => "10100001",
6763 => "11110110",
6764 => "11110110",
6765 => "10011001",
6766 => "10100000",
6767 => "10100000",
6768 => "10100000",
6769 => "10011000",
6770 => "10011000",
6771 => "10010000",
6772 => "10010000",
6784 => "11101011",
6785 => "11101011",
6786 => "11101011",
6787 => "11101011",
6788 => "11101011",
6789 => "10011011",
6790 => "00001010",
6791 => "01011011",
6792 => "01011011",
6793 => "01011100",
6794 => "01011100",
6795 => "01100101",
6796 => "10100100",
6797 => "10100011",
6798 => "10011011",
6799 => "11101100",
6800 => "11101100",
6801 => "11101100",
6802 => "11101011",
6803 => "11101011",
6804 => "11101011",
6805 => "11101011",
6806 => "11100011",
6807 => "11110101",
6808 => "11111111",
6809 => "11111111",
6810 => "01011011",
6811 => "01011011",
6812 => "01011011",
6813 => "01011011",
6814 => "01011011",
6815 => "01011011",
6816 => "01011011",
6817 => "01011011",
6818 => "01011011",
6819 => "01011011",
6820 => "01011011",
6821 => "01011011",
6822 => "01011011",
6823 => "01011011",
6824 => "01011011",
6825 => "01011011",
6826 => "01011011",
6827 => "01011011",
6828 => "01011011",
6829 => "01011011",
6830 => "01011011",
6831 => "01011100",
6832 => "01100101",
6833 => "01100110",
6834 => "01101111",
6835 => "01101111",
6836 => "01101111",
6837 => "01101111",
6838 => "01101111",
6839 => "01101111",
6840 => "01101111",
6841 => "01101111",
6842 => "01101111",
6843 => "01101111",
6844 => "01101111",
6845 => "01101111",
6846 => "01100110",
6847 => "01100101",
6848 => "01100100",
6849 => "01011011",
6850 => "01011011",
6851 => "01011011",
6852 => "01011011",
6853 => "01011011",
6854 => "01011011",
6855 => "01011011",
6856 => "01011011",
6857 => "01011011",
6858 => "01011011",
6859 => "01011011",
6860 => "01011011",
6861 => "01011011",
6862 => "01011011",
6863 => "01011011",
6864 => "01011011",
6865 => "10101101",
6866 => "10100100",
6867 => "01001000",
6868 => "10010000",
6869 => "10010000",
6870 => "10011000",
6871 => "10011000",
6872 => "10011000",
6873 => "10100000",
6874 => "10100000",
6875 => "10100000",
6876 => "10100000",
6877 => "11101000",
6878 => "11100000",
6879 => "10100010",
6880 => "11111111",
6881 => "10101101",
6882 => "10100000",
6883 => "11110000",
6884 => "11110000",
6885 => "11110000",
6886 => "11101000",
6887 => "11101000",
6888 => "11101000",
6889 => "11101000",
6890 => "10100000",
6891 => "11110110",
6892 => "11110110",
6893 => "10011000",
6894 => "10100000",
6895 => "10100000",
6896 => "10011000",
6897 => "10011000",
6898 => "10011000",
6899 => "10010000",
6900 => "10010000",
6912 => "11101011",
6913 => "11101100",
6914 => "11101011",
6915 => "11100011",
6916 => "11101011",
6917 => "11101011",
6918 => "01010010",
6919 => "01010010",
6920 => "01010011",
6921 => "01010011",
6922 => "01100100",
6923 => "10110110",
6924 => "01011011",
6925 => "00000001",
6926 => "01010010",
6927 => "11101011",
6928 => "11101011",
6929 => "11101011",
6930 => "11101011",
6931 => "11101011",
6932 => "11101011",
6933 => "11101011",
6934 => "11100011",
6935 => "11101100",
6936 => "11111111",
6937 => "11111111",
6938 => "10101101",
6939 => "01011011",
6940 => "01011011",
6941 => "01011011",
6942 => "01011011",
6943 => "01011011",
6944 => "01011011",
6945 => "01011011",
6946 => "01011011",
6947 => "01011011",
6948 => "01011011",
6949 => "01011011",
6950 => "01011011",
6951 => "01011011",
6952 => "01011011",
6953 => "01011011",
6954 => "01011011",
6955 => "01011011",
6956 => "01011011",
6957 => "01011011",
6958 => "01011011",
6959 => "01011011",
6960 => "01011011",
6961 => "01100111",
6962 => "01100111",
6963 => "01101111",
6964 => "01101111",
6965 => "01101111",
6966 => "01101111",
6967 => "01101111",
6968 => "01101111",
6969 => "01101111",
6970 => "01101111",
6971 => "01101111",
6972 => "01101111",
6973 => "01100111",
6974 => "01100110",
6975 => "01011011",
6976 => "01011011",
6977 => "01011011",
6978 => "01011011",
6979 => "01011011",
6980 => "01011011",
6981 => "01011011",
6982 => "01011011",
6983 => "01011011",
6984 => "01011011",
6985 => "01011011",
6986 => "01011011",
6987 => "01011011",
6988 => "01011011",
6989 => "01011011",
6990 => "01011011",
6991 => "01011011",
6992 => "01011011",
6993 => "10101101",
6994 => "10100100",
6995 => "01001000",
6996 => "10010000",
6997 => "10010000",
6998 => "10011000",
6999 => "10011000",
7000 => "10011000",
7001 => "10100000",
7002 => "10100000",
7003 => "10100000",
7004 => "11100000",
7005 => "11101000",
7006 => "11100000",
7007 => "10100010",
7008 => "11111111",
7009 => "10101101",
7010 => "10100000",
7011 => "11110000",
7012 => "11110000",
7013 => "11110000",
7014 => "11110000",
7015 => "11101000",
7016 => "11101000",
7017 => "11101000",
7018 => "10100001",
7019 => "11110110",
7020 => "11110110",
7021 => "10011000",
7022 => "10100000",
7023 => "10100000",
7024 => "10011000",
7025 => "10011000",
7026 => "10011000",
7027 => "10010000",
7028 => "10010000",
7040 => "11100011",
7041 => "11101011",
7042 => "11101011",
7043 => "11100011",
7044 => "11100011",
7045 => "11101011",
7046 => "10100011",
7047 => "01001001",
7048 => "01010010",
7049 => "01100100",
7050 => "10101110",
7051 => "10101101",
7052 => "01100100",
7053 => "00010010",
7054 => "10100011",
7055 => "11101100",
7056 => "11101011",
7057 => "11101011",
7058 => "11101011",
7059 => "11101011",
7060 => "11101011",
7061 => "11101011",
7062 => "11100011",
7063 => "11101100",
7064 => "11111111",
7065 => "11111111",
7066 => "11111111",
7067 => "10100100",
7068 => "01011011",
7069 => "01011011",
7070 => "01011011",
7071 => "01011011",
7072 => "01011011",
7073 => "01011011",
7074 => "01011011",
7075 => "01011011",
7076 => "01011011",
7077 => "01011011",
7078 => "01011011",
7079 => "01011011",
7080 => "01011011",
7081 => "01011011",
7082 => "01011011",
7083 => "01011011",
7084 => "01011011",
7085 => "01011011",
7086 => "01011011",
7087 => "01011011",
7088 => "01100101",
7089 => "01101111",
7090 => "01100110",
7091 => "01100110",
7092 => "01100110",
7093 => "01100110",
7094 => "01100110",
7095 => "01100110",
7096 => "01100110",
7097 => "01100110",
7098 => "01100110",
7099 => "01100110",
7100 => "01100110",
7101 => "01100110",
7102 => "01101111",
7103 => "01011101",
7104 => "01011011",
7105 => "01011011",
7106 => "01011011",
7107 => "01011011",
7108 => "01011011",
7109 => "01011011",
7110 => "01011011",
7111 => "01011011",
7112 => "01011011",
7113 => "01011011",
7114 => "01011011",
7115 => "01011011",
7116 => "01011011",
7117 => "01011011",
7118 => "01011011",
7119 => "01011011",
7120 => "01011011",
7121 => "10101101",
7122 => "10100100",
7123 => "01001000",
7124 => "10010000",
7125 => "10010000",
7126 => "10011000",
7127 => "10011000",
7128 => "10011000",
7129 => "10100000",
7130 => "10100000",
7131 => "10100000",
7132 => "11100000",
7133 => "11101000",
7134 => "11100000",
7135 => "10100010",
7136 => "11110111",
7137 => "10101101",
7138 => "10100000",
7139 => "11110000",
7140 => "11110000",
7141 => "11110000",
7142 => "11110000",
7143 => "11101000",
7144 => "11101000",
7145 => "11100000",
7146 => "10011000",
7147 => "11110110",
7148 => "11110110",
7149 => "10011000",
7150 => "10100000",
7151 => "10100000",
7152 => "10011000",
7153 => "10011000",
7154 => "10011000",
7155 => "10010000",
7156 => "10010000",
7168 => "11100011",
7169 => "11101011",
7170 => "11101011",
7171 => "11101011",
7172 => "11100011",
7173 => "11100011",
7174 => "11101011",
7175 => "10100011",
7176 => "01011011",
7177 => "01100101",
7178 => "01010011",
7179 => "00010010",
7180 => "01011100",
7181 => "00010011",
7182 => "01010010",
7183 => "10100011",
7184 => "11101011",
7185 => "11100011",
7186 => "11100011",
7187 => "11101011",
7188 => "11101011",
7189 => "11101011",
7190 => "11101011",
7191 => "11101011",
7192 => "11111110",
7193 => "11111111",
7194 => "10101101",
7195 => "01011011",
7196 => "01011011",
7197 => "01011011",
7198 => "01011011",
7199 => "01011011",
7200 => "01011011",
7201 => "01011011",
7202 => "01011011",
7203 => "01011011",
7204 => "01011011",
7205 => "01011011",
7206 => "01011011",
7207 => "01011011",
7208 => "01011011",
7209 => "01011011",
7210 => "01011011",
7211 => "01011011",
7212 => "01011011",
7213 => "01011011",
7214 => "01011011",
7215 => "01011010",
7216 => "01100100",
7217 => "01100101",
7218 => "00011101",
7219 => "00011101",
7220 => "00011101",
7221 => "01011110",
7222 => "01011110",
7223 => "01100110",
7224 => "01100110",
7225 => "01011110",
7226 => "01011101",
7227 => "00011101",
7228 => "00011101",
7229 => "00011101",
7230 => "01100101",
7231 => "01011100",
7232 => "01011011",
7233 => "01011011",
7234 => "01011011",
7235 => "01011011",
7236 => "01011011",
7237 => "01011011",
7238 => "01011011",
7239 => "01011011",
7240 => "01011011",
7241 => "01011011",
7242 => "01011011",
7243 => "01011011",
7244 => "01011011",
7245 => "01011011",
7246 => "01011011",
7247 => "01011011",
7248 => "01011011",
7249 => "10101101",
7250 => "10101100",
7251 => "01001000",
7252 => "10010000",
7253 => "10010000",
7254 => "10011000",
7255 => "10011000",
7256 => "10011000",
7257 => "10100000",
7258 => "10100000",
7259 => "10100000",
7260 => "11100000",
7261 => "11101000",
7262 => "11100000",
7263 => "10100010",
7264 => "11110110",
7265 => "10101101",
7266 => "10100000",
7267 => "11110000",
7268 => "11110000",
7269 => "11110000",
7270 => "11101000",
7271 => "11101000",
7272 => "10101010",
7273 => "10101011",
7274 => "10100011",
7275 => "11110110",
7276 => "10110110",
7277 => "10011000",
7278 => "10100000",
7279 => "10100000",
7280 => "10011000",
7281 => "10011000",
7282 => "10011000",
7283 => "10010000",
7284 => "10010000",
7296 => "11100011",
7297 => "11100011",
7298 => "11100011",
7299 => "11100011",
7300 => "11100011",
7301 => "10100011",
7302 => "10011011",
7303 => "01011011",
7304 => "01100101",
7305 => "01011011",
7306 => "01011011",
7307 => "01010011",
7308 => "00010011",
7309 => "01011011",
7310 => "00010011",
7311 => "00001001",
7312 => "10011010",
7313 => "11101011",
7314 => "11101011",
7315 => "11101011",
7316 => "11101011",
7317 => "11101011",
7318 => "11101011",
7319 => "11100011",
7320 => "11110110",
7321 => "11111111",
7322 => "11111111",
7323 => "10101101",
7324 => "01011011",
7325 => "01011011",
7326 => "10100011",
7327 => "10100011",
7328 => "10100011",
7329 => "10100011",
7330 => "10100011",
7331 => "10100011",
7332 => "10100011",
7333 => "10100011",
7334 => "10100011",
7335 => "01011011",
7336 => "01011011",
7337 => "01011011",
7338 => "01011011",
7339 => "01011011",
7340 => "01011011",
7341 => "01011011",
7342 => "01010010",
7343 => "01101010",
7344 => "01101011",
7345 => "01100010",
7346 => "01100011",
7347 => "00011101",
7348 => "01011100",
7349 => "01011100",
7350 => "01011011",
7351 => "01011011",
7352 => "01011011",
7353 => "01100011",
7354 => "01011100",
7355 => "01011100",
7356 => "00011100",
7357 => "01100011",
7358 => "01101010",
7359 => "01101011",
7360 => "01100010",
7361 => "01011011",
7362 => "01011011",
7363 => "01011011",
7364 => "01011011",
7365 => "01011011",
7366 => "01011011",
7367 => "01011011",
7368 => "01011011",
7369 => "01011011",
7370 => "10100011",
7371 => "01100011",
7372 => "01011011",
7373 => "01011011",
7374 => "01011011",
7375 => "01011011",
7376 => "01011011",
7377 => "10101100",
7378 => "10101101",
7379 => "01010000",
7380 => "10010000",
7381 => "10010000",
7382 => "10011000",
7383 => "10011000",
7384 => "10011000",
7385 => "10100000",
7386 => "10100000",
7387 => "10100000",
7388 => "11101000",
7389 => "11101000",
7390 => "11100000",
7391 => "10100010",
7392 => "10110110",
7393 => "10101100",
7394 => "10100000",
7395 => "11110000",
7396 => "11110000",
7397 => "11101000",
7398 => "10100001",
7399 => "10101101",
7400 => "10110110",
7401 => "11110110",
7402 => "11110110",
7403 => "11110110",
7404 => "10110110",
7405 => "10011001",
7406 => "10100000",
7407 => "10100000",
7408 => "10011000",
7409 => "10011000",
7410 => "10011000",
7411 => "10010000",
7412 => "10010000",
7424 => "11101011",
7425 => "11101011",
7426 => "11101011",
7427 => "11101011",
7428 => "01011011",
7429 => "00010011",
7430 => "01010011",
7431 => "01011011",
7432 => "01010011",
7433 => "00010010",
7434 => "00010011",
7435 => "00001010",
7436 => "00010010",
7437 => "01011011",
7438 => "01011011",
7439 => "01010011",
7440 => "00001001",
7441 => "01010010",
7442 => "10100011",
7443 => "10100011",
7444 => "11101011",
7445 => "11100011",
7446 => "11101011",
7447 => "11100011",
7448 => "11110101",
7449 => "11111111",
7450 => "11111111",
7451 => "10101101",
7452 => "01011011",
7453 => "01011011",
7454 => "10100011",
7455 => "10100011",
7456 => "10100011",
7457 => "10100011",
7458 => "10100011",
7459 => "10100011",
7460 => "10100011",
7461 => "10100011",
7462 => "10100011",
7463 => "10100011",
7464 => "10100011",
7465 => "01011011",
7466 => "01011011",
7467 => "01011011",
7468 => "01011011",
7469 => "01011011",
7470 => "01100010",
7471 => "01101011",
7472 => "01100010",
7473 => "01100010",
7474 => "01100010",
7475 => "01100010",
7476 => "01100001",
7477 => "01100001",
7478 => "01100001",
7479 => "01100001",
7480 => "01100001",
7481 => "01100001",
7482 => "01100001",
7483 => "01100001",
7484 => "01100010",
7485 => "01100010",
7486 => "01100010",
7487 => "01101011",
7488 => "01101011",
7489 => "01011010",
7490 => "01011011",
7491 => "01011011",
7492 => "01011011",
7493 => "01011011",
7494 => "01011011",
7495 => "01011011",
7496 => "10100011",
7497 => "10100011",
7498 => "10100011",
7499 => "10100011",
7500 => "01100011",
7501 => "01011011",
7502 => "01011011",
7503 => "01011011",
7504 => "01011011",
7505 => "10100100",
7506 => "10110110",
7507 => "01010001",
7508 => "10010000",
7509 => "10010000",
7510 => "10011000",
7511 => "10011000",
7512 => "10011000",
7513 => "10100000",
7514 => "10100000",
7515 => "10100000",
7516 => "10100000",
7517 => "10100000",
7518 => "10100000",
7519 => "10100011",
7520 => "10110110",
7521 => "10100100",
7522 => "10100000",
7523 => "11110000",
7524 => "11101000",
7525 => "10101000",
7526 => "10101101",
7527 => "10110110",
7528 => "10101101",
7529 => "10101101",
7530 => "10101101",
7531 => "10110110",
7532 => "10101110",
7533 => "10011001",
7534 => "10100000",
7535 => "10100000",
7536 => "10011000",
7537 => "10011000",
7538 => "10011000",
7539 => "10010000",
7540 => "10010000",
7552 => "11101011",
7553 => "11101011",
7554 => "11100011",
7555 => "11101011",
7556 => "01011100",
7557 => "00010011",
7558 => "01010011",
7559 => "01011011",
7560 => "01011011",
7561 => "01011100",
7562 => "00010010",
7563 => "01001010",
7564 => "01010010",
7565 => "01010011",
7566 => "01011011",
7567 => "01011011",
7568 => "01011100",
7569 => "01011011",
7570 => "01011100",
7571 => "01010011",
7572 => "10011010",
7573 => "11101011",
7574 => "11101011",
7575 => "11100011",
7576 => "11101101",
7577 => "11111111",
7578 => "11111111",
7579 => "01011011",
7580 => "01011011",
7581 => "10100011",
7582 => "10100011",
7583 => "10100011",
7584 => "10100011",
7585 => "10100011",
7586 => "10100011",
7587 => "10100100",
7588 => "10100100",
7589 => "10100011",
7590 => "10100011",
7591 => "10100011",
7592 => "10100011",
7593 => "10100011",
7594 => "01011011",
7595 => "01011011",
7596 => "01011011",
7597 => "01011010",
7598 => "01110011",
7599 => "01100010",
7600 => "01100010",
7601 => "01101011",
7602 => "01101011",
7603 => "01100010",
7604 => "01100010",
7605 => "01100010",
7606 => "01101011",
7607 => "01100010",
7608 => "01100011",
7609 => "01100010",
7610 => "01100010",
7611 => "01100010",
7612 => "01100010",
7613 => "01100010",
7614 => "01100010",
7615 => "01100010",
7616 => "01101011",
7617 => "01101011",
7618 => "01011011",
7619 => "01011011",
7620 => "01011011",
7621 => "01011011",
7622 => "01011011",
7623 => "10100011",
7624 => "10100011",
7625 => "10100011",
7626 => "10100011",
7627 => "10100011",
7628 => "10100011",
7629 => "10100011",
7630 => "01011011",
7631 => "01011011",
7632 => "01011011",
7633 => "01011011",
7634 => "11110110",
7635 => "01011010",
7636 => "01010000",
7637 => "10010000",
7638 => "10010000",
7639 => "10011000",
7640 => "10011000",
7641 => "10100000",
7642 => "10100000",
7643 => "10011000",
7644 => "10100100",
7645 => "10101101",
7646 => "10101101",
7647 => "10101101",
7648 => "10101101",
7649 => "10100100",
7650 => "10100000",
7651 => "11101000",
7652 => "11101000",
7653 => "10100001",
7654 => "10101101",
7655 => "10101101",
7656 => "10101101",
7657 => "10101101",
7658 => "10101101",
7659 => "10110110",
7660 => "10101110",
7661 => "10011000",
7662 => "10100000",
7663 => "10100000",
7664 => "10011000",
7665 => "10011000",
7666 => "10011000",
7667 => "10010000",
7668 => "10010000",
7680 => "11101011",
7681 => "11100011",
7682 => "10100010",
7683 => "11101011",
7684 => "10100100",
7685 => "01011100",
7686 => "00010011",
7687 => "01010010",
7688 => "01011100",
7689 => "01011100",
7690 => "01010011",
7691 => "00001001",
7692 => "01010010",
7693 => "01010010",
7694 => "01010010",
7695 => "01010010",
7696 => "01010010",
7697 => "01010011",
7698 => "01011100",
7699 => "01010011",
7700 => "01010010",
7701 => "10100011",
7702 => "10100011",
7703 => "11100011",
7704 => "11101100",
7705 => "11111111",
7706 => "11111111",
7707 => "11110110",
7708 => "10100100",
7709 => "10100011",
7710 => "10100100",
7711 => "10100100",
7712 => "10100100",
7713 => "10100100",
7714 => "10100100",
7715 => "10100100",
7716 => "10100100",
7717 => "10100100",
7718 => "10100100",
7719 => "10100100",
7720 => "10100011",
7721 => "10100011",
7722 => "01011011",
7723 => "01011011",
7724 => "01011011",
7725 => "01101010",
7726 => "01101011",
7727 => "01100010",
7728 => "01101011",
7729 => "01101011",
7730 => "01100010",
7731 => "01100010",
7732 => "01100010",
7733 => "01101011",
7734 => "01101011",
7735 => "01100010",
7736 => "01101011",
7737 => "01101011",
7738 => "01101011",
7739 => "01100010",
7740 => "01100010",
7741 => "01100010",
7742 => "01100010",
7743 => "01100010",
7744 => "01100010",
7745 => "01101011",
7746 => "01100010",
7747 => "01011011",
7748 => "01011011",
7749 => "01011011",
7750 => "10100011",
7751 => "10100100",
7752 => "10100100",
7753 => "10100100",
7754 => "10100100",
7755 => "10100100",
7756 => "10100100",
7757 => "10100011",
7758 => "10100011",
7759 => "01011011",
7760 => "01011011",
7761 => "01011011",
7762 => "10101101",
7763 => "10100100",
7764 => "01010000",
7765 => "10010000",
7766 => "10010000",
7767 => "10011000",
7768 => "10011000",
7769 => "10011000",
7770 => "10011000",
7771 => "10101101",
7772 => "10110110",
7773 => "10101101",
7774 => "10101101",
7775 => "10101101",
7776 => "10101101",
7777 => "10100100",
7778 => "10100000",
7779 => "11101000",
7780 => "11101000",
7781 => "10100001",
7782 => "10101101",
7783 => "10101101",
7784 => "10101101",
7785 => "10101101",
7786 => "10101101",
7787 => "10110110",
7788 => "10100100",
7789 => "10011000",
7790 => "10100000",
7791 => "10100000",
7792 => "10011000",
7793 => "10011000",
7794 => "10010000",
7795 => "10010000",
7796 => "10010000",
7808 => "11100010",
7809 => "11100010",
7810 => "11100010",
7811 => "11100011",
7812 => "11101011",
7813 => "10100011",
7814 => "01010011",
7815 => "01010011",
7816 => "01010011",
7817 => "01011100",
7818 => "01100100",
7819 => "01011011",
7820 => "00001001",
7821 => "01010010",
7822 => "01011011",
7823 => "01011011",
7824 => "01011011",
7825 => "01010011",
7826 => "01010011",
7827 => "01010010",
7828 => "01010011",
7829 => "01011100",
7830 => "10011011",
7831 => "10100011",
7832 => "11101011",
7833 => "11111111",
7834 => "11111111",
7835 => "11110110",
7836 => "10100100",
7837 => "10100011",
7838 => "10100100",
7839 => "10100100",
7840 => "10100100",
7841 => "10100100",
7842 => "10100100",
7843 => "10100100",
7844 => "10100100",
7845 => "10100100",
7846 => "10100100",
7847 => "10100100",
7848 => "10100100",
7849 => "10100011",
7850 => "01011011",
7851 => "01011011",
7852 => "01011010",
7853 => "01101011",
7854 => "01100010",
7855 => "01100010",
7856 => "01101011",
7857 => "01101011",
7858 => "01100010",
7859 => "01100010",
7860 => "01100011",
7861 => "01101011",
7862 => "01101011",
7863 => "01101011",
7864 => "01101011",
7865 => "01101011",
7866 => "01101011",
7867 => "01101011",
7868 => "01100010",
7869 => "01100010",
7870 => "01101011",
7871 => "01100010",
7872 => "01100010",
7873 => "01101011",
7874 => "01101010",
7875 => "01011011",
7876 => "01011011",
7877 => "10100011",
7878 => "10100011",
7879 => "10100100",
7880 => "10100100",
7881 => "10100100",
7882 => "10100100",
7883 => "10100100",
7884 => "10100100",
7885 => "10100100",
7886 => "10100100",
7887 => "10100011",
7888 => "01011011",
7889 => "01011011",
7890 => "10100100",
7891 => "10110110",
7892 => "01010001",
7893 => "10010000",
7894 => "10010000",
7895 => "10011000",
7896 => "10011000",
7897 => "10011000",
7898 => "10011010",
7899 => "10110110",
7900 => "10101101",
7901 => "10101101",
7902 => "10101101",
7903 => "10101101",
7904 => "10101101",
7905 => "10100100",
7906 => "10100000",
7907 => "11101000",
7908 => "11101000",
7909 => "10100000",
7910 => "10011011",
7911 => "10101101",
7912 => "10101101",
7913 => "10101101",
7914 => "10101110",
7915 => "10100100",
7916 => "10011000",
7917 => "10100000",
7918 => "10100000",
7919 => "10011000",
7920 => "10011000",
7921 => "10011000",
7922 => "10010000",
7923 => "10010000",
7924 => "01010000",
7936 => "10011001",
7937 => "10100010",
7938 => "10100010",
7939 => "10011001",
7940 => "11100010",
7941 => "11101011",
7942 => "10100011",
7943 => "10100100",
7944 => "01011011",
7945 => "01011100",
7946 => "10100100",
7947 => "11100011",
7948 => "10100010",
7949 => "01001010",
7950 => "00001010",
7951 => "01010010",
7952 => "01010010",
7953 => "01010010",
7954 => "01010010",
7955 => "01010010",
7956 => "01011011",
7957 => "01011011",
7958 => "01011010",
7959 => "10100011",
7960 => "11100011",
7961 => "11110110",
7962 => "11111111",
7963 => "10101101",
7964 => "01011011",
7965 => "10100100",
7966 => "10100100",
7967 => "10100100",
7968 => "10100100",
7969 => "10100100",
7970 => "10100100",
7971 => "10100100",
7972 => "10100100",
7973 => "10100100",
7974 => "10100100",
7975 => "10100100",
7976 => "10100100",
7977 => "10100100",
7978 => "01011011",
7979 => "01011011",
7980 => "01100010",
7981 => "01101011",
7982 => "01100010",
7983 => "01100010",
7984 => "01101011",
7985 => "01100010",
7986 => "01100010",
7987 => "01100010",
7988 => "01101011",
7989 => "01101011",
7990 => "01101011",
7991 => "01101011",
7992 => "01101011",
7993 => "01101011",
7994 => "01101011",
7995 => "01101011",
7996 => "01100010",
7997 => "01100010",
7998 => "01100010",
7999 => "01101011",
8000 => "01100010",
8001 => "01100010",
8002 => "01101011",
8003 => "01100011",
8004 => "01011011",
8005 => "10100100",
8006 => "10100100",
8007 => "10100100",
8008 => "10100100",
8009 => "10100100",
8010 => "10100100",
8011 => "10100100",
8012 => "10100100",
8013 => "10100100",
8014 => "10100100",
8015 => "10100011",
8016 => "01011011",
8017 => "01011011",
8018 => "01011011",
8019 => "10110110",
8020 => "10100011",
8021 => "01010000",
8022 => "10010000",
8023 => "10010000",
8024 => "10011000",
8025 => "10010000",
8026 => "10011011",
8027 => "10101110",
8028 => "10101101",
8029 => "10101101",
8030 => "10101101",
8031 => "10101101",
8032 => "10101101",
8033 => "10100011",
8034 => "10100000",
8035 => "11101000",
8036 => "11101000",
8037 => "11101000",
8038 => "10100000",
8039 => "10011001",
8040 => "10011011",
8041 => "10011011",
8042 => "10011010",
8043 => "10011000",
8044 => "10100000",
8045 => "10100000",
8046 => "10100000",
8047 => "10011000",
8048 => "10011000",
8049 => "10011000",
8050 => "10010000",
8051 => "10010000",
8052 => "01010001",
8064 => "10011001",
8065 => "10100010",
8066 => "10011001",
8067 => "10100010",
8068 => "11100011",
8069 => "11100011",
8070 => "11101011",
8071 => "11101011",
8072 => "11100010",
8073 => "11100011",
8074 => "11101011",
8075 => "11100011",
8076 => "11100010",
8077 => "10100011",
8078 => "01010010",
8079 => "01010010",
8080 => "01011011",
8081 => "01010011",
8082 => "01010011",
8083 => "01010011",
8084 => "01011011",
8085 => "01011011",
8086 => "01011010",
8087 => "10100011",
8088 => "11100011",
8089 => "11110110",
8090 => "11111111",
8091 => "11111111",
8092 => "10101101",
8093 => "10100011",
8094 => "10100100",
8095 => "10100100",
8096 => "10100100",
8097 => "10100100",
8098 => "10100100",
8099 => "10100100",
8100 => "10100100",
8101 => "10100100",
8102 => "10100100",
8103 => "10100100",
8104 => "10100100",
8105 => "10100100",
8106 => "10100011",
8107 => "01011011",
8108 => "01101010",
8109 => "01101010",
8110 => "01100010",
8111 => "01100010",
8112 => "01100010",
8113 => "01100010",
8114 => "01100010",
8115 => "01101011",
8116 => "01101011",
8117 => "01101011",
8118 => "01101011",
8119 => "01101011",
8120 => "01101011",
8121 => "01101011",
8122 => "01101011",
8123 => "01101011",
8124 => "01101011",
8125 => "01100010",
8126 => "01100010",
8127 => "01100010",
8128 => "01100010",
8129 => "01100010",
8130 => "01101011",
8131 => "01100011",
8132 => "10100011",
8133 => "10100100",
8134 => "10100100",
8135 => "10100100",
8136 => "10100100",
8137 => "10100100",
8138 => "10100100",
8139 => "10100100",
8140 => "10100100",
8141 => "10100100",
8142 => "10100100",
8143 => "10100100",
8144 => "01011011",
8145 => "01011011",
8146 => "01011011",
8147 => "10100100",
8148 => "10110110",
8149 => "01010010",
8150 => "10010000",
8151 => "10010000",
8152 => "10011000",
8153 => "10011000",
8154 => "01010001",
8155 => "10101101",
8156 => "10101101",
8157 => "10101101",
8158 => "10101101",
8159 => "10101101",
8160 => "10100101",
8161 => "10011001",
8162 => "11101000",
8163 => "11101000",
8164 => "11101000",
8165 => "11101000",
8166 => "11101000",
8167 => "11100000",
8168 => "10100000",
8169 => "10100000",
8170 => "10100000",
8171 => "10100000",
8172 => "10100000",
8173 => "10100000",
8174 => "10011000",
8175 => "10011000",
8176 => "10011000",
8177 => "10010000",
8178 => "10010000",
8179 => "01010000",
8180 => "01011011",
8192 => "10011001",
8193 => "10100010",
8194 => "10011001",
8195 => "10100010",
8196 => "11100011",
8197 => "11101011",
8198 => "11100011",
8199 => "11100011",
8200 => "11100010",
8201 => "11100011",
8202 => "11100011",
8203 => "11100011",
8204 => "10100010",
8205 => "11100010",
8206 => "11100011",
8207 => "10100010",
8208 => "10011010",
8209 => "01011010",
8210 => "01010010",
8211 => "01010010",
8212 => "01010010",
8213 => "01010010",
8214 => "10011010",
8215 => "10100011",
8216 => "11100010",
8217 => "11101101",
8218 => "11111111",
8219 => "11111110",
8220 => "10100100",
8221 => "10100011",
8222 => "10100100",
8223 => "10100100",
8224 => "10100100",
8225 => "10100100",
8226 => "10100100",
8227 => "10100100",
8228 => "10100100",
8229 => "10100100",
8230 => "10100100",
8231 => "10100100",
8232 => "10100100",
8233 => "10100100",
8234 => "10100100",
8235 => "01011011",
8236 => "01101010",
8237 => "01101010",
8238 => "01100010",
8239 => "01100010",
8240 => "01100010",
8241 => "01100010",
8242 => "01100011",
8243 => "01101011",
8244 => "01101011",
8245 => "01101011",
8246 => "01101011",
8247 => "01101011",
8248 => "01101011",
8249 => "01101011",
8250 => "01101011",
8251 => "01101011",
8252 => "01100010",
8253 => "01100010",
8254 => "01100010",
8255 => "01100010",
8256 => "01100010",
8257 => "01100010",
8258 => "01101011",
8259 => "01100011",
8260 => "10100100",
8261 => "10100100",
8262 => "10100100",
8263 => "10100100",
8264 => "10100100",
8265 => "10100100",
8266 => "10100100",
8267 => "10100100",
8268 => "10100100",
8269 => "10100100",
8270 => "10100100",
8271 => "10100100",
8272 => "10100011",
8273 => "01011011",
8274 => "01011011",
8275 => "01011011",
8276 => "10110101",
8277 => "10100100",
8278 => "01010001",
8279 => "10011000",
8280 => "10011000",
8281 => "10011000",
8282 => "10010000",
8283 => "01010001",
8284 => "10100100",
8285 => "10100101",
8286 => "10100100",
8287 => "10011011",
8288 => "10011001",
8289 => "10100000",
8290 => "11101000",
8291 => "11101000",
8292 => "11101000",
8293 => "11101000",
8294 => "11101000",
8295 => "11101000",
8296 => "11101000",
8297 => "11101000",
8298 => "10100000",
8299 => "10100000",
8300 => "10100000",
8301 => "10100000",
8302 => "10011000",
8303 => "10011000",
8304 => "10011000",
8305 => "10010000",
8306 => "10010000",
8307 => "01010001",
8308 => "10110110",
8320 => "10011010",
8321 => "10011001",
8322 => "10011001",
8323 => "10011001",
8324 => "10100010",
8325 => "11100011",
8326 => "11100011",
8327 => "11100011",
8328 => "10100010",
8329 => "11100011",
8330 => "11100011",
8331 => "11100011",
8332 => "11100010",
8333 => "11100010",
8334 => "11100011",
8335 => "11100011",
8336 => "11101011",
8337 => "11101011",
8338 => "11100011",
8339 => "10100010",
8340 => "10100010",
8341 => "10100010",
8342 => "10100010",
8343 => "11100011",
8344 => "10100010",
8345 => "11101100",
8346 => "11111111",
8347 => "11110110",
8348 => "01011011",
8349 => "10100100",
8350 => "10100100",
8351 => "10100100",
8352 => "10100100",
8353 => "10100100",
8354 => "10100100",
8355 => "10100100",
8356 => "10100100",
8357 => "10100100",
8358 => "10100100",
8359 => "10100100",
8360 => "10100100",
8361 => "10100100",
8362 => "10100100",
8363 => "01011011",
8364 => "01101010",
8365 => "01100010",
8366 => "01100010",
8367 => "00011001",
8368 => "01100010",
8369 => "01100010",
8370 => "01101011",
8371 => "01100010",
8372 => "01100010",
8373 => "01101011",
8374 => "01100010",
8375 => "01101011",
8376 => "01101011",
8377 => "01100010",
8378 => "01101011",
8379 => "01101011",
8380 => "01100010",
8381 => "01100011",
8382 => "01100010",
8383 => "00011010",
8384 => "01100010",
8385 => "01100010",
8386 => "01101010",
8387 => "01101011",
8388 => "10100100",
8389 => "10100100",
8390 => "10100100",
8391 => "10100100",
8392 => "10100100",
8393 => "10100100",
8394 => "10100100",
8395 => "10100100",
8396 => "10100100",
8397 => "10100100",
8398 => "10100100",
8399 => "10100100",
8400 => "10100100",
8401 => "10100011",
8402 => "01011011",
8403 => "01011011",
8404 => "01011011",
8405 => "11110110",
8406 => "01011011",
8407 => "01010000",
8408 => "10011000",
8409 => "10011000",
8410 => "10011000",
8411 => "10011000",
8412 => "10010000",
8413 => "10010000",
8414 => "10011000",
8415 => "10011000",
8416 => "10100000",
8417 => "11101000",
8418 => "11101000",
8419 => "11101000",
8420 => "11101000",
8421 => "11101000",
8422 => "11101000",
8423 => "10101000",
8424 => "10100000",
8425 => "10100000",
8426 => "10100000",
8427 => "10100000",
8428 => "10100000",
8429 => "10011000",
8430 => "10011000",
8431 => "10011000",
8432 => "10010000",
8433 => "10010000",
8434 => "01010001",
8435 => "10101101",
8436 => "10101101",
8448 => "10011010",
8449 => "10011001",
8450 => "10011001",
8451 => "10011001",
8452 => "10100010",
8453 => "11100011",
8454 => "11100011",
8455 => "11100010",
8456 => "11100010",
8457 => "11100011",
8458 => "11101011",
8459 => "11100011",
8460 => "11100010",
8461 => "11100010",
8462 => "11100010",
8463 => "10100010",
8464 => "10100010",
8465 => "10100010",
8466 => "11100010",
8467 => "11100011",
8468 => "11101011",
8469 => "11101100",
8470 => "11101101",
8471 => "11110101",
8472 => "11110110",
8473 => "11110110",
8474 => "11110110",
8475 => "11111111",
8476 => "11110110",
8477 => "10100100",
8478 => "10100100",
8479 => "10100100",
8480 => "10100100",
8481 => "10100100",
8482 => "10100100",
8483 => "10100100",
8484 => "10100100",
8485 => "10100100",
8486 => "10100100",
8487 => "10100100",
8488 => "10100100",
8489 => "10100100",
8490 => "10100100",
8491 => "01011011",
8492 => "01101010",
8493 => "01100010",
8494 => "01100010",
8495 => "00011001",
8496 => "01100010",
8497 => "01100010",
8498 => "01100010",
8499 => "01100010",
8500 => "01100011",
8501 => "01100010",
8502 => "01100011",
8503 => "01100011",
8504 => "01101011",
8505 => "01101011",
8506 => "01101011",
8507 => "01101011",
8508 => "01100010",
8509 => "01100010",
8510 => "01100010",
8511 => "01100010",
8512 => "01100001",
8513 => "01100010",
8514 => "01101010",
8515 => "01100011",
8516 => "10100100",
8517 => "10100100",
8518 => "10100100",
8519 => "10100100",
8520 => "10100100",
8521 => "10100100",
8522 => "10100100",
8523 => "10100100",
8524 => "10100100",
8525 => "10100100",
8526 => "10100100",
8527 => "10100100",
8528 => "10100100",
8529 => "10100100",
8530 => "01011011",
8531 => "01011011",
8532 => "01011011",
8533 => "10100100",
8534 => "11110110",
8535 => "01011010",
8536 => "01010000",
8537 => "10011000",
8538 => "10011000",
8539 => "10011000",
8540 => "10011000",
8541 => "10100000",
8542 => "10100000",
8543 => "10100000",
8544 => "10100000",
8545 => "10100000",
8546 => "10100000",
8547 => "10101000",
8548 => "10101000",
8549 => "10101000",
8550 => "10100000",
8551 => "10100000",
8552 => "10100000",
8553 => "10100000",
8554 => "10100000",
8555 => "10100000",
8556 => "10011000",
8557 => "10011000",
8558 => "10011000",
8559 => "10011000",
8560 => "10010000",
8561 => "01010001",
8562 => "10100100",
8563 => "11110110",
8564 => "01011011",
8576 => "10011010",
8577 => "11011010",
8578 => "10011010",
8579 => "10011010",
8580 => "11100011",
8581 => "11101011",
8582 => "11100011",
8583 => "10100010",
8584 => "11100010",
8585 => "11100011",
8586 => "11100010",
8587 => "10100010",
8588 => "10100010",
8589 => "11100011",
8590 => "11101011",
8591 => "11101100",
8592 => "11101101",
8593 => "11110101",
8594 => "11110110",
8595 => "11111111",
8596 => "11111111",
8597 => "11111111",
8598 => "11111111",
8599 => "11111111",
8600 => "11111111",
8601 => "11111111",
8602 => "11111111",
8603 => "11110110",
8604 => "11111111",
8605 => "10101101",
8606 => "10100100",
8607 => "10100100",
8608 => "10100100",
8609 => "10100100",
8610 => "10100100",
8611 => "10100100",
8612 => "10100100",
8613 => "10100100",
8614 => "10100100",
8615 => "10100100",
8616 => "10100100",
8617 => "10100100",
8618 => "10100100",
8619 => "10100011",
8620 => "01100010",
8621 => "01101010",
8622 => "01011010",
8623 => "00011001",
8624 => "01100010",
8625 => "01100010",
8626 => "01100010",
8627 => "01100010",
8628 => "01100010",
8629 => "01101011",
8630 => "01101011",
8631 => "01101011",
8632 => "01101011",
8633 => "01101011",
8634 => "01101011",
8635 => "01101011",
8636 => "01100011",
8637 => "01100010",
8638 => "01100010",
8639 => "01100010",
8640 => "01011001",
8641 => "01011010",
8642 => "01101010",
8643 => "01100011",
8644 => "10100100",
8645 => "10100100",
8646 => "10100100",
8647 => "10100100",
8648 => "10100100",
8649 => "10100100",
8650 => "10100100",
8651 => "10100100",
8652 => "10100100",
8653 => "10100100",
8654 => "10100100",
8655 => "10100100",
8656 => "10100100",
8657 => "10100100",
8658 => "10100011",
8659 => "01011011",
8660 => "01011011",
8661 => "01010010",
8662 => "10100100",
8663 => "11110110",
8664 => "01011010",
8665 => "01010000",
8666 => "10011000",
8667 => "10011000",
8668 => "10011000",
8669 => "10011000",
8670 => "10100000",
8671 => "10100000",
8672 => "10100000",
8673 => "10100000",
8674 => "10100000",
8675 => "10100000",
8676 => "10100000",
8677 => "10100000",
8678 => "10100000",
8679 => "10100000",
8680 => "10100000",
8681 => "10100000",
8682 => "10100000",
8683 => "10011000",
8684 => "10011000",
8685 => "10011000",
8686 => "10011000",
8687 => "10010000",
8688 => "01010001",
8689 => "10100100",
8690 => "11110110",
8691 => "01011011",
8692 => "01011011",
8704 => "11101100",
8705 => "11100010",
8706 => "11100011",
8707 => "11100010",
8708 => "11100011",
8709 => "11100010",
8710 => "10100010",
8711 => "10100010",
8712 => "11100011",
8713 => "11101100",
8714 => "11101100",
8715 => "10101100",
8716 => "10101101",
8717 => "11110110",
8718 => "11110110",
8719 => "11110110",
8720 => "11110110",
8721 => "11110110",
8722 => "11110110",
8723 => "11110110",
8724 => "11110110",
8725 => "11110110",
8726 => "10110101",
8727 => "11110110",
8728 => "11110110",
8729 => "10100100",
8730 => "11111111",
8731 => "10100100",
8732 => "01011011",
8733 => "10100100",
8734 => "10100100",
8735 => "10100100",
8736 => "10100100",
8737 => "10100100",
8738 => "10100100",
8739 => "10100100",
8740 => "10100100",
8741 => "10100100",
8742 => "10100100",
8743 => "10100100",
8744 => "10100100",
8745 => "10100100",
8746 => "10100100",
8747 => "10100011",
8748 => "01100010",
8749 => "01101010",
8750 => "01011010",
8751 => "00011001",
8752 => "01100010",
8753 => "01100010",
8754 => "01100010",
8755 => "01100010",
8756 => "01100010",
8757 => "01101011",
8758 => "01101011",
8759 => "01101011",
8760 => "01101011",
8761 => "01101011",
8762 => "01101011",
8763 => "01101011",
8764 => "01100011",
8765 => "01100010",
8766 => "01100010",
8767 => "01100010",
8768 => "00011001",
8769 => "01100010",
8770 => "01101010",
8771 => "01100011",
8772 => "10100100",
8773 => "10100100",
8774 => "10100100",
8775 => "10100100",
8776 => "10100100",
8777 => "10100100",
8778 => "10100100",
8779 => "10100100",
8780 => "10100100",
8781 => "10100100",
8782 => "10100100",
8783 => "10100100",
8784 => "10100100",
8785 => "10100100",
8786 => "10100100",
8787 => "10100011",
8788 => "01011011",
8789 => "01011011",
8790 => "01010010",
8791 => "10100100",
8792 => "11110110",
8793 => "10011011",
8794 => "01010001",
8795 => "10011000",
8796 => "10011000",
8797 => "10011000",
8798 => "10011000",
8799 => "10011000",
8800 => "10100000",
8801 => "10100000",
8802 => "10100000",
8803 => "10100000",
8804 => "10100000",
8805 => "10100000",
8806 => "10100000",
8807 => "10100000",
8808 => "10100000",
8809 => "10011000",
8810 => "10011000",
8811 => "10011000",
8812 => "10011000",
8813 => "10011000",
8814 => "01010000",
8815 => "01010001",
8816 => "10100100",
8817 => "11110110",
8818 => "01011011",
8819 => "01011011",
8820 => "01011011",
8832 => "11110101",
8833 => "11100010",
8834 => "11101011",
8835 => "11101011",
8836 => "10101100",
8837 => "10100100",
8838 => "10101101",
8839 => "11110110",
8840 => "10101101",
8841 => "11110110",
8842 => "11110110",
8843 => "10110110",
8844 => "11110110",
8845 => "11111111",
8846 => "11110110",
8847 => "11110110",
8848 => "11111110",
8849 => "10110101",
8850 => "11110110",
8851 => "11111111",
8852 => "10100100",
8853 => "11110110",
8854 => "10100100",
8855 => "10100100",
8856 => "10101101",
8857 => "01011011",
8858 => "10100100",
8859 => "10100011",
8860 => "10100100",
8861 => "10100100",
8862 => "10100100",
8863 => "10100100",
8864 => "10100100",
8865 => "10100100",
8866 => "10100100",
8867 => "10100100",
8868 => "10100100",
8869 => "10100100",
8870 => "10100100",
8871 => "10100100",
8872 => "10100100",
8873 => "10100100",
8874 => "10100100",
8875 => "10100100",
8876 => "01100010",
8877 => "01101010",
8878 => "01010010",
8879 => "01011010",
8880 => "01100010",
8881 => "01100010",
8882 => "01100010",
8883 => "01100010",
8884 => "01100010",
8885 => "01101011",
8886 => "01101011",
8887 => "01101011",
8888 => "01101011",
8889 => "01101011",
8890 => "01101011",
8891 => "01101011",
8892 => "01100011",
8893 => "01100010",
8894 => "01100010",
8895 => "01100010",
8896 => "01011010",
8897 => "01011010",
8898 => "01101010",
8899 => "01100011",
8900 => "10100100",
8901 => "10100100",
8902 => "10100100",
8903 => "10100100",
8904 => "10100100",
8905 => "10100100",
8906 => "10100100",
8907 => "10100100",
8908 => "10100100",
8909 => "10100100",
8910 => "10100100",
8911 => "10100100",
8912 => "10100100",
8913 => "10100100",
8914 => "10100100",
8915 => "10100100",
8916 => "10100100",
8917 => "01011011",
8918 => "01011011",
8919 => "01010010",
8920 => "10100100",
8921 => "11110110",
8922 => "10100100",
8923 => "01010010",
8924 => "01010000",
8925 => "10011000",
8926 => "10011000",
8927 => "10011000",
8928 => "10011000",
8929 => "10011000",
8930 => "10011000",
8931 => "10011000",
8932 => "10011000",
8933 => "10011000",
8934 => "10011000",
8935 => "10011000",
8936 => "10011000",
8937 => "10011000",
8938 => "10011000",
8939 => "10011000",
8940 => "10011000",
8941 => "01010001",
8942 => "01011010",
8943 => "10101101",
8944 => "10110110",
8945 => "01011011",
8946 => "01011011",
8947 => "01011011",
8948 => "10100100",
8960 => "10101101",
8961 => "10101101",
8962 => "10110101",
8963 => "10110101",
8964 => "10110110",
8965 => "11110110",
8966 => "11110110",
8967 => "11110110",
8968 => "11110110",
8969 => "11110110",
8970 => "10101101",
8971 => "11110110",
8972 => "10101101",
8973 => "10101101",
8974 => "11110110",
8975 => "01011011",
8976 => "10101101",
8977 => "01011011",
8978 => "01011011",
8979 => "10100100",
8980 => "01011011",
8981 => "01011011",
8982 => "01011011",
8983 => "01011011",
8984 => "01011011",
8985 => "10011011",
8986 => "01011011",
8987 => "10100011",
8988 => "10100100",
8989 => "10100100",
8990 => "10100100",
8991 => "10100100",
8992 => "10100100",
8993 => "10100100",
8994 => "10100100",
8995 => "10100100",
8996 => "10100100",
8997 => "10100100",
8998 => "10100100",
8999 => "10100100",
9000 => "10100100",
9001 => "10100100",
9002 => "10100100",
9003 => "10100100",
9004 => "01100010",
9005 => "01100010",
9006 => "01010010",
9007 => "01011010",
9008 => "01100010",
9009 => "01100010",
9010 => "01100010",
9011 => "01100010",
9012 => "01100010",
9013 => "01101011",
9014 => "01101011",
9015 => "01101011",
9016 => "01101011",
9017 => "01101011",
9018 => "01101011",
9019 => "01101011",
9020 => "01100011",
9021 => "01100010",
9022 => "01100010",
9023 => "01100010",
9024 => "01011010",
9025 => "01011010",
9026 => "01100010",
9027 => "01100011",
9028 => "10100100",
9029 => "10100100",
9030 => "10100100",
9031 => "10100100",
9032 => "10100100",
9033 => "10100100",
9034 => "10100100",
9035 => "10100100",
9036 => "10100100",
9037 => "10100100",
9038 => "10100100",
9039 => "10100100",
9040 => "10100100",
9041 => "10100100",
9042 => "10100100",
9043 => "10100100",
9044 => "10100100",
9045 => "10100100",
9046 => "01100011",
9047 => "01011011",
9048 => "01011011",
9049 => "01011011",
9050 => "10110101",
9051 => "10110110",
9052 => "10100011",
9053 => "01010010",
9054 => "01010001",
9055 => "10011000",
9056 => "10011000",
9057 => "10011000",
9058 => "10011000",
9059 => "10011000",
9060 => "10011000",
9061 => "10011000",
9062 => "10011000",
9063 => "10011000",
9064 => "10011000",
9065 => "10011000",
9066 => "10010000",
9067 => "01010001",
9068 => "01011010",
9069 => "10100100",
9070 => "11110110",
9071 => "10101101",
9072 => "01011011",
9073 => "01011011",
9074 => "01011011",
9075 => "10100100",
9076 => "10100100",
9088 => "11110110",
9089 => "11110110",
9090 => "11110110",
9091 => "11110110",
9092 => "11110110",
9093 => "10101101",
9094 => "11110110",
9095 => "10101101",
9096 => "10100100",
9097 => "11110110",
9098 => "01011010",
9099 => "10100100",
9100 => "10100100",
9101 => "01011011",
9102 => "01011011",
9103 => "01011011",
9104 => "01011011",
9105 => "01011011",
9106 => "01011011",
9107 => "01011011",
9108 => "01011011",
9109 => "01011011",
9110 => "01011011",
9111 => "01011011",
9112 => "01011011",
9113 => "01011011",
9114 => "10100100",
9115 => "10100100",
9116 => "10100100",
9117 => "10100100",
9118 => "10100100",
9119 => "10100100",
9120 => "10100100",
9121 => "10100100",
9122 => "10100100",
9123 => "10100100",
9124 => "10100100",
9125 => "10100100",
9126 => "10100100",
9127 => "10100100",
9128 => "10100100",
9129 => "10100100",
9130 => "10100100",
9131 => "10100100",
9132 => "01011011",
9133 => "01011010",
9134 => "01010010",
9135 => "01010010",
9136 => "01100010",
9137 => "01100010",
9138 => "01100010",
9139 => "01100010",
9140 => "01100010",
9141 => "01101011",
9142 => "01101011",
9143 => "01101011",
9144 => "01101011",
9145 => "01101011",
9146 => "01101011",
9147 => "01101011",
9148 => "01100010",
9149 => "01100010",
9150 => "01100010",
9151 => "01100010",
9152 => "01010010",
9153 => "01010010",
9154 => "01011010",
9155 => "01100011",
9156 => "10100100",
9157 => "10100100",
9158 => "10100100",
9159 => "10100100",
9160 => "10100100",
9161 => "10100100",
9162 => "10100100",
9163 => "10100100",
9164 => "10100100",
9165 => "10101100",
9166 => "10100100",
9167 => "10100100",
9168 => "10100100",
9169 => "10100100",
9170 => "10100100",
9171 => "10100100",
9172 => "10100100",
9173 => "10100100",
9174 => "10100100",
9175 => "10100100",
9176 => "01011011",
9177 => "01011011",
9178 => "01010010",
9179 => "10100100",
9180 => "10110110",
9181 => "10110110",
9182 => "10100100",
9183 => "01011010",
9184 => "01010001",
9185 => "01010001",
9186 => "01010001",
9187 => "01010000",
9188 => "01010000",
9189 => "01010000",
9190 => "01010001",
9191 => "01010001",
9192 => "01010001",
9193 => "01010010",
9194 => "01011011",
9195 => "10101101",
9196 => "11110110",
9197 => "10101101",
9198 => "01011011",
9199 => "01010010",
9200 => "01011011",
9201 => "10100100",
9202 => "10100100",
9203 => "10100100",
9204 => "10100100",
9216 => "10100100",
9217 => "10101101",
9218 => "10101101",
9219 => "01011011",
9220 => "10101101",
9221 => "01010010",
9222 => "10100011",
9223 => "10100011",
9224 => "01010010",
9225 => "01011011",
9226 => "01011011",
9227 => "01011010",
9228 => "01011011",
9229 => "01011011",
9230 => "01011011",
9231 => "01011011",
9232 => "01011011",
9233 => "01011011",
9234 => "01011011",
9235 => "01011011",
9236 => "01011011",
9237 => "01011011",
9238 => "10011011",
9239 => "10100011",
9240 => "10100011",
9241 => "10100100",
9242 => "10100100",
9243 => "10100100",
9244 => "10100100",
9245 => "10100100",
9246 => "10100100",
9247 => "10100100",
9248 => "10101100",
9249 => "10101100",
9250 => "10101100",
9251 => "10101100",
9252 => "10101100",
9253 => "10101101",
9254 => "10101100",
9255 => "10101100",
9256 => "10100100",
9257 => "10100100",
9258 => "10100100",
9259 => "10100100",
9260 => "10100100",
9261 => "01011011",
9262 => "01010010",
9263 => "01010010",
9264 => "01010010",
9265 => "01011010",
9266 => "01100010",
9267 => "01100010",
9268 => "01100010",
9269 => "01100010",
9270 => "01100011",
9271 => "01100011",
9272 => "01100011",
9273 => "01100011",
9274 => "01100010",
9275 => "01100010",
9276 => "01100010",
9277 => "01100010",
9278 => "01011010",
9279 => "01011010",
9280 => "01010010",
9281 => "01011011",
9282 => "01011011",
9283 => "10100100",
9284 => "10100100",
9285 => "10100100",
9286 => "10100100",
9287 => "10101100",
9288 => "10101100",
9289 => "10101101",
9290 => "10101101",
9291 => "10101100",
9292 => "10101100",
9293 => "10101100",
9294 => "10101101",
9295 => "10101100",
9296 => "10101101",
9297 => "10101100",
9298 => "10101100",
9299 => "10100100",
9300 => "10100100",
9301 => "10100100",
9302 => "10100100",
9303 => "10100100",
9304 => "10100100",
9305 => "10100100",
9306 => "10100011",
9307 => "01011011",
9308 => "01011010",
9309 => "10100100",
9310 => "10101101",
9311 => "11110110",
9312 => "10110101",
9313 => "10101101",
9314 => "10100100",
9315 => "10100100",
9316 => "10100011",
9317 => "10100011",
9318 => "10100100",
9319 => "10101100",
9320 => "10101101",
9321 => "10110110",
9322 => "10110110",
9323 => "10101101",
9324 => "01011011",
9325 => "01010010",
9326 => "01011011",
9327 => "10100100",
9328 => "10100100",
9329 => "10100100",
9330 => "10100100",
9331 => "10100100",
9332 => "10100100",
9344 => "01010010",
9345 => "01011011",
9346 => "01011011",
9347 => "01011011",
9348 => "01011011",
9349 => "01011011",
9350 => "01011011",
9351 => "01011011",
9352 => "01011011",
9353 => "01011011",
9354 => "10100100",
9355 => "10100011",
9356 => "10011011",
9357 => "10100011",
9358 => "10100011",
9359 => "10100011",
9360 => "10100100",
9361 => "10100100",
9362 => "10100100",
9363 => "10100100",
9364 => "10100100",
9365 => "10100100",
9366 => "10100100",
9367 => "10100100",
9368 => "10100100",
9369 => "10100100",
9370 => "10100100",
9371 => "10100100",
9372 => "10100100",
9373 => "10100100",
9374 => "10100100",
9375 => "10100100",
9376 => "10101100",
9377 => "10101101",
9378 => "10101101",
9379 => "10101101",
9380 => "10101101",
9381 => "10101101",
9382 => "10101101",
9383 => "10101100",
9384 => "10101100",
9385 => "10101100",
9386 => "10100100",
9387 => "10100100",
9388 => "10100100",
9389 => "10100100",
9390 => "01011011",
9391 => "01011011",
9392 => "01011011",
9393 => "01011010",
9394 => "01011010",
9395 => "01011010",
9396 => "01011010",
9397 => "01100010",
9398 => "01100010",
9399 => "01100010",
9400 => "01100010",
9401 => "01100010",
9402 => "01011010",
9403 => "01011010",
9404 => "01011010",
9405 => "01011010",
9406 => "01011010",
9407 => "01011011",
9408 => "01011011",
9409 => "10100011",
9410 => "10100100",
9411 => "10100100",
9412 => "10100100",
9413 => "10101100",
9414 => "10101101",
9415 => "10101101",
9416 => "10101101",
9417 => "10101101",
9418 => "10101101",
9419 => "10101101",
9420 => "10101101",
9421 => "10101101",
9422 => "10101101",
9423 => "10101101",
9424 => "10101101",
9425 => "10101101",
9426 => "10101101",
9427 => "10101101",
9428 => "10101101",
9429 => "10101100",
9430 => "10100100",
9431 => "10100100",
9432 => "10100100",
9433 => "10100100",
9434 => "10100100",
9435 => "10100100",
9436 => "10100100",
9437 => "01011011",
9438 => "01010010",
9439 => "01011011",
9440 => "10100011",
9441 => "10100100",
9442 => "10101101",
9443 => "10101101",
9444 => "10101101",
9445 => "10101101",
9446 => "10101101",
9447 => "10101101",
9448 => "10100100",
9449 => "01011011",
9450 => "01011011",
9451 => "01011011",
9452 => "01011011",
9453 => "10100100",
9454 => "10100100",
9455 => "10100100",
9456 => "10100100",
9457 => "10100100",
9458 => "10100100",
9459 => "10101100",
9460 => "10101101",
9472 => "10011011",
9473 => "01011011",
9474 => "01011011",
9475 => "10100011",
9476 => "10011011",
9477 => "10011011",
9478 => "10100011",
9479 => "10100011",
9480 => "10100100",
9481 => "10100100",
9482 => "10100100",
9483 => "10100100",
9484 => "10100100",
9485 => "10100100",
9486 => "10100100",
9487 => "10100100",
9488 => "10100100",
9489 => "10100100",
9490 => "10100100",
9491 => "10100100",
9492 => "10100100",
9493 => "10100100",
9494 => "10100100",
9495 => "10100100",
9496 => "10100100",
9497 => "10100100",
9498 => "10100100",
9499 => "10100100",
9500 => "10100100",
9501 => "10101100",
9502 => "10101100",
9503 => "10101100",
9504 => "10101101",
9505 => "10101101",
9506 => "10101101",
9507 => "10101101",
9508 => "10101101",
9509 => "10101101",
9510 => "10101101",
9511 => "10101101",
9512 => "10101101",
9513 => "10101101",
9514 => "10101101",
9515 => "10101101",
9516 => "10100100",
9517 => "10100100",
9518 => "10100100",
9519 => "10100100",
9520 => "10100100",
9521 => "01100011",
9522 => "01100011",
9523 => "01011011",
9524 => "01011011",
9525 => "01011011",
9526 => "01011010",
9527 => "01011010",
9528 => "01011010",
9529 => "01011010",
9530 => "01011011",
9531 => "01011011",
9532 => "01011011",
9533 => "01100011",
9534 => "10100100",
9535 => "10100100",
9536 => "10100100",
9537 => "10100100",
9538 => "10100100",
9539 => "10101100",
9540 => "10101101",
9541 => "10101101",
9542 => "10101101",
9543 => "10101101",
9544 => "10101101",
9545 => "10101101",
9546 => "10101101",
9547 => "10101101",
9548 => "10101101",
9549 => "10101101",
9550 => "10101101",
9551 => "10101101",
9552 => "10101101",
9553 => "10101101",
9554 => "10101101",
9555 => "10101101",
9556 => "10101101",
9557 => "10101101",
9558 => "10101101",
9559 => "10101101",
9560 => "10101101",
9561 => "10101101",
9562 => "10101100",
9563 => "10100100",
9564 => "10100100",
9565 => "10100100",
9566 => "10100100",
9567 => "10100100",
9568 => "01011011",
9569 => "01011011",
9570 => "01011011",
9571 => "01011011",
9572 => "01011011",
9573 => "01011011",
9574 => "01011011",
9575 => "01011011",
9576 => "01011011",
9577 => "10100100",
9578 => "10100100",
9579 => "10100100",
9580 => "10100100",
9581 => "10100100",
9582 => "10100100",
9583 => "10101101",
9584 => "10101101",
9585 => "10101101",
9586 => "10101101",
9587 => "10101101",
9588 => "10101101",
9600 => "10100100",
9601 => "10100100",
9602 => "10100100",
9603 => "10100100",
9604 => "10100100",
9605 => "10100100",
9606 => "10101100",
9607 => "10101101",
9608 => "10101100",
9609 => "10101100",
9610 => "10100100",
9611 => "10100100",
9612 => "10100100",
9613 => "10100100",
9614 => "10100100",
9615 => "10100100",
9616 => "10100100",
9617 => "10100100",
9618 => "10100100",
9619 => "10100100",
9620 => "10101100",
9621 => "10101100",
9622 => "10101100",
9623 => "10101101",
9624 => "10101101",
9625 => "10101100",
9626 => "10101100",
9627 => "10100100",
9628 => "10100100",
9629 => "10101100",
9630 => "10101100",
9631 => "10101100",
9632 => "10101101",
9633 => "10101101",
9634 => "10101101",
9635 => "10101101",
9636 => "10101101",
9637 => "10101101",
9638 => "10101101",
9639 => "10101101",
9640 => "10101101",
9641 => "10101101",
9642 => "10101101",
9643 => "10101101",
9644 => "10101100",
9645 => "10101100",
9646 => "10101100",
9647 => "10100100",
9648 => "10101100",
9649 => "10101100",
9650 => "10101100",
9651 => "10101100",
9652 => "10101100",
9653 => "10101100",
9654 => "10101100",
9655 => "10101100",
9656 => "10101100",
9657 => "10101100",
9658 => "10101100",
9659 => "10101100",
9660 => "10101100",
9661 => "10101100",
9662 => "10101100",
9663 => "10100100",
9664 => "10101100",
9665 => "10101100",
9666 => "10101100",
9667 => "10101101",
9668 => "10101101",
9669 => "10101101",
9670 => "10101101",
9671 => "10101101",
9672 => "10101101",
9673 => "10101101",
9674 => "10101101",
9675 => "10101101",
9676 => "10101101",
9677 => "10101101",
9678 => "10101101",
9679 => "10101101",
9680 => "10101101",
9681 => "10101101",
9682 => "10101101",
9683 => "10101101",
9684 => "10101101",
9685 => "10101101",
9686 => "10101101",
9687 => "10101101",
9688 => "10101101",
9689 => "10101101",
9690 => "10101101",
9691 => "10101101",
9692 => "10101101",
9693 => "10101101",
9694 => "10101101",
9695 => "10101101",
9696 => "10101101",
9697 => "10101101",
9698 => "10101101",
9699 => "10101101",
9700 => "10101101",
9701 => "10101101",
9702 => "10101101",
9703 => "10101101",
9704 => "10101101",
9705 => "10101101",
9706 => "10101101",
9707 => "10101101",
9708 => "10101101",
9709 => "10101101",
9710 => "10101101",
9711 => "10101101",
9712 => "10101101",
9713 => "10101101",
9714 => "10101101",
9715 => "10101101",
9716 => "10101101",
9728 => "10101101",
9729 => "10101101",
9730 => "10101101",
9731 => "10101101",
9732 => "10101101",
9733 => "10101101",
9734 => "10101101",
9735 => "10101101",
9736 => "10101101",
9737 => "10101101",
9738 => "10101101",
9739 => "10101101",
9740 => "10101101",
9741 => "10101101",
9742 => "10101101",
9743 => "10101101",
9744 => "10101101",
9745 => "10101101",
9746 => "10101101",
9747 => "10101101",
9748 => "10101101",
9749 => "10101101",
9750 => "10101101",
9751 => "10101101",
9752 => "10101101",
9753 => "10101101",
9754 => "10101101",
9755 => "10101101",
9756 => "10101101",
9757 => "10101101",
9758 => "10101101",
9759 => "10101101",
9760 => "10101101",
9761 => "10101101",
9762 => "10101101",
9763 => "10101101",
9764 => "10101101",
9765 => "10101101",
9766 => "10101101",
9767 => "10101101",
9768 => "10101101",
9769 => "10101101",
9770 => "10101101",
9771 => "10101100",
9772 => "10101100",
9773 => "10101100",
9774 => "10101100",
9775 => "10101100",
9776 => "10101100",
9777 => "10101100",
9778 => "10101100",
9779 => "10101100",
9780 => "10101100",
9781 => "10101100",
9782 => "10101100",
9783 => "10101100",
9784 => "10101100",
9785 => "10101100",
9786 => "10101100",
9787 => "10101100",
9788 => "10101100",
9789 => "10101100",
9790 => "10101100",
9791 => "10101100",
9792 => "10101100",
9793 => "10101100",
9794 => "10101100",
9795 => "10101100",
9796 => "10101101",
9797 => "10101101",
9798 => "10101101",
9799 => "10101101",
9800 => "10101101",
9801 => "10101101",
9802 => "10101101",
9803 => "10101101",
9804 => "10101101",
9805 => "10101101",
9806 => "10101101",
9807 => "10101101",
9808 => "10101101",
9809 => "10101101",
9810 => "10101101",
9811 => "10101101",
9812 => "10101101",
9813 => "10101101",
9814 => "10101101",
9815 => "10101101",
9816 => "10101101",
9817 => "10101101",
9818 => "10101101",
9819 => "10101101",
9820 => "10101101",
9821 => "10101101",
9822 => "10101101",
9823 => "10101101",
9824 => "10101101",
9825 => "10101100",
9826 => "10101100",
9827 => "10101100",
9828 => "10101100",
9829 => "10101100",
9830 => "10101100",
9831 => "10101100",
9832 => "10101100",
9833 => "10101101",
9834 => "10101101",
9835 => "10101101",
9836 => "10101101",
9837 => "10101101",
9838 => "10101101",
9839 => "10101101",
9840 => "10101101",
9841 => "10101101",
9842 => "10101101",
9843 => "10101101",
9844 => "10101101",
9856 => "10101101",
9857 => "10101101",
9858 => "10101101",
9859 => "10101101",
9860 => "10101101",
9861 => "10101101",
9862 => "10101101",
9863 => "10101101",
9864 => "10101101",
9865 => "10101101",
9866 => "10101101",
9867 => "10101101",
9868 => "10101101",
9869 => "10101101",
9870 => "10101101",
9871 => "10101101",
9872 => "10101101",
9873 => "10101101",
9874 => "10101101",
9875 => "10101101",
9876 => "10101101",
9877 => "10101101",
9878 => "10101101",
9879 => "10101101",
9880 => "10101101",
9881 => "10101101",
9882 => "10101101",
9883 => "10101101",
9884 => "10101101",
9885 => "10101101",
9886 => "10101101",
9887 => "10101101",
9888 => "10101101",
9889 => "10101101",
9890 => "10101101",
9891 => "10101101",
9892 => "10101101",
9893 => "10101101",
9894 => "10101101",
9895 => "10101101",
9896 => "10101101",
9897 => "10101101",
9898 => "10101101",
9899 => "10101101",
9900 => "10101100",
9901 => "10101100",
9902 => "10101100",
9903 => "10101100",
9904 => "10101100",
9905 => "10101100",
9906 => "10101100",
9907 => "10101100",
9908 => "10101100",
9909 => "10101100",
9910 => "10101100",
9911 => "10101100",
9912 => "10101100",
9913 => "10101100",
9914 => "10101100",
9915 => "10101100",
9916 => "10101100",
9917 => "10101100",
9918 => "10101100",
9919 => "10101100",
9920 => "10101100",
9921 => "10101100",
9922 => "10101100",
9923 => "10101101",
9924 => "10101101",
9925 => "10101101",
9926 => "10101101",
9927 => "10101101",
9928 => "10101101",
9929 => "10101101",
9930 => "10101101",
9931 => "10101101",
9932 => "10101101",
9933 => "10101101",
9934 => "10101101",
9935 => "10101101",
9936 => "10101101",
9937 => "10101101",
9938 => "10101101",
9939 => "10101101",
9940 => "10101101",
9941 => "10101101",
9942 => "10101101",
9943 => "10101101",
9944 => "10101101",
9945 => "10101101",
9946 => "10101101",
9947 => "10101101",
9948 => "10101101",
9949 => "10101100",
9950 => "10101100",
9951 => "10101100",
9952 => "10101100",
9953 => "10101100",
9954 => "10101100",
9955 => "10101100",
9956 => "10101100",
9957 => "10101100",
9958 => "10101100",
9959 => "10101100",
9960 => "10101100",
9961 => "10101100",
9962 => "10101100",
9963 => "10101100",
9964 => "10101101",
9965 => "10101101",
9966 => "10101101",
9967 => "10101101",
9968 => "10101101",
9969 => "10101101",
9970 => "10101101",
9971 => "10101101",
9972 => "10101101",
9984 => "10110101",
9985 => "10110101",
9986 => "10110101",
9987 => "10110101",
9988 => "10110101",
9989 => "10110101",
9990 => "10110101",
9991 => "10110101",
9992 => "10110110",
9993 => "10110110",
9994 => "10110101",
9995 => "10110110",
9996 => "10110101",
9997 => "10110101",
9998 => "10110101",
9999 => "10101101",
10000 => "10101101",
10001 => "10101101",
10002 => "10101101",
10003 => "10101101",
10004 => "10101101",
10005 => "10101101",
10006 => "10101101",
10007 => "10101101",
10008 => "10101101",
10009 => "10101101",
10010 => "10101101",
10011 => "10101101",
10012 => "10101101",
10013 => "10101101",
10014 => "10101101",
10015 => "10101101",
10016 => "10101101",
10017 => "10101101",
10018 => "10101101",
10019 => "10101101",
10020 => "10101101",
10021 => "10101101",
10022 => "10101101",
10023 => "10101101",
10024 => "10101101",
10025 => "10101101",
10026 => "10101101",
10027 => "10101101",
10028 => "10101101",
10029 => "10101100",
10030 => "10101100",
10031 => "10101100",
10032 => "10101100",
10033 => "10101100",
10034 => "10101100",
10035 => "10101100",
10036 => "10101100",
10037 => "10101101",
10038 => "10101101",
10039 => "10101101",
10040 => "10101101",
10041 => "10101101",
10042 => "10101101",
10043 => "10101100",
10044 => "10101100",
10045 => "10101100",
10046 => "10101100",
10047 => "10101100",
10048 => "10101100",
10049 => "10101100",
10050 => "10101101",
10051 => "10101101",
10052 => "10101101",
10053 => "10101101",
10054 => "10101101",
10055 => "10101101",
10056 => "10101101",
10057 => "10101101",
10058 => "10101101",
10059 => "10101101",
10060 => "10101101",
10061 => "10101101",
10062 => "10101101",
10063 => "10101101",
10064 => "10101101",
10065 => "10101101",
10066 => "10101101",
10067 => "10101101",
10068 => "10101101",
10069 => "10101101",
10070 => "10101101",
10071 => "10101101",
10072 => "10101101",
10073 => "10101101",
10074 => "10101101",
10075 => "10101100",
10076 => "10101100",
10077 => "10101100",
10078 => "10101100",
10079 => "10101100",
10080 => "10101100",
10081 => "10101011",
10082 => "10101011",
10083 => "10101011",
10084 => "10101011",
10085 => "10101011",
10086 => "10101011",
10087 => "10101011",
10088 => "10101100",
10089 => "10101100",
10090 => "10101100",
10091 => "10101100",
10092 => "10101100",
10093 => "10101100",
10094 => "10101101",
10095 => "10101101",
10096 => "10101101",
10097 => "10101101",
10098 => "10101101",
10099 => "10101101",
10100 => "10101101",
10112 => "10110101",
10113 => "10101101",
10114 => "10101101",
10115 => "10101101",
10116 => "10101101",
10117 => "10101101",
10118 => "10110101",
10119 => "10110101",
10120 => "10110101",
10121 => "10110101",
10122 => "10110101",
10123 => "10110101",
10124 => "10110110",
10125 => "10110110",
10126 => "10110110",
10127 => "10110110",
10128 => "10110110",
10129 => "10110101",
10130 => "10110101",
10131 => "10110101",
10132 => "10110101",
10133 => "10101101",
10134 => "10101101",
10135 => "10101101",
10136 => "10101101",
10137 => "10101101",
10138 => "10101101",
10139 => "10101101",
10140 => "10101101",
10141 => "10101101",
10142 => "10101101",
10143 => "10101101",
10144 => "10101101",
10145 => "10101101",
10146 => "10101101",
10147 => "10101101",
10148 => "10101101",
10149 => "10101101",
10150 => "10101101",
10151 => "10101101",
10152 => "10101101",
10153 => "10101101",
10154 => "10101101",
10155 => "10101101",
10156 => "10101101",
10157 => "10101100",
10158 => "10101100",
10159 => "10101100",
10160 => "10101100",
10161 => "10101100",
10162 => "10101100",
10163 => "10101100",
10164 => "10101100",
10165 => "10101100",
10166 => "10101101",
10167 => "10101101",
10168 => "10101101",
10169 => "10101101",
10170 => "10101101",
10171 => "10101101",
10172 => "10101100",
10173 => "10101100",
10174 => "10101100",
10175 => "10101100",
10176 => "10101100",
10177 => "10101100",
10178 => "10101101",
10179 => "10101101",
10180 => "10101101",
10181 => "10101101",
10182 => "10101101",
10183 => "10101101",
10184 => "10101101",
10185 => "10101101",
10186 => "10101101",
10187 => "10101101",
10188 => "10101101",
10189 => "10101101",
10190 => "10101101",
10191 => "10101101",
10192 => "10101101",
10193 => "10101101",
10194 => "10101101",
10195 => "10101101",
10196 => "10101101",
10197 => "10101101",
10198 => "10101101",
10199 => "10101101",
10200 => "10101101",
10201 => "10101101",
10202 => "10101100",
10203 => "10101100",
10204 => "10101100",
10205 => "10101100",
10206 => "10101011",
10207 => "10101011",
10208 => "10101011",
10209 => "10101011",
10210 => "10101011",
10211 => "10101011",
10212 => "10101011",
10213 => "10101011",
10214 => "10101011",
10215 => "10101011",
10216 => "10101011",
10217 => "10101011",
10218 => "10101011",
10219 => "10101100",
10220 => "10101100",
10221 => "10101100",
10222 => "10101100",
10223 => "10101101",
10224 => "10101101",
10225 => "10101101",
10226 => "10101101",
10227 => "10101101",
10228 => "10101101",
10240 => "10101101",
10241 => "10101101",
10242 => "10101101",
10243 => "10101101",
10244 => "10101101",
10245 => "10101101",
10246 => "10101101",
10247 => "10101101",
10248 => "10101101",
10249 => "10101101",
10250 => "10110101",
10251 => "10110101",
10252 => "10110101",
10253 => "10110101",
10254 => "10110101",
10255 => "10110101",
10256 => "10110110",
10257 => "10110110",
10258 => "10110110",
10259 => "10110110",
10260 => "10110110",
10261 => "10110110",
10262 => "10110110",
10263 => "10110110",
10264 => "10110110",
10265 => "10110101",
10266 => "10101101",
10267 => "10101101",
10268 => "10101101",
10269 => "10101101",
10270 => "10101101",
10271 => "10101101",
10272 => "10101101",
10273 => "10101101",
10274 => "10101101",
10275 => "10101101",
10276 => "10101101",
10277 => "10101101",
10278 => "10101101",
10279 => "10101101",
10280 => "10101101",
10281 => "10101101",
10282 => "10101101",
10283 => "10101101",
10284 => "10101101",
10285 => "10101101",
10286 => "10101100",
10287 => "10101100",
10288 => "10101100",
10289 => "10101100",
10290 => "10101100",
10291 => "10101100",
10292 => "10101101",
10293 => "10101101",
10294 => "10101101",
10295 => "10110101",
10296 => "10110101",
10297 => "10110101",
10298 => "10110101",
10299 => "10101101",
10300 => "10101101",
10301 => "10101100",
10302 => "10101100",
10303 => "10101100",
10304 => "10101100",
10305 => "10101101",
10306 => "10101101",
10307 => "10101101",
10308 => "10101101",
10309 => "10101101",
10310 => "10101101",
10311 => "10101101",
10312 => "10101101",
10313 => "10101101",
10314 => "10101101",
10315 => "10101101",
10316 => "10101101",
10317 => "10101101",
10318 => "10101101",
10319 => "10101101",
10320 => "10101101",
10321 => "10101101",
10322 => "10101101",
10323 => "10101101",
10324 => "10101101",
10325 => "10101101",
10326 => "10101101",
10327 => "10101101",
10328 => "10101101",
10329 => "10101100",
10330 => "10101100",
10331 => "10101100",
10332 => "10101100",
10333 => "10101011",
10334 => "10101011",
10335 => "10101011",
10336 => "10101011",
10337 => "10101011",
10338 => "10101011",
10339 => "10101011",
10340 => "10101011",
10341 => "10101011",
10342 => "10101011",
10343 => "10101011",
10344 => "10101011",
10345 => "10101011",
10346 => "10101011",
10347 => "10101011",
10348 => "10101100",
10349 => "10101100",
10350 => "10101100",
10351 => "10101100",
10352 => "10101100",
10353 => "10101101",
10354 => "10101101",
10355 => "10101101",
10356 => "10101101",
10368 => "10101101",
10369 => "10101101",
10370 => "10101101",
10371 => "10101101",
10372 => "10101101",
10373 => "10101101",
10374 => "10101101",
10375 => "10101101",
10376 => "10101101",
10377 => "10101101",
10378 => "10101101",
10379 => "10101101",
10380 => "10101101",
10381 => "10101101",
10382 => "10110101",
10383 => "10110101",
10384 => "10110101",
10385 => "10110101",
10386 => "10110101",
10387 => "10110101",
10388 => "10110110",
10389 => "10110110",
10390 => "10110110",
10391 => "10110110",
10392 => "10110110",
10393 => "10110110",
10394 => "10110101",
10395 => "10101101",
10396 => "10101101",
10397 => "10101101",
10398 => "10101101",
10399 => "10101101",
10400 => "10101101",
10401 => "10101101",
10402 => "10101101",
10403 => "10101101",
10404 => "10101101",
10405 => "10101101",
10406 => "10101101",
10407 => "10101101",
10408 => "10101101",
10409 => "10101101",
10410 => "10101101",
10411 => "10101101",
10412 => "10101101",
10413 => "10101101",
10414 => "10101100",
10415 => "10101100",
10416 => "10101100",
10417 => "10101100",
10418 => "10101100",
10419 => "10101101",
10420 => "10101101",
10421 => "10101101",
10422 => "10110101",
10423 => "10101101",
10424 => "10110101",
10425 => "10110101",
10426 => "10110101",
10427 => "10101101",
10428 => "10101101",
10429 => "10101100",
10430 => "10101100",
10431 => "10101100",
10432 => "10101100",
10433 => "10101101",
10434 => "10101101",
10435 => "10101101",
10436 => "10101101",
10437 => "10101101",
10438 => "10101101",
10439 => "10101101",
10440 => "10101101",
10441 => "10101101",
10442 => "10101101",
10443 => "10101101",
10444 => "10101101",
10445 => "10101101",
10446 => "10101101",
10447 => "10101101",
10448 => "10101101",
10449 => "10101101",
10450 => "10101101",
10451 => "10101101",
10452 => "10101101",
10453 => "10101101",
10454 => "10101101",
10455 => "10101100",
10456 => "10101100",
10457 => "10101100",
10458 => "10101100",
10459 => "10101100",
10460 => "10101011",
10461 => "10101011",
10462 => "10101011",
10463 => "10101011",
10464 => "10101011",
10465 => "10101011",
10466 => "10101011",
10467 => "10101011",
10468 => "10101011",
10469 => "10101011",
10470 => "10101011",
10471 => "10101011",
10472 => "10101011",
10473 => "10101011",
10474 => "10101011",
10475 => "10101011",
10476 => "10101011",
10477 => "10101011",
10478 => "10101100",
10479 => "10101100",
10480 => "10101100",
10481 => "10101100",
10482 => "10101101",
10483 => "10101101",
10484 => "10101101",
10496 => "10101101",
10497 => "10101101",
10498 => "10101101",
10499 => "10101101",
10500 => "10101101",
10501 => "10101101",
10502 => "10101101",
10503 => "10101101",
10504 => "10101101",
10505 => "10101101",
10506 => "10101101",
10507 => "10101101",
10508 => "10101101",
10509 => "10101101",
10510 => "10101101",
10511 => "10101101",
10512 => "10101101",
10513 => "10101101",
10514 => "10101101",
10515 => "10101101",
10516 => "10110101",
10517 => "10110101",
10518 => "10110101",
10519 => "10110110",
10520 => "10110110",
10521 => "10110110",
10522 => "10110110",
10523 => "10110110",
10524 => "10101101",
10525 => "10101101",
10526 => "10101101",
10527 => "10101101",
10528 => "10101101",
10529 => "10101101",
10530 => "10101101",
10531 => "10101101",
10532 => "10101101",
10533 => "10101101",
10534 => "10101101",
10535 => "10101101",
10536 => "10101101",
10537 => "10101101",
10538 => "10101101",
10539 => "10101101",
10540 => "10101101",
10541 => "10101101",
10542 => "10101101",
10543 => "10101101",
10544 => "10101101",
10545 => "10101101",
10546 => "10101101",
10547 => "10101101",
10548 => "10110101",
10549 => "10110101",
10550 => "10110101",
10551 => "10110101",
10552 => "10110101",
10553 => "10110101",
10554 => "10110101",
10555 => "10110101",
10556 => "10110101",
10557 => "10110101",
10558 => "10101101",
10559 => "10101101",
10560 => "10101101",
10561 => "10101101",
10562 => "10101101",
10563 => "10101101",
10564 => "10101101",
10565 => "10101101",
10566 => "10101101",
10567 => "10101101",
10568 => "10101101",
10569 => "10101101",
10570 => "10101101",
10571 => "10101101",
10572 => "10101101",
10573 => "10101101",
10574 => "10101101",
10575 => "10101101",
10576 => "10101101",
10577 => "10101101",
10578 => "10101101",
10579 => "10101101",
10580 => "10101101",
10581 => "10101101",
10582 => "10101101",
10583 => "10101100",
10584 => "10101100",
10585 => "10101100",
10586 => "10101100",
10587 => "10101100",
10588 => "10101100",
10589 => "10101100",
10590 => "10101100",
10591 => "10101100",
10592 => "10101100",
10593 => "10101100",
10594 => "10101100",
10595 => "10101100",
10596 => "10101100",
10597 => "10101100",
10598 => "10101100",
10599 => "10101100",
10600 => "10101100",
10601 => "10101100",
10602 => "10101100",
10603 => "10101100",
10604 => "10101100",
10605 => "10101100",
10606 => "10101100",
10607 => "10101100",
10608 => "10101100",
10609 => "10101100",
10610 => "10101101",
10611 => "10101101",
10612 => "10101101",
10624 => "10101101",
10625 => "10101101",
10626 => "10101101",
10627 => "10101101",
10628 => "10101101",
10629 => "10101101",
10630 => "10101101",
10631 => "10101101",
10632 => "10101101",
10633 => "10101101",
10634 => "10101101",
10635 => "10101101",
10636 => "10101101",
10637 => "10101101",
10638 => "10101101",
10639 => "10101101",
10640 => "10101101",
10641 => "10101101",
10642 => "10101101",
10643 => "10101101",
10644 => "10101101",
10645 => "10101101",
10646 => "10110101",
10647 => "10110101",
10648 => "10110101",
10649 => "10110110",
10650 => "10110110",
10651 => "10110101",
10652 => "10110101",
10653 => "10101101",
10654 => "10101101",
10655 => "10101101",
10656 => "10101101",
10657 => "10101101",
10658 => "10101101",
10659 => "10101101",
10660 => "10101101",
10661 => "10101101",
10662 => "10101101",
10663 => "10101101",
10664 => "10101101",
10665 => "10101101",
10666 => "10101101",
10667 => "10101101",
10668 => "10101101",
10669 => "10101101",
10670 => "10101101",
10671 => "10101101",
10672 => "10101101",
10673 => "10101101",
10674 => "10110101",
10675 => "10110101",
10676 => "10110101",
10677 => "10110101",
10678 => "10110101",
10679 => "10110101",
10680 => "10110101",
10681 => "10110101",
10682 => "10110101",
10683 => "10110101",
10684 => "10110101",
10685 => "10110101",
10686 => "10101101",
10687 => "10101101",
10688 => "10101101",
10689 => "10101101",
10690 => "10101101",
10691 => "10101101",
10692 => "10101101",
10693 => "10101101",
10694 => "10101101",
10695 => "10101101",
10696 => "10101101",
10697 => "10101101",
10698 => "10101101",
10699 => "10101101",
10700 => "10101101",
10701 => "10101101",
10702 => "10101101",
10703 => "10101101",
10704 => "10101101",
10705 => "10101101",
10706 => "10101101",
10707 => "10101101",
10708 => "10101101",
10709 => "10101101",
10710 => "10101101",
10711 => "10101100",
10712 => "10101100",
10713 => "10101100",
10714 => "10101100",
10715 => "10101100",
10716 => "10101100",
10717 => "10101100",
10718 => "10101100",
10719 => "10101100",
10720 => "10101100",
10721 => "10101100",
10722 => "10101100",
10723 => "10110100",
10724 => "10110100",
10725 => "10101100",
10726 => "10101100",
10727 => "10101100",
10728 => "10101100",
10729 => "10101100",
10730 => "10101100",
10731 => "10101100",
10732 => "10101100",
10733 => "10101100",
10734 => "10101100",
10735 => "10101100",
10736 => "10101100",
10737 => "10101100",
10738 => "10101100",
10739 => "10101101",
10740 => "10101101",
10752 => "11111110",
10753 => "11111110",
10754 => "11111110",
10755 => "11111110",
10756 => "11111110",
10757 => "11111110",
10758 => "11111110",
10759 => "11111110",
10760 => "11111110",
10761 => "11110110",
10762 => "11110110",
10763 => "11110110",
10764 => "11110110",
10765 => "11110110",
10766 => "11110110",
10767 => "11110110",
10768 => "11110110",
10769 => "11110110",
10770 => "11110110",
10771 => "11110110",
10772 => "11110110",
10773 => "11110110",
10774 => "11111110",
10775 => "11111111",
10776 => "11111111",
10777 => "11111111",
10778 => "11111111",
10779 => "11111111",
10780 => "11111111",
10781 => "11111111",
10782 => "11111111",
10783 => "11111111",
10784 => "11111111",
10785 => "11111111",
10786 => "11111111",
10787 => "11111111",
10788 => "11111111",
10789 => "11111111",
10790 => "11111111",
10791 => "11111111",
10792 => "11111111",
10793 => "11111111",
10794 => "11111111",
10795 => "11111110",
10796 => "11111110",
10797 => "11111110",
10798 => "11111110",
10799 => "10111110",
10800 => "10111110",
10801 => "10111110",
10802 => "10111110",
10803 => "10111110",
10804 => "10111110",
10805 => "10111110",
10806 => "10111110",
10807 => "10111110",
10808 => "10111110",
10809 => "10111110",
10810 => "10111110",
10811 => "10111110",
10812 => "10111110",
10813 => "10111110",
10814 => "10111110",
10815 => "10111110",
10816 => "11111110",
10817 => "11111110",
10818 => "11111110",
10819 => "11111110",
10820 => "11111111",
10821 => "11111111",
10822 => "11111111",
10823 => "11111111",
10824 => "11111111",
10825 => "11111111",
10826 => "11111111",
10827 => "11111111",
10828 => "11111111",
10829 => "11111111",
10830 => "11111111",
10831 => "11111111",
10832 => "11111111",
10833 => "11111111",
10834 => "11111111",
10835 => "11111110",
10836 => "11110110",
10837 => "11110110",
10838 => "11110110",
10839 => "11110110",
10840 => "11110110",
10841 => "11110110",
10842 => "11110110",
10843 => "11110110",
10844 => "11110110",
10845 => "11111110",
10846 => "11111110",
10847 => "11111110",
10848 => "11111110",
10849 => "11111110",
10850 => "11111110",
10851 => "11111101",
10852 => "11111101",
10853 => "11111101",
10854 => "11111101",
10855 => "11111101",
10856 => "11111101",
10857 => "11111101",
10858 => "11110101",
10859 => "11110101",
10860 => "11110101",
10861 => "11110101",
10862 => "11110101",
10863 => "11110101",
10864 => "11110101",
10865 => "11110101",
10866 => "11110110",
10867 => "11110110",
10868 => "11110110",
10880 => "10100100",
10881 => "10100100",
10882 => "10100100",
10883 => "10100100",
10884 => "10100100",
10885 => "10100100",
10886 => "10100100",
10887 => "10100100",
10888 => "10100100",
10889 => "10100100",
10890 => "10100100",
10891 => "10100100",
10892 => "10100100",
10893 => "10100100",
10894 => "10100100",
10895 => "10100100",
10896 => "10100100",
10897 => "10100100",
10898 => "10100100",
10899 => "10100100",
10900 => "10100100",
10901 => "10100100",
10902 => "10100100",
10903 => "10100100",
10904 => "10100100",
10905 => "10100100",
10906 => "10100100",
10907 => "10100100",
10908 => "10100100",
10909 => "10100100",
10910 => "10100100",
10911 => "10100100",
10912 => "10100100",
10913 => "10100100",
10914 => "10100100",
10915 => "10100100",
10916 => "10100100",
10917 => "10100100",
10918 => "10100100",
10919 => "10100100",
10920 => "10100100",
10921 => "10100100",
10922 => "10100100",
10923 => "10100100",
10924 => "10100100",
10925 => "10100100",
10926 => "10100100",
10927 => "10100100",
10928 => "10100100",
10929 => "10100100",
10930 => "10100100",
10931 => "10100100",
10932 => "10100100",
10933 => "10100100",
10934 => "10100100",
10935 => "10100100",
10936 => "10100100",
10937 => "10100100",
10938 => "10100100",
10939 => "10100100",
10940 => "10100100",
10941 => "10100100",
10942 => "10100100",
10943 => "10100100",
10944 => "10100100",
10945 => "10100100",
10946 => "10100100",
10947 => "10100100",
10948 => "10100100",
10949 => "10100100",
10950 => "10100100",
10951 => "10100100",
10952 => "10100100",
10953 => "10100100",
10954 => "10100100",
10955 => "10100100",
10956 => "10100100",
10957 => "10100100",
10958 => "10100100",
10959 => "10100100",
10960 => "10100100",
10961 => "10100100",
10962 => "10100100",
10963 => "10100100",
10964 => "10100100",
10965 => "10100100",
10966 => "10100100",
10967 => "10100100",
10968 => "10100100",
10969 => "10100100",
10970 => "10100100",
10971 => "10100100",
10972 => "10100100",
10973 => "10100100",
10974 => "10100100",
10975 => "10100100",
10976 => "10100100",
10977 => "10100100",
10978 => "10100100",
10979 => "10100100",
10980 => "10100100",
10981 => "10100100",
10982 => "10100100",
10983 => "10100100",
10984 => "10100100",
10985 => "10100100",
10986 => "10100100",
10987 => "10100100",
10988 => "10100100",
10989 => "10100100",
10990 => "10100100",
10991 => "10100100",
10992 => "10100100",
10993 => "10100100",
10994 => "10100100",
10995 => "10100100",
10996 => "10100100",
11008 => "10100100",
11009 => "10100100",
11010 => "10100100",
11011 => "10100100",
11012 => "10100100",
11013 => "10100100",
11014 => "10100100",
11015 => "10100100",
11016 => "10100100",
11017 => "10100100",
11018 => "10100100",
11019 => "10100100",
11020 => "10100100",
11021 => "10100100",
11022 => "10100100",
11023 => "10100100",
11024 => "10100100",
11025 => "10100100",
11026 => "10100100",
11027 => "10100100",
11028 => "10100100",
11029 => "10100100",
11030 => "10100100",
11031 => "10100100",
11032 => "10100100",
11033 => "10100100",
11034 => "10100100",
11035 => "10100100",
11036 => "10100100",
11037 => "10100100",
11038 => "10100100",
11039 => "10100100",
11040 => "10100100",
11041 => "10100100",
11042 => "10100100",
11043 => "10100100",
11044 => "10100100",
11045 => "10100100",
11046 => "10100100",
11047 => "10100100",
11048 => "10100100",
11049 => "10100100",
11050 => "10100100",
11051 => "10100100",
11052 => "10100100",
11053 => "10100100",
11054 => "10100100",
11055 => "10100100",
11056 => "10100100",
11057 => "10100100",
11058 => "10100100",
11059 => "10100100",
11060 => "10100100",
11061 => "10100100",
11062 => "10100100",
11063 => "10100100",
11064 => "10100100",
11065 => "10100100",
11066 => "10100100",
11067 => "10100100",
11068 => "10100100",
11069 => "10100100",
11070 => "10100100",
11071 => "10100100",
11072 => "10100100",
11073 => "10100100",
11074 => "10100100",
11075 => "10100100",
11076 => "10100100",
11077 => "10100100",
11078 => "10100100",
11079 => "10100100",
11080 => "10100100",
11081 => "10100100",
11082 => "10100100",
11083 => "10100100",
11084 => "10100100",
11085 => "10100100",
11086 => "10100100",
11087 => "10100100",
11088 => "10100100",
11089 => "10100100",
11090 => "10100100",
11091 => "10100100",
11092 => "10100100",
11093 => "10100100",
11094 => "10100100",
11095 => "10100100",
11096 => "10100100",
11097 => "10100100",
11098 => "10100100",
11099 => "10100100",
11100 => "10100100",
11101 => "10100100",
11102 => "10100100",
11103 => "10100100",
11104 => "10100100",
11105 => "10100100",
11106 => "10100100",
11107 => "10100100",
11108 => "10100100",
11109 => "10100100",
11110 => "10100100",
11111 => "10100100",
11112 => "10100100",
11113 => "10100100",
11114 => "10100100",
11115 => "10100100",
11116 => "10100100",
11117 => "10100100",
11118 => "10100100",
11119 => "10100100",
11120 => "10100100",
11121 => "10100100",
11122 => "10100100",
11123 => "10100100",
11124 => "10100100",
11136 => "10100100",
11137 => "10100100",
11138 => "10100100",
11139 => "10100100",
11140 => "10100100",
11141 => "10100100",
11142 => "10100100",
11143 => "10100100",
11144 => "10100100",
11145 => "10100100",
11146 => "10100100",
11147 => "10100100",
11148 => "10100100",
11149 => "10100100",
11150 => "10100100",
11151 => "10100100",
11152 => "10100100",
11153 => "10100100",
11154 => "10100100",
11155 => "10100100",
11156 => "10100100",
11157 => "10100100",
11158 => "10100100",
11159 => "10100100",
11160 => "10100100",
11161 => "10100100",
11162 => "10100100",
11163 => "10100100",
11164 => "10100100",
11165 => "10100100",
11166 => "10100100",
11167 => "10100100",
11168 => "10100100",
11169 => "10100100",
11170 => "10100100",
11171 => "10100100",
11172 => "10100100",
11173 => "10100100",
11174 => "10100100",
11175 => "10100100",
11176 => "10100100",
11177 => "10100100",
11178 => "10100100",
11179 => "10100100",
11180 => "10100100",
11181 => "10100100",
11182 => "10100100",
11183 => "10100100",
11184 => "10100100",
11185 => "10100100",
11186 => "10100100",
11187 => "10100100",
11188 => "10100100",
11189 => "10100100",
11190 => "10100100",
11191 => "10100100",
11192 => "10100100",
11193 => "10100100",
11194 => "10100100",
11195 => "10100100",
11196 => "10100100",
11197 => "10100100",
11198 => "10100100",
11199 => "10100100",
11200 => "10100100",
11201 => "10100100",
11202 => "10100100",
11203 => "10100100",
11204 => "10100100",
11205 => "10100100",
11206 => "10100100",
11207 => "10100100",
11208 => "10100100",
11209 => "10100100",
11210 => "10100100",
11211 => "10100100",
11212 => "10100100",
11213 => "10100100",
11214 => "10100100",
11215 => "10100100",
11216 => "10100100",
11217 => "10100100",
11218 => "10100100",
11219 => "10100100",
11220 => "10100100",
11221 => "10100100",
11222 => "10100100",
11223 => "10100100",
11224 => "10100100",
11225 => "10100100",
11226 => "10100100",
11227 => "10100100",
11228 => "10100100",
11229 => "10100100",
11230 => "10100100",
11231 => "10100100",
11232 => "10100100",
11233 => "10100100",
11234 => "10100100",
11235 => "10100100",
11236 => "10100100",
11237 => "10100100",
11238 => "10100100",
11239 => "10100100",
11240 => "10100100",
11241 => "10100100",
11242 => "10100100",
11243 => "10100100",
11244 => "10100100",
11245 => "10100100",
11246 => "10100100",
11247 => "10100100",
11248 => "10100100",
11249 => "10100100",
11250 => "10100100",
11251 => "10100100",
11252 => "10100100",
