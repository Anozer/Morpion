library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM_vide_sel is
	port (CLK : in std_logic;
		  EN : in std_logic;
		  ADDR : in std_logic_vector(13 downto 0);
		  DATA : out std_logic_vector(7 downto 0));
end ROM_vide_sel;

architecture Behavioral of ROM_vide_sel is

type zone_memoire is array ((2**14)-1 downto 0) of std_logic_vector (7 downto 0);
constant ROM: zone_memoire := (
	0 => "11111111",
	1 => "11111111",
	2 => "11111111",
	3 => "11111111",
	4 => "11111111",
	5 => "11111111",
	6 => "11111111",
	7 => "11111111",
	8 => "11111111",
	9 => "11111111",
	10 => "11111111",
	11 => "11111111",
	12 => "11111111",
	13 => "11111111",
	14 => "11111111",
	15 => "11111111",
	16 => "11111111",
	17 => "11111111",
	18 => "11111111",
	19 => "11111111",
	20 => "11111111",
	21 => "11111111",
	22 => "11111111",
	23 => "11111111",
	24 => "11111111",
	25 => "11111111",
	26 => "11111111",
	27 => "11111111",
	28 => "11111111",
	29 => "11111111",
	30 => "11111111",
	31 => "11111111",
	32 => "11111111",
	33 => "11111111",
	34 => "11111111",
	35 => "11111111",
	36 => "11111111",
	37 => "11111111",
	38 => "11111111",
	39 => "11111111",
	40 => "11111111",
	41 => "11111111",
	42 => "11111111",
	43 => "11111111",
	44 => "11111111",
	45 => "11111111",
	46 => "11111111",
	47 => "11111111",
	48 => "11111111",
	49 => "11111111",
	50 => "11111111",
	51 => "11111111",
	52 => "11111111",
	53 => "11111111",
	54 => "11111111",
	55 => "11111111",
	56 => "11111111",
	57 => "11111111",
	58 => "11111111",
	59 => "11111111",
	60 => "11111111",
	61 => "11111111",
	62 => "11111111",
	63 => "11111111",
	64 => "11111111",
	65 => "11111111",
	66 => "11111111",
	67 => "11111111",
	68 => "11111111",
	69 => "11111111",
	70 => "11111111",
	71 => "11111111",
	72 => "11111111",
	73 => "11111111",
	74 => "11111111",
	75 => "11111111",
	76 => "11111111",
	77 => "11111111",
	78 => "11111111",
	79 => "11111111",
	80 => "11111111",
	81 => "11111111",
	82 => "11111111",
	83 => "11111111",
	84 => "11111111",
	85 => "11111111",
	86 => "11111111",
	87 => "11111111",
	88 => "11111111",
	89 => "11111111",
	90 => "11111111",
	91 => "11111111",
	92 => "11111111",
	93 => "11111111",
	94 => "11111111",
	95 => "11111111",
	96 => "11111111",
	97 => "11111111",
	98 => "11111111",
	99 => "11111111",
	100 => "11111111",
	101 => "11111111",
	102 => "11111111",
	103 => "11111111",
	104 => "11111111",
	105 => "11111111",
	106 => "11111111",
	107 => "11111111",
	108 => "11111111",
	109 => "11111111",
	110 => "11111111",
	111 => "11111111",
	112 => "11111111",
	113 => "11111111",
	114 => "11111111",
	115 => "11111111",
	116 => "11111111",
	117 => "11111111",
	118 => "11111111",
	119 => "11111111",
	128 => "11111111",
	129 => "11111111",
	130 => "11111111",
	131 => "11111111",
	132 => "11111111",
	133 => "11111111",
	134 => "11111111",
	135 => "11111111",
	136 => "11111111",
	137 => "11111111",
	138 => "11111111",
	139 => "11111111",
	140 => "11111111",
	141 => "11111111",
	142 => "11111111",
	143 => "11111111",
	144 => "11111111",
	145 => "11111111",
	146 => "11111111",
	147 => "11111111",
	148 => "11111111",
	149 => "11111111",
	150 => "11111111",
	151 => "11111111",
	152 => "11111111",
	153 => "11111111",
	154 => "11111111",
	155 => "11111111",
	156 => "11111111",
	157 => "11111111",
	158 => "11111111",
	159 => "11111111",
	160 => "11111111",
	161 => "11111111",
	162 => "11111111",
	163 => "11111111",
	164 => "11111111",
	165 => "11111111",
	166 => "11111111",
	167 => "11111111",
	168 => "11111111",
	169 => "11111111",
	170 => "11111111",
	171 => "11111111",
	172 => "11111111",
	173 => "11111111",
	174 => "11111111",
	175 => "11111111",
	176 => "11111111",
	177 => "11111111",
	178 => "11111111",
	179 => "11111111",
	180 => "11111111",
	181 => "11111111",
	182 => "11111111",
	183 => "11111111",
	184 => "11111111",
	185 => "11111111",
	186 => "11111111",
	187 => "11111111",
	188 => "11111111",
	189 => "11111111",
	190 => "11111111",
	191 => "11111111",
	192 => "11111111",
	193 => "11111111",
	194 => "11111111",
	195 => "11111111",
	196 => "11111111",
	197 => "11111111",
	198 => "11111111",
	199 => "11111111",
	200 => "11111111",
	201 => "11111111",
	202 => "11111111",
	203 => "11111111",
	204 => "11111111",
	205 => "11111111",
	206 => "11111111",
	207 => "11111111",
	208 => "11111111",
	209 => "11111111",
	210 => "11111111",
	211 => "11111111",
	212 => "11111111",
	213 => "11111111",
	214 => "11111111",
	215 => "11111111",
	216 => "11111111",
	217 => "11111111",
	218 => "11111111",
	219 => "11111111",
	220 => "11111111",
	221 => "11111111",
	222 => "11111111",
	223 => "11111111",
	224 => "11111111",
	225 => "11111111",
	226 => "11111111",
	227 => "11111111",
	228 => "11111111",
	229 => "11111111",
	230 => "11111111",
	231 => "11111111",
	232 => "11111111",
	233 => "11111111",
	234 => "11111111",
	235 => "11111111",
	236 => "11111111",
	237 => "11111111",
	238 => "11111111",
	239 => "11111111",
	240 => "11111111",
	241 => "11111111",
	242 => "11111111",
	243 => "11111111",
	244 => "11111111",
	245 => "11111111",
	246 => "11111111",
	247 => "11111111",
	256 => "11111111",
	257 => "11111111",
	258 => "11111111",
	259 => "11111111",
	260 => "11111111",
	261 => "11111111",
	262 => "11111111",
	263 => "11111111",
	264 => "11111111",
	265 => "11111111",
	266 => "11111111",
	267 => "11111111",
	268 => "11111111",
	269 => "11111111",
	270 => "11111111",
	271 => "11111111",
	272 => "11111111",
	273 => "11111111",
	274 => "11111111",
	275 => "11111111",
	276 => "11111111",
	277 => "11111111",
	278 => "11111111",
	279 => "11111111",
	280 => "11111111",
	281 => "11111111",
	282 => "11111111",
	283 => "11111111",
	284 => "11111111",
	285 => "11111111",
	286 => "11111111",
	287 => "11111111",
	288 => "11111111",
	289 => "11111111",
	290 => "11111111",
	291 => "11111111",
	292 => "11111111",
	293 => "11111111",
	294 => "11111111",
	295 => "11111111",
	296 => "11111111",
	297 => "11111111",
	298 => "11111111",
	299 => "11111111",
	300 => "11111111",
	301 => "11111111",
	302 => "11111111",
	303 => "11111111",
	304 => "11111111",
	305 => "11111111",
	306 => "11111111",
	307 => "11111111",
	308 => "11111111",
	309 => "11111111",
	310 => "11111111",
	311 => "11111111",
	312 => "11111111",
	313 => "11111111",
	314 => "11111111",
	315 => "11111111",
	316 => "11111111",
	317 => "11111111",
	318 => "11111111",
	319 => "11111111",
	320 => "11111111",
	321 => "11111111",
	322 => "11111111",
	323 => "11111111",
	324 => "11111111",
	325 => "11111111",
	326 => "11111111",
	327 => "11111111",
	328 => "11111111",
	329 => "11111111",
	330 => "11111111",
	331 => "11111111",
	332 => "11111111",
	333 => "11111111",
	334 => "11111111",
	335 => "11111111",
	336 => "11111111",
	337 => "11111111",
	338 => "11111111",
	339 => "11111111",
	340 => "11111111",
	341 => "11111111",
	342 => "11111111",
	343 => "11111111",
	344 => "11111111",
	345 => "11111111",
	346 => "11111111",
	347 => "11111111",
	348 => "11111111",
	349 => "11111111",
	350 => "11111111",
	351 => "11111111",
	352 => "11111111",
	353 => "11111111",
	354 => "11111111",
	355 => "11111111",
	356 => "11111111",
	357 => "11111111",
	358 => "11111111",
	359 => "11111111",
	360 => "11111111",
	361 => "11111111",
	362 => "11111111",
	363 => "11111111",
	364 => "11111111",
	365 => "11111111",
	366 => "11111111",
	367 => "11111111",
	368 => "11111111",
	369 => "11111111",
	370 => "11111111",
	371 => "11111111",
	372 => "11111111",
	373 => "11111111",
	374 => "11111111",
	375 => "11111111",
	384 => "11111111",
	385 => "11111111",
	386 => "11111111",
	387 => "11111111",
	388 => "11111111",
	389 => "11111111",
	390 => "11111111",
	391 => "11111111",
	392 => "11111111",
	393 => "11111111",
	394 => "11111111",
	395 => "11111111",
	396 => "11111111",
	397 => "11111111",
	398 => "11111111",
	399 => "11111111",
	400 => "11111111",
	401 => "11111111",
	402 => "11111111",
	403 => "11111111",
	404 => "11111111",
	405 => "11111111",
	406 => "11111111",
	407 => "11111111",
	408 => "11111111",
	409 => "11111111",
	410 => "11111111",
	411 => "11111111",
	412 => "11111111",
	413 => "11111111",
	414 => "11111111",
	415 => "11111111",
	416 => "11111111",
	417 => "11111111",
	418 => "11111111",
	419 => "11111111",
	420 => "11111111",
	421 => "11111111",
	422 => "11111111",
	423 => "11111111",
	424 => "11111111",
	425 => "11111111",
	426 => "11111111",
	427 => "11111111",
	428 => "11111111",
	429 => "11111111",
	430 => "11111111",
	431 => "11111111",
	432 => "11111111",
	433 => "11111111",
	434 => "11111111",
	435 => "11111111",
	436 => "11111111",
	437 => "11111111",
	438 => "11111111",
	439 => "11111111",
	440 => "11111111",
	441 => "11111111",
	442 => "11111111",
	443 => "11111111",
	444 => "11111111",
	445 => "11111111",
	446 => "11111111",
	447 => "11111111",
	448 => "11111111",
	449 => "11111111",
	450 => "11111111",
	451 => "11111111",
	452 => "11111111",
	453 => "11111111",
	454 => "11111111",
	455 => "11111111",
	456 => "11111111",
	457 => "11111111",
	458 => "11111111",
	459 => "11111111",
	460 => "11111111",
	461 => "11111111",
	462 => "11111111",
	463 => "11111111",
	464 => "11111111",
	465 => "11111111",
	466 => "11111111",
	467 => "11111111",
	468 => "11111111",
	469 => "11111111",
	470 => "11111111",
	471 => "11111111",
	472 => "11111111",
	473 => "11111111",
	474 => "11111111",
	475 => "11111111",
	476 => "11111111",
	477 => "11111111",
	478 => "11111111",
	479 => "11111111",
	480 => "11111111",
	481 => "11111111",
	482 => "11111111",
	483 => "11111111",
	484 => "11111111",
	485 => "11111111",
	486 => "11111111",
	487 => "11111111",
	488 => "11111111",
	489 => "11111111",
	490 => "11111111",
	491 => "11111111",
	492 => "11111111",
	493 => "11111111",
	494 => "11111111",
	495 => "11111111",
	496 => "11111111",
	497 => "11111111",
	498 => "11111111",
	499 => "11111111",
	500 => "11111111",
	501 => "11111111",
	502 => "11111111",
	503 => "11111111",
	512 => "11111111",
	513 => "11111111",
	514 => "11111111",
	515 => "11111111",
	516 => "11111111",
	517 => "11111111",
	518 => "11111111",
	519 => "11111111",
	520 => "11111111",
	521 => "11111111",
	522 => "11111111",
	523 => "11111111",
	524 => "11111111",
	525 => "11111111",
	526 => "11111111",
	527 => "11111111",
	528 => "11111111",
	529 => "11111111",
	530 => "11111111",
	531 => "11111111",
	532 => "11111111",
	533 => "11111111",
	534 => "11111111",
	535 => "11111111",
	536 => "11111111",
	537 => "11111111",
	538 => "11111111",
	539 => "11111111",
	540 => "11111111",
	541 => "11111111",
	542 => "11111111",
	543 => "11111111",
	544 => "11111111",
	545 => "11111111",
	546 => "11111111",
	547 => "11111111",
	548 => "11111111",
	549 => "11111111",
	550 => "11111111",
	551 => "11111111",
	552 => "11111111",
	553 => "11111111",
	554 => "11111111",
	555 => "11111111",
	556 => "11111111",
	557 => "11111111",
	558 => "11111111",
	559 => "11111111",
	560 => "11111111",
	561 => "11111111",
	562 => "11111111",
	563 => "11111111",
	564 => "11111111",
	565 => "11111111",
	566 => "11111111",
	567 => "11111111",
	568 => "11111111",
	569 => "11111111",
	570 => "11111111",
	571 => "11111111",
	572 => "11111111",
	573 => "11111111",
	574 => "11111111",
	575 => "11111111",
	576 => "11111111",
	577 => "11111111",
	578 => "11111111",
	579 => "11111111",
	580 => "11111111",
	581 => "11111111",
	582 => "11111111",
	583 => "11111111",
	584 => "11111111",
	585 => "11111111",
	586 => "11111111",
	587 => "11111111",
	588 => "11111111",
	589 => "11111111",
	590 => "11111111",
	591 => "11111111",
	592 => "11111111",
	593 => "11111111",
	594 => "11111111",
	595 => "11111111",
	596 => "11111111",
	597 => "11111111",
	598 => "11111111",
	599 => "11111111",
	600 => "11111111",
	601 => "11111111",
	602 => "11111111",
	603 => "11111111",
	604 => "11111111",
	605 => "11111111",
	606 => "11111111",
	607 => "11111111",
	608 => "11111111",
	609 => "11111111",
	610 => "11111111",
	611 => "11111111",
	612 => "11111111",
	613 => "11111111",
	614 => "11111111",
	615 => "11111111",
	616 => "11111111",
	617 => "11111111",
	618 => "11111111",
	619 => "11111111",
	620 => "11111111",
	621 => "11111111",
	622 => "11111111",
	623 => "11111111",
	624 => "11111111",
	625 => "11111111",
	626 => "11111111",
	627 => "11111111",
	628 => "11111111",
	629 => "11111111",
	630 => "11111111",
	631 => "11111111",
	640 => "11111111",
	641 => "11111111",
	642 => "11111111",
	643 => "11111111",
	644 => "11111111",
	645 => "11111111",
	646 => "11111111",
	647 => "11111111",
	648 => "11111111",
	649 => "11111111",
	650 => "11111111",
	651 => "11111111",
	652 => "11111111",
	653 => "11111111",
	654 => "11111111",
	655 => "11111111",
	656 => "11111111",
	657 => "11111111",
	658 => "11111111",
	659 => "11111111",
	660 => "11111111",
	661 => "11111111",
	662 => "11111111",
	663 => "11111111",
	664 => "11111111",
	665 => "11111111",
	666 => "11111111",
	667 => "11111111",
	668 => "11111111",
	669 => "11111111",
	670 => "11111111",
	671 => "11111111",
	672 => "11111111",
	673 => "11111111",
	674 => "11111111",
	675 => "11111111",
	676 => "11111111",
	677 => "11111111",
	678 => "11111111",
	679 => "11111111",
	680 => "11111111",
	681 => "11111111",
	682 => "11111111",
	683 => "11111111",
	684 => "11111111",
	685 => "11111111",
	686 => "11111111",
	687 => "11111111",
	688 => "11111111",
	689 => "11111111",
	690 => "11111111",
	691 => "11111111",
	692 => "11111111",
	693 => "11111111",
	694 => "11111111",
	695 => "11111111",
	696 => "11111111",
	697 => "11111111",
	698 => "11111111",
	699 => "11111111",
	700 => "11111111",
	701 => "11111111",
	702 => "11111111",
	703 => "11111111",
	704 => "11111111",
	705 => "11111111",
	706 => "11111111",
	707 => "11111111",
	708 => "11111111",
	709 => "11111111",
	710 => "11111111",
	711 => "11111111",
	712 => "11111111",
	713 => "11111111",
	714 => "11111111",
	715 => "11111111",
	716 => "11111111",
	717 => "11111111",
	718 => "11111111",
	719 => "11111111",
	720 => "11111111",
	721 => "11111111",
	722 => "11111111",
	723 => "11111111",
	724 => "11111111",
	725 => "11111111",
	726 => "11111111",
	727 => "11111111",
	728 => "11111111",
	729 => "11111111",
	730 => "11111111",
	731 => "11111111",
	732 => "11111111",
	733 => "11111111",
	734 => "11111111",
	735 => "11111111",
	736 => "11111111",
	737 => "11111111",
	738 => "11111111",
	739 => "11111111",
	740 => "11111111",
	741 => "11111111",
	742 => "11111111",
	743 => "11111111",
	744 => "11111111",
	745 => "11111111",
	746 => "11111111",
	747 => "11111111",
	748 => "11111111",
	749 => "11111111",
	750 => "11111111",
	751 => "11111111",
	752 => "11111111",
	753 => "11111111",
	754 => "11111111",
	755 => "11111111",
	756 => "11111111",
	757 => "11111111",
	758 => "11111111",
	759 => "11111111",
	768 => "11111111",
	769 => "11111111",
	770 => "11111111",
	771 => "11111111",
	772 => "11111111",
	773 => "11111111",
	774 => "11111111",
	775 => "11111111",
	776 => "11111111",
	777 => "11111111",
	778 => "11111111",
	779 => "11111111",
	780 => "11111111",
	781 => "11111111",
	782 => "11111111",
	783 => "11111111",
	784 => "11111111",
	785 => "11111111",
	786 => "11111111",
	787 => "11111111",
	788 => "11111111",
	789 => "11111111",
	790 => "11111111",
	791 => "11111111",
	792 => "11111111",
	793 => "11111111",
	794 => "11111111",
	795 => "11111111",
	796 => "11111111",
	797 => "11111111",
	798 => "11111111",
	799 => "11111111",
	800 => "11111111",
	801 => "11111111",
	802 => "11111111",
	803 => "11111111",
	804 => "11111111",
	805 => "11111111",
	806 => "11111111",
	807 => "11111111",
	808 => "11111111",
	809 => "11111111",
	810 => "11111111",
	811 => "11111111",
	812 => "11111111",
	813 => "11111111",
	814 => "11111111",
	815 => "11111111",
	816 => "11111111",
	817 => "11111111",
	818 => "11111111",
	819 => "11111111",
	820 => "11111111",
	821 => "11111111",
	822 => "11111111",
	823 => "11111111",
	824 => "11111111",
	825 => "11111111",
	826 => "11111111",
	827 => "11111111",
	828 => "11111111",
	829 => "11111111",
	830 => "11111111",
	831 => "11111111",
	832 => "11111111",
	833 => "11111111",
	834 => "11111111",
	835 => "11111111",
	836 => "11111111",
	837 => "11111111",
	838 => "11111111",
	839 => "11111111",
	840 => "11111111",
	841 => "11111111",
	842 => "11111111",
	843 => "11111111",
	844 => "11111111",
	845 => "11111111",
	846 => "11111111",
	847 => "11111111",
	848 => "11111111",
	849 => "11111111",
	850 => "11111111",
	851 => "11111111",
	852 => "11111111",
	853 => "11111111",
	854 => "11111111",
	855 => "11111111",
	856 => "11111111",
	857 => "11111111",
	858 => "11111111",
	859 => "11111111",
	860 => "11111111",
	861 => "11111111",
	862 => "11111111",
	863 => "11111111",
	864 => "11111111",
	865 => "11111111",
	866 => "11111111",
	867 => "11111111",
	868 => "11111111",
	869 => "11111111",
	870 => "11111111",
	871 => "11111111",
	872 => "11111111",
	873 => "11111111",
	874 => "11111111",
	875 => "11111111",
	876 => "11111111",
	877 => "11111111",
	878 => "11111111",
	879 => "11111111",
	880 => "11111111",
	881 => "11111111",
	882 => "11111111",
	883 => "11111111",
	884 => "11111111",
	885 => "11111111",
	886 => "11111111",
	887 => "11111111",
	896 => "11111111",
	897 => "11111111",
	898 => "11111111",
	899 => "11111111",
	900 => "11111111",
	901 => "11111111",
	902 => "11111111",
	903 => "11111111",
	904 => "11111111",
	905 => "11111111",
	906 => "11111111",
	907 => "11111111",
	908 => "11111111",
	909 => "11111111",
	910 => "11111111",
	911 => "11111111",
	912 => "11111111",
	913 => "11111111",
	914 => "11111111",
	915 => "11111111",
	916 => "11111111",
	917 => "11111111",
	918 => "11111111",
	919 => "11111111",
	920 => "11111111",
	921 => "11111111",
	922 => "11111111",
	923 => "11111111",
	924 => "11111111",
	925 => "11111111",
	926 => "11111111",
	927 => "11111111",
	928 => "11111111",
	929 => "11111111",
	930 => "11111111",
	931 => "11111111",
	932 => "11111111",
	933 => "11111111",
	934 => "11111111",
	935 => "11111111",
	936 => "11111111",
	937 => "11111111",
	938 => "11111111",
	939 => "11111111",
	940 => "11111111",
	941 => "11111111",
	942 => "11111111",
	943 => "11111111",
	944 => "11111111",
	945 => "11111111",
	946 => "11111111",
	947 => "11111111",
	948 => "11111111",
	949 => "11111111",
	950 => "11111111",
	951 => "11111111",
	952 => "11111111",
	953 => "11111111",
	954 => "11111111",
	955 => "11111111",
	956 => "11111111",
	957 => "11111111",
	958 => "11111111",
	959 => "11111111",
	960 => "11111111",
	961 => "11111111",
	962 => "11111111",
	963 => "11111111",
	964 => "11111111",
	965 => "11111111",
	966 => "11111111",
	967 => "11111111",
	968 => "11111111",
	969 => "11111111",
	970 => "11111111",
	971 => "11111111",
	972 => "11111111",
	973 => "11111111",
	974 => "11111111",
	975 => "11111111",
	976 => "11111111",
	977 => "11111111",
	978 => "11111111",
	979 => "11111111",
	980 => "11111111",
	981 => "11111111",
	982 => "11111111",
	983 => "11111111",
	984 => "11111111",
	985 => "11111111",
	986 => "11111111",
	987 => "11111111",
	988 => "11111111",
	989 => "11111111",
	990 => "11111111",
	991 => "11111111",
	992 => "11111111",
	993 => "11111111",
	994 => "11111111",
	995 => "11111111",
	996 => "11111111",
	997 => "11111111",
	998 => "11111111",
	999 => "11111111",
	1000 => "11111111",
	1001 => "11111111",
	1002 => "11111111",
	1003 => "11111111",
	1004 => "11111111",
	1005 => "11111111",
	1006 => "11111111",
	1007 => "11111111",
	1008 => "11111111",
	1009 => "11111111",
	1010 => "11111111",
	1011 => "11111111",
	1012 => "11111111",
	1013 => "11111111",
	1014 => "11111111",
	1015 => "11111111",
	1024 => "11111111",
	1025 => "11111111",
	1026 => "11111111",
	1027 => "11111111",
	1028 => "11111111",
	1029 => "11111111",
	1030 => "11111111",
	1031 => "11111111",
	1032 => "11111111",
	1033 => "11111111",
	1034 => "11111111",
	1035 => "11111111",
	1036 => "11111111",
	1037 => "11111111",
	1038 => "11111111",
	1039 => "11111111",
	1040 => "11111111",
	1041 => "11111111",
	1042 => "11111111",
	1043 => "11111111",
	1044 => "11111111",
	1045 => "11111111",
	1046 => "11111111",
	1047 => "11111111",
	1048 => "11111111",
	1049 => "11111111",
	1050 => "11111111",
	1051 => "11111111",
	1052 => "11111111",
	1053 => "11111111",
	1054 => "11111111",
	1055 => "11111111",
	1056 => "11111111",
	1057 => "11111111",
	1058 => "11111111",
	1059 => "11111111",
	1060 => "11111111",
	1061 => "11111111",
	1062 => "11111111",
	1063 => "11111111",
	1064 => "11111111",
	1065 => "11111111",
	1066 => "11111111",
	1067 => "11111111",
	1068 => "11111111",
	1069 => "11111111",
	1070 => "11111111",
	1071 => "11111111",
	1072 => "11111111",
	1073 => "11111111",
	1074 => "11111111",
	1075 => "11111111",
	1076 => "11111111",
	1077 => "11111111",
	1078 => "11111111",
	1079 => "11111111",
	1080 => "11111111",
	1081 => "11111111",
	1082 => "11111111",
	1083 => "11111111",
	1084 => "11111111",
	1085 => "11111111",
	1086 => "11111111",
	1087 => "11111111",
	1088 => "11111111",
	1089 => "11111111",
	1090 => "11111111",
	1091 => "11111111",
	1092 => "11111111",
	1093 => "11111111",
	1094 => "11111111",
	1095 => "11111111",
	1096 => "11111111",
	1097 => "11111111",
	1098 => "11111111",
	1099 => "11111111",
	1100 => "11111111",
	1101 => "11111111",
	1102 => "11111111",
	1103 => "11111111",
	1104 => "11111111",
	1105 => "11111111",
	1106 => "11111111",
	1107 => "11111111",
	1108 => "11111111",
	1109 => "11111111",
	1110 => "11111111",
	1111 => "11111111",
	1112 => "11111111",
	1113 => "11111111",
	1114 => "11111111",
	1115 => "11111111",
	1116 => "11111111",
	1117 => "11111111",
	1118 => "11111111",
	1119 => "11111111",
	1120 => "11111111",
	1121 => "11111111",
	1122 => "11111111",
	1123 => "11111111",
	1124 => "11111111",
	1125 => "11111111",
	1126 => "11111111",
	1127 => "11111111",
	1128 => "11111111",
	1129 => "11111111",
	1130 => "11111111",
	1131 => "11111111",
	1132 => "11111111",
	1133 => "11111111",
	1134 => "11111111",
	1135 => "11111111",
	1136 => "11111111",
	1137 => "11111111",
	1138 => "11111111",
	1139 => "11111111",
	1140 => "11111111",
	1141 => "11111111",
	1142 => "11111111",
	1143 => "11111111",
	1152 => "11111111",
	1153 => "11111111",
	1154 => "11111111",
	1155 => "11111111",
	1156 => "11111111",
	1157 => "11111111",
	1158 => "11111111",
	1159 => "11111111",
	1160 => "11111111",
	1161 => "11111111",
	1162 => "11111111",
	1163 => "11111111",
	1164 => "11111111",
	1165 => "11111111",
	1166 => "11111111",
	1167 => "11111111",
	1168 => "11111111",
	1169 => "11111111",
	1170 => "11111111",
	1171 => "11111111",
	1172 => "11111111",
	1173 => "11111111",
	1174 => "11111111",
	1175 => "11111111",
	1176 => "11111111",
	1177 => "11111111",
	1178 => "11111111",
	1179 => "11111111",
	1180 => "11111111",
	1181 => "11111111",
	1182 => "11111111",
	1183 => "11111111",
	1184 => "11111111",
	1185 => "11111111",
	1186 => "11111111",
	1187 => "11111111",
	1188 => "11111111",
	1189 => "11111111",
	1190 => "11111111",
	1191 => "11111111",
	1192 => "11111111",
	1193 => "11111111",
	1194 => "11111111",
	1195 => "11111111",
	1196 => "11111111",
	1197 => "11111111",
	1198 => "11111111",
	1199 => "11111111",
	1200 => "11111111",
	1201 => "11111111",
	1202 => "11111111",
	1203 => "11111111",
	1204 => "11111111",
	1205 => "11111111",
	1206 => "11111111",
	1207 => "11111111",
	1208 => "11111111",
	1209 => "11111111",
	1210 => "11111111",
	1211 => "11111111",
	1212 => "11111111",
	1213 => "11111111",
	1214 => "11111111",
	1215 => "11111111",
	1216 => "11111111",
	1217 => "11111111",
	1218 => "11111111",
	1219 => "11111111",
	1220 => "11111111",
	1221 => "11111111",
	1222 => "11111111",
	1223 => "11111111",
	1224 => "11111111",
	1225 => "11111111",
	1226 => "11111111",
	1227 => "11111111",
	1228 => "11111111",
	1229 => "11111111",
	1230 => "11111111",
	1231 => "11111111",
	1232 => "11111111",
	1233 => "11111111",
	1234 => "11111111",
	1235 => "11111111",
	1236 => "11111111",
	1237 => "11111111",
	1238 => "11111111",
	1239 => "11111111",
	1240 => "11111111",
	1241 => "11111111",
	1242 => "11111111",
	1243 => "11111111",
	1244 => "11111111",
	1245 => "11111111",
	1246 => "11111111",
	1247 => "11111111",
	1248 => "11111111",
	1249 => "11111111",
	1250 => "11111111",
	1251 => "11111111",
	1252 => "11111111",
	1253 => "11111111",
	1254 => "11111111",
	1255 => "11111111",
	1256 => "11111111",
	1257 => "11111111",
	1258 => "11111111",
	1259 => "11111111",
	1260 => "11111111",
	1261 => "11111111",
	1262 => "11111111",
	1263 => "11111111",
	1264 => "11111111",
	1265 => "11111111",
	1266 => "11111111",
	1267 => "11111111",
	1268 => "11111111",
	1269 => "11111111",
	1270 => "11111111",
	1271 => "11111111",
	1280 => "11111111",
	1281 => "11111111",
	1282 => "11111111",
	1283 => "11111111",
	1284 => "11111111",
	1285 => "11111111",
	1286 => "11111111",
	1287 => "11111111",
	1288 => "11111111",
	1289 => "11111111",
	1290 => "11111111",
	1291 => "11111111",
	1292 => "11111111",
	1293 => "11111111",
	1294 => "11111111",
	1295 => "11111111",
	1296 => "11111111",
	1297 => "11111111",
	1298 => "11111111",
	1299 => "11111111",
	1300 => "11111111",
	1301 => "11111111",
	1302 => "11111111",
	1303 => "11111111",
	1304 => "11111111",
	1305 => "11111111",
	1306 => "11111111",
	1307 => "11111111",
	1308 => "11111111",
	1309 => "11111111",
	1310 => "11111111",
	1311 => "11111111",
	1312 => "11111111",
	1313 => "11111111",
	1314 => "11111111",
	1315 => "11111111",
	1316 => "11111111",
	1317 => "11111111",
	1318 => "11111111",
	1319 => "11111111",
	1320 => "11111111",
	1321 => "11111111",
	1322 => "11111111",
	1323 => "11111111",
	1324 => "11111111",
	1325 => "11111111",
	1326 => "11111111",
	1327 => "11111111",
	1328 => "11111111",
	1329 => "11111111",
	1330 => "11111111",
	1331 => "11111111",
	1332 => "11111111",
	1333 => "11111111",
	1334 => "11111111",
	1335 => "11111111",
	1336 => "11111111",
	1337 => "11111111",
	1338 => "11111111",
	1339 => "11111111",
	1340 => "11111111",
	1341 => "11111111",
	1342 => "11111111",
	1343 => "11111111",
	1344 => "11111111",
	1345 => "11111111",
	1346 => "11111111",
	1347 => "11111111",
	1348 => "11111111",
	1349 => "11111111",
	1350 => "11111111",
	1351 => "11111111",
	1352 => "11111111",
	1353 => "11111111",
	1354 => "11111111",
	1355 => "11111111",
	1356 => "11111111",
	1357 => "11111111",
	1358 => "11111111",
	1359 => "11111111",
	1360 => "11111111",
	1361 => "11111111",
	1362 => "11111111",
	1363 => "11111111",
	1364 => "11111111",
	1365 => "11111111",
	1366 => "11111111",
	1367 => "11111111",
	1368 => "11111111",
	1369 => "11111111",
	1370 => "11111111",
	1371 => "11111111",
	1372 => "11111111",
	1373 => "11111111",
	1374 => "11111111",
	1375 => "11111111",
	1376 => "11111111",
	1377 => "11111111",
	1378 => "11111111",
	1379 => "11111111",
	1380 => "11111111",
	1381 => "11111111",
	1382 => "11111111",
	1383 => "11111111",
	1384 => "11111111",
	1385 => "11111111",
	1386 => "11111111",
	1387 => "11111111",
	1388 => "11111111",
	1389 => "11111111",
	1390 => "11111111",
	1391 => "11111111",
	1392 => "11111111",
	1393 => "11111111",
	1394 => "11111111",
	1395 => "11111111",
	1396 => "11111111",
	1397 => "11111111",
	1398 => "11111111",
	1399 => "11111111",
	1408 => "11111111",
	1409 => "11111111",
	1410 => "11111111",
	1411 => "11111111",
	1412 => "11111111",
	1413 => "11111111",
	1414 => "11111111",
	1415 => "11111111",
	1416 => "11111111",
	1417 => "11111111",
	1418 => "11111111",
	1419 => "11111111",
	1420 => "11111111",
	1421 => "11111111",
	1422 => "11111111",
	1423 => "11111111",
	1424 => "11111111",
	1425 => "11111111",
	1426 => "11111111",
	1427 => "11111111",
	1428 => "11111111",
	1429 => "11111111",
	1430 => "11111111",
	1431 => "11111111",
	1432 => "11111111",
	1433 => "11111111",
	1434 => "11111111",
	1435 => "11111111",
	1436 => "11111111",
	1437 => "11111111",
	1438 => "11111111",
	1439 => "11111111",
	1440 => "11111111",
	1441 => "11111111",
	1442 => "11111111",
	1443 => "11111111",
	1444 => "11111111",
	1445 => "11111111",
	1446 => "11111111",
	1447 => "11111111",
	1448 => "11111111",
	1449 => "11111111",
	1450 => "11111111",
	1451 => "11111111",
	1452 => "11111111",
	1453 => "11111111",
	1454 => "11111111",
	1455 => "11111111",
	1456 => "11111111",
	1457 => "11111111",
	1458 => "11111111",
	1459 => "11111111",
	1460 => "11111111",
	1461 => "11111111",
	1462 => "11111111",
	1463 => "11111111",
	1464 => "11111111",
	1465 => "11111111",
	1466 => "11111111",
	1467 => "11111111",
	1468 => "11111111",
	1469 => "11111111",
	1470 => "11111111",
	1471 => "11111111",
	1472 => "11111111",
	1473 => "11111111",
	1474 => "11111111",
	1475 => "11111111",
	1476 => "11111111",
	1477 => "11111111",
	1478 => "11111111",
	1479 => "11111111",
	1480 => "11111111",
	1481 => "11111111",
	1482 => "11111111",
	1483 => "11111111",
	1484 => "11111111",
	1485 => "11111111",
	1486 => "11111111",
	1487 => "11111111",
	1488 => "11111111",
	1489 => "11111111",
	1490 => "11111111",
	1491 => "11111111",
	1492 => "11111111",
	1493 => "11111111",
	1494 => "11111111",
	1495 => "11111111",
	1496 => "11111111",
	1497 => "11111111",
	1498 => "11111111",
	1499 => "11111111",
	1500 => "11111111",
	1501 => "11111111",
	1502 => "11111111",
	1503 => "11111111",
	1504 => "11111111",
	1505 => "11111111",
	1506 => "11111111",
	1507 => "11111111",
	1508 => "11111111",
	1509 => "11111111",
	1510 => "11111111",
	1511 => "11111111",
	1512 => "11111111",
	1513 => "11111111",
	1514 => "11111111",
	1515 => "11111111",
	1516 => "11111111",
	1517 => "11111111",
	1518 => "11111111",
	1519 => "11111111",
	1520 => "11111111",
	1521 => "11111111",
	1522 => "11111111",
	1523 => "11111111",
	1524 => "11111111",
	1525 => "11111111",
	1526 => "11111111",
	1527 => "11111111",
	1536 => "11111111",
	1537 => "11111111",
	1538 => "11111111",
	1539 => "11111111",
	1540 => "11111111",
	1541 => "11111111",
	1542 => "11111111",
	1543 => "11111111",
	1544 => "11111111",
	1545 => "11111111",
	1546 => "11111111",
	1547 => "11111111",
	1548 => "11111111",
	1549 => "11111111",
	1550 => "11111111",
	1551 => "11111111",
	1552 => "11111111",
	1553 => "11111111",
	1554 => "11111111",
	1555 => "11111111",
	1556 => "11111111",
	1557 => "11111111",
	1558 => "11111111",
	1559 => "11111111",
	1560 => "11111111",
	1561 => "11111111",
	1562 => "11111111",
	1563 => "11111111",
	1564 => "11111111",
	1565 => "11111111",
	1566 => "11111111",
	1567 => "11111111",
	1568 => "11111111",
	1569 => "11111111",
	1570 => "11111111",
	1571 => "11111111",
	1572 => "11111111",
	1573 => "11111111",
	1574 => "11111111",
	1575 => "11111111",
	1576 => "11111111",
	1577 => "11111111",
	1578 => "11111111",
	1579 => "11111111",
	1580 => "11111111",
	1581 => "11111111",
	1582 => "11111111",
	1583 => "11111111",
	1584 => "11111111",
	1585 => "11111111",
	1586 => "11111111",
	1587 => "11111111",
	1588 => "11111111",
	1589 => "11111111",
	1590 => "11111111",
	1591 => "11111111",
	1592 => "11111111",
	1593 => "11111111",
	1594 => "11111111",
	1595 => "11111111",
	1596 => "11111111",
	1597 => "11111111",
	1598 => "11111111",
	1599 => "11111111",
	1600 => "11111111",
	1601 => "11111111",
	1602 => "11111111",
	1603 => "11111111",
	1604 => "11111111",
	1605 => "11111111",
	1606 => "11111111",
	1607 => "11111111",
	1608 => "11111111",
	1609 => "11111111",
	1610 => "11111111",
	1611 => "11111111",
	1612 => "11111111",
	1613 => "11111111",
	1614 => "11111111",
	1615 => "11111111",
	1616 => "11111111",
	1617 => "11111111",
	1618 => "11111111",
	1619 => "11111111",
	1620 => "11111111",
	1621 => "11111111",
	1622 => "11111111",
	1623 => "11111111",
	1624 => "11111111",
	1625 => "11111111",
	1626 => "11111111",
	1627 => "11111111",
	1628 => "11111111",
	1629 => "11111111",
	1630 => "11111111",
	1631 => "11111111",
	1632 => "11111111",
	1633 => "11111111",
	1634 => "11111111",
	1635 => "11111111",
	1636 => "11111111",
	1637 => "11111111",
	1638 => "11111111",
	1639 => "11111111",
	1640 => "11111111",
	1641 => "11111111",
	1642 => "11111111",
	1643 => "11111111",
	1644 => "11111111",
	1645 => "11111111",
	1646 => "11111111",
	1647 => "11111111",
	1648 => "11111111",
	1649 => "11111111",
	1650 => "11111111",
	1651 => "11111111",
	1652 => "11111111",
	1653 => "11111111",
	1654 => "11111111",
	1655 => "11111111",
	1664 => "11111111",
	1665 => "11111111",
	1666 => "11111111",
	1667 => "11111111",
	1668 => "11111111",
	1669 => "11111111",
	1670 => "11111111",
	1671 => "11111111",
	1672 => "11111111",
	1673 => "11111111",
	1674 => "11111111",
	1675 => "11111111",
	1676 => "11111111",
	1677 => "11111111",
	1678 => "11111111",
	1679 => "11111111",
	1680 => "11111111",
	1681 => "11111111",
	1682 => "11111111",
	1683 => "11111111",
	1684 => "11111111",
	1685 => "11111111",
	1686 => "11111111",
	1687 => "11111111",
	1688 => "11111111",
	1689 => "11111111",
	1690 => "11111111",
	1691 => "11111111",
	1692 => "11111111",
	1693 => "11111111",
	1694 => "11111111",
	1695 => "11111111",
	1696 => "11111111",
	1697 => "11111111",
	1698 => "11111111",
	1699 => "11111111",
	1700 => "11111111",
	1701 => "11111111",
	1702 => "11111111",
	1703 => "11111111",
	1704 => "11111111",
	1705 => "11111111",
	1706 => "11111111",
	1707 => "11111111",
	1708 => "11111111",
	1709 => "11111111",
	1710 => "11111111",
	1711 => "11111111",
	1712 => "11111111",
	1713 => "11111111",
	1714 => "11111111",
	1715 => "11111111",
	1716 => "11111111",
	1717 => "11111111",
	1718 => "11111111",
	1719 => "11111111",
	1720 => "11111111",
	1721 => "11111111",
	1722 => "11111111",
	1723 => "11111111",
	1724 => "11111111",
	1725 => "11111111",
	1726 => "11111111",
	1727 => "11111111",
	1728 => "11111111",
	1729 => "11111111",
	1730 => "11111111",
	1731 => "11111111",
	1732 => "11111111",
	1733 => "11111111",
	1734 => "11111111",
	1735 => "11111111",
	1736 => "11111111",
	1737 => "11111111",
	1738 => "11111111",
	1739 => "11111111",
	1740 => "11111111",
	1741 => "11111111",
	1742 => "11111111",
	1743 => "11111111",
	1744 => "11111111",
	1745 => "11111111",
	1746 => "11111111",
	1747 => "11111111",
	1748 => "11111111",
	1749 => "11111111",
	1750 => "11111111",
	1751 => "11111111",
	1752 => "11111111",
	1753 => "11111111",
	1754 => "11111111",
	1755 => "11111111",
	1756 => "11111111",
	1757 => "11111111",
	1758 => "11111111",
	1759 => "11111111",
	1760 => "11111111",
	1761 => "11111111",
	1762 => "11111111",
	1763 => "11111111",
	1764 => "11111111",
	1765 => "11111111",
	1766 => "11111111",
	1767 => "11111111",
	1768 => "11111111",
	1769 => "11111111",
	1770 => "11111111",
	1771 => "11111111",
	1772 => "11111111",
	1773 => "11111111",
	1774 => "11111111",
	1775 => "11111111",
	1776 => "11111111",
	1777 => "11111111",
	1778 => "11111111",
	1779 => "11111111",
	1780 => "11111111",
	1781 => "11111111",
	1782 => "11111111",
	1783 => "11111111",
	1792 => "11111111",
	1793 => "11111111",
	1794 => "11111111",
	1795 => "11111111",
	1796 => "11111111",
	1797 => "11111111",
	1798 => "11111111",
	1799 => "11111111",
	1800 => "11111111",
	1801 => "11111111",
	1802 => "11111111",
	1803 => "11111111",
	1804 => "11111111",
	1805 => "11111111",
	1806 => "11111111",
	1807 => "11111111",
	1808 => "11111111",
	1809 => "11111111",
	1810 => "11111111",
	1811 => "11111111",
	1812 => "11111111",
	1813 => "11111111",
	1814 => "11111111",
	1815 => "11111111",
	1816 => "11111111",
	1817 => "11111111",
	1818 => "11111111",
	1819 => "11111111",
	1820 => "11111111",
	1821 => "11111111",
	1822 => "11111111",
	1823 => "11111111",
	1824 => "11111111",
	1825 => "11111111",
	1826 => "11111111",
	1827 => "11111111",
	1828 => "11111111",
	1829 => "11111111",
	1830 => "11111111",
	1831 => "11111111",
	1832 => "11111111",
	1833 => "11111111",
	1834 => "11111111",
	1835 => "11111111",
	1836 => "11111111",
	1837 => "11111111",
	1838 => "11111111",
	1839 => "11111111",
	1840 => "11111111",
	1841 => "11111111",
	1842 => "11111111",
	1843 => "11111111",
	1844 => "11111111",
	1845 => "11111111",
	1846 => "11111111",
	1847 => "11111111",
	1848 => "11111111",
	1849 => "11111111",
	1850 => "11111111",
	1851 => "11111111",
	1852 => "11111111",
	1853 => "11111111",
	1854 => "11111111",
	1855 => "11111111",
	1856 => "11111111",
	1857 => "11111111",
	1858 => "11111111",
	1859 => "11111111",
	1860 => "11111111",
	1861 => "11111111",
	1862 => "11111111",
	1863 => "11111111",
	1864 => "11111111",
	1865 => "11111111",
	1866 => "11111111",
	1867 => "11111111",
	1868 => "11111111",
	1869 => "11111111",
	1870 => "11111111",
	1871 => "11111111",
	1872 => "11111111",
	1873 => "11111111",
	1874 => "11111111",
	1875 => "11111111",
	1876 => "11111111",
	1877 => "11111111",
	1878 => "11111111",
	1879 => "11111111",
	1880 => "11111111",
	1881 => "11111111",
	1882 => "11111111",
	1883 => "11111111",
	1884 => "11111111",
	1885 => "11111111",
	1886 => "11111111",
	1887 => "11111111",
	1888 => "11111111",
	1889 => "11111111",
	1890 => "11111111",
	1891 => "11111111",
	1892 => "11111111",
	1893 => "11111111",
	1894 => "11111111",
	1895 => "11111111",
	1896 => "11111111",
	1897 => "11111111",
	1898 => "11111111",
	1899 => "11111111",
	1900 => "11111111",
	1901 => "11111111",
	1902 => "11111111",
	1903 => "11111111",
	1904 => "11111111",
	1905 => "11111111",
	1906 => "11111111",
	1907 => "11111111",
	1908 => "11111111",
	1909 => "11111111",
	1910 => "11111111",
	1911 => "11111111",
	1920 => "11111111",
	1921 => "11111111",
	1922 => "11111111",
	1923 => "11111111",
	1924 => "11111111",
	1925 => "11111111",
	1926 => "11111111",
	1927 => "11111111",
	1928 => "11111111",
	1929 => "11111111",
	1930 => "11111111",
	1931 => "11111111",
	1932 => "11111111",
	1933 => "11111111",
	1934 => "11111111",
	1935 => "11111111",
	1936 => "11111111",
	1937 => "11111111",
	1938 => "11111111",
	1939 => "11111111",
	1940 => "11111111",
	1941 => "11111111",
	1942 => "11111111",
	1943 => "11111111",
	1944 => "11111111",
	1945 => "11111111",
	1946 => "11111111",
	1947 => "11111111",
	1948 => "11111111",
	1949 => "11111111",
	1950 => "11111111",
	1951 => "11111111",
	1952 => "11111111",
	1953 => "11111111",
	1954 => "11111111",
	1955 => "11111111",
	1956 => "11111111",
	1957 => "11111111",
	1958 => "11111111",
	1959 => "11111111",
	1960 => "11111111",
	1961 => "11111111",
	1962 => "11111111",
	1963 => "11111111",
	1964 => "11111111",
	1965 => "11111111",
	1966 => "11111111",
	1967 => "11111111",
	1968 => "11111111",
	1969 => "11111111",
	1970 => "11111111",
	1971 => "11111111",
	1972 => "11111111",
	1973 => "11111111",
	1974 => "11111111",
	1975 => "11111111",
	1976 => "11111111",
	1977 => "11111111",
	1978 => "11111111",
	1979 => "11111111",
	1980 => "11111111",
	1981 => "11111111",
	1982 => "11111111",
	1983 => "11111111",
	1984 => "11111111",
	1985 => "11111111",
	1986 => "11111111",
	1987 => "11111111",
	1988 => "11111111",
	1989 => "11111111",
	1990 => "11111111",
	1991 => "11111111",
	1992 => "11111111",
	1993 => "11111111",
	1994 => "11111111",
	1995 => "11111111",
	1996 => "11111111",
	1997 => "11111111",
	1998 => "11111111",
	1999 => "11111111",
	2000 => "11111111",
	2001 => "11111111",
	2002 => "11111111",
	2003 => "11111111",
	2004 => "11111111",
	2005 => "11111111",
	2006 => "11111111",
	2007 => "11111111",
	2008 => "11111111",
	2009 => "11111111",
	2010 => "11111111",
	2011 => "11111111",
	2012 => "11111111",
	2013 => "11111111",
	2014 => "11111111",
	2015 => "11111111",
	2016 => "11111111",
	2017 => "11111111",
	2018 => "11111111",
	2019 => "11111111",
	2020 => "11111111",
	2021 => "11111111",
	2022 => "11111111",
	2023 => "11111111",
	2024 => "11111111",
	2025 => "11111111",
	2026 => "11111111",
	2027 => "11111111",
	2028 => "11111111",
	2029 => "11111111",
	2030 => "11111111",
	2031 => "11111111",
	2032 => "11111111",
	2033 => "11111111",
	2034 => "11111111",
	2035 => "11111111",
	2036 => "11111111",
	2037 => "11111111",
	2038 => "11111111",
	2039 => "11111111",
	2048 => "11111111",
	2049 => "11111111",
	2050 => "11111111",
	2051 => "11111111",
	2052 => "11111111",
	2053 => "11111111",
	2054 => "11111111",
	2055 => "11111111",
	2056 => "11111111",
	2057 => "11111111",
	2058 => "11111111",
	2059 => "11111111",
	2060 => "11111111",
	2061 => "11111111",
	2062 => "11111111",
	2063 => "11111111",
	2064 => "11111111",
	2065 => "11111111",
	2066 => "11111111",
	2067 => "11111111",
	2068 => "11111111",
	2069 => "11111111",
	2070 => "11111111",
	2071 => "11111111",
	2072 => "11111111",
	2073 => "11111111",
	2074 => "11111111",
	2075 => "11111111",
	2076 => "11111111",
	2077 => "11111111",
	2078 => "11111111",
	2079 => "11111111",
	2080 => "11111111",
	2081 => "11111111",
	2082 => "11111111",
	2083 => "11111111",
	2084 => "11111111",
	2085 => "11111111",
	2086 => "11111111",
	2087 => "11111111",
	2088 => "11111111",
	2089 => "11111111",
	2090 => "11111111",
	2091 => "11111111",
	2092 => "11111111",
	2093 => "11111111",
	2094 => "11111111",
	2095 => "11111111",
	2096 => "11111111",
	2097 => "11111111",
	2098 => "11111111",
	2099 => "11111111",
	2100 => "11111111",
	2101 => "11111111",
	2102 => "11111111",
	2103 => "11111111",
	2104 => "11111111",
	2105 => "11111111",
	2106 => "11111111",
	2107 => "11111111",
	2108 => "11111111",
	2109 => "11111111",
	2110 => "11111111",
	2111 => "11111111",
	2112 => "11111111",
	2113 => "11111111",
	2114 => "11111111",
	2115 => "11111111",
	2116 => "11111111",
	2117 => "11111111",
	2118 => "11111111",
	2119 => "11111111",
	2120 => "11111111",
	2121 => "11111111",
	2122 => "11111111",
	2123 => "11111111",
	2124 => "11111111",
	2125 => "11111111",
	2126 => "11111111",
	2127 => "11111111",
	2128 => "11111111",
	2129 => "11111111",
	2130 => "11111111",
	2131 => "11111111",
	2132 => "11111111",
	2133 => "11111111",
	2134 => "11111111",
	2135 => "11111111",
	2136 => "11111111",
	2137 => "11111111",
	2138 => "11111111",
	2139 => "11111111",
	2140 => "11111111",
	2141 => "11111111",
	2142 => "11111111",
	2143 => "11111111",
	2144 => "11111111",
	2145 => "11111111",
	2146 => "11111111",
	2147 => "11111111",
	2148 => "11111111",
	2149 => "11111111",
	2150 => "11111111",
	2151 => "11111111",
	2152 => "11111111",
	2153 => "11111111",
	2154 => "11111111",
	2155 => "11111111",
	2156 => "11111111",
	2157 => "11111111",
	2158 => "11111111",
	2159 => "11111111",
	2160 => "11111111",
	2161 => "11111111",
	2162 => "11111111",
	2163 => "11111111",
	2164 => "11111111",
	2165 => "11111111",
	2166 => "11111111",
	2167 => "11111111",
	2176 => "11111111",
	2177 => "11111111",
	2178 => "11111111",
	2179 => "11111111",
	2180 => "11111111",
	2181 => "11111111",
	2182 => "11111111",
	2183 => "11111111",
	2184 => "11111111",
	2185 => "11111111",
	2186 => "11111111",
	2187 => "11111111",
	2188 => "11111111",
	2189 => "11111111",
	2190 => "11111111",
	2191 => "11111111",
	2192 => "11111111",
	2193 => "11111111",
	2194 => "11111111",
	2195 => "11111111",
	2196 => "11111111",
	2197 => "11111111",
	2198 => "11111111",
	2199 => "11111111",
	2200 => "11111111",
	2201 => "11111111",
	2202 => "11111111",
	2203 => "11111111",
	2204 => "11111111",
	2205 => "11111111",
	2206 => "11111111",
	2207 => "11111111",
	2208 => "11111111",
	2209 => "11111111",
	2210 => "11111111",
	2211 => "11111111",
	2212 => "11111111",
	2213 => "11111111",
	2214 => "11111111",
	2215 => "11111111",
	2216 => "11111111",
	2217 => "11111111",
	2218 => "11111111",
	2219 => "11111111",
	2220 => "11111111",
	2221 => "11111111",
	2222 => "11111111",
	2223 => "11111111",
	2224 => "11111111",
	2225 => "11111111",
	2226 => "11111111",
	2227 => "11111111",
	2228 => "11111111",
	2229 => "11111111",
	2230 => "11111111",
	2231 => "11111111",
	2232 => "11111111",
	2233 => "11111111",
	2234 => "11111111",
	2235 => "11111111",
	2236 => "11111111",
	2237 => "11111111",
	2238 => "11111111",
	2239 => "11111111",
	2240 => "11111111",
	2241 => "11111111",
	2242 => "11111111",
	2243 => "11111111",
	2244 => "11111111",
	2245 => "11111111",
	2246 => "11111111",
	2247 => "11111111",
	2248 => "11111111",
	2249 => "11111111",
	2250 => "11111111",
	2251 => "11111111",
	2252 => "11111111",
	2253 => "11111111",
	2254 => "11111111",
	2255 => "11111111",
	2256 => "11111111",
	2257 => "11111111",
	2258 => "11111111",
	2259 => "11111111",
	2260 => "11111111",
	2261 => "11111111",
	2262 => "11111111",
	2263 => "11111111",
	2264 => "11111111",
	2265 => "11111111",
	2266 => "11111111",
	2267 => "11111111",
	2268 => "11111111",
	2269 => "11111111",
	2270 => "11111111",
	2271 => "11111111",
	2272 => "11111111",
	2273 => "11111111",
	2274 => "11111111",
	2275 => "11111111",
	2276 => "11111111",
	2277 => "11111111",
	2278 => "11111111",
	2279 => "11111111",
	2280 => "11111111",
	2281 => "11111111",
	2282 => "11111111",
	2283 => "11111111",
	2284 => "11111111",
	2285 => "11111111",
	2286 => "11111111",
	2287 => "11111111",
	2288 => "11111111",
	2289 => "11111111",
	2290 => "11111111",
	2291 => "11111111",
	2292 => "11111111",
	2293 => "11111111",
	2294 => "11111111",
	2295 => "11111111",
	2304 => "11111111",
	2305 => "11111111",
	2306 => "11111111",
	2307 => "11111111",
	2308 => "11111111",
	2309 => "11111111",
	2310 => "11111111",
	2311 => "11111111",
	2312 => "11111111",
	2313 => "11111111",
	2314 => "11111111",
	2315 => "11111111",
	2316 => "11111111",
	2317 => "11111111",
	2318 => "11111111",
	2319 => "11111111",
	2320 => "11111111",
	2321 => "11111111",
	2322 => "11111111",
	2323 => "11111111",
	2324 => "11111111",
	2325 => "11111111",
	2326 => "11111111",
	2327 => "11111111",
	2328 => "11111111",
	2329 => "11111111",
	2330 => "11111111",
	2331 => "11111111",
	2332 => "11111111",
	2333 => "11111111",
	2334 => "11111111",
	2335 => "11111111",
	2336 => "11111111",
	2337 => "11111111",
	2338 => "11111111",
	2339 => "11111111",
	2340 => "11111111",
	2341 => "11111111",
	2342 => "11111111",
	2343 => "11111111",
	2344 => "11111111",
	2345 => "11111111",
	2346 => "11111111",
	2347 => "11111111",
	2348 => "11111111",
	2349 => "11111111",
	2350 => "11111111",
	2351 => "11111111",
	2352 => "11111111",
	2353 => "11111111",
	2354 => "11111111",
	2355 => "11111111",
	2356 => "11111111",
	2357 => "11111111",
	2358 => "11111111",
	2359 => "11111111",
	2360 => "11111111",
	2361 => "11111111",
	2362 => "11111111",
	2363 => "11111111",
	2364 => "11111111",
	2365 => "11111111",
	2366 => "11111111",
	2367 => "11111111",
	2368 => "11111111",
	2369 => "11111111",
	2370 => "11111111",
	2371 => "11111111",
	2372 => "11111111",
	2373 => "11111111",
	2374 => "11111111",
	2375 => "11111111",
	2376 => "11111111",
	2377 => "11111111",
	2378 => "11111111",
	2379 => "11111111",
	2380 => "11111111",
	2381 => "11111111",
	2382 => "11111111",
	2383 => "11111111",
	2384 => "11111111",
	2385 => "11111111",
	2386 => "11111111",
	2387 => "11111111",
	2388 => "11111111",
	2389 => "11111111",
	2390 => "11111111",
	2391 => "11111111",
	2392 => "11111111",
	2393 => "11111111",
	2394 => "11111111",
	2395 => "11111111",
	2396 => "11111111",
	2397 => "11111111",
	2398 => "11111111",
	2399 => "11111111",
	2400 => "11111111",
	2401 => "11111111",
	2402 => "11111111",
	2403 => "11111111",
	2404 => "11111111",
	2405 => "11111111",
	2406 => "11111111",
	2407 => "11111111",
	2408 => "11111111",
	2409 => "11111111",
	2410 => "11111111",
	2411 => "11111111",
	2412 => "11111111",
	2413 => "11111111",
	2414 => "11111111",
	2415 => "11111111",
	2416 => "11111111",
	2417 => "11111111",
	2418 => "11111111",
	2419 => "11111111",
	2420 => "11111111",
	2421 => "11111111",
	2422 => "11111111",
	2423 => "11111111",
	2432 => "11111111",
	2433 => "11111111",
	2434 => "11111111",
	2435 => "11111111",
	2436 => "11111111",
	2437 => "11111111",
	2438 => "11111111",
	2439 => "11111111",
	2440 => "11111111",
	2441 => "11111111",
	2442 => "11111111",
	2443 => "11111111",
	2444 => "11111111",
	2445 => "11111111",
	2446 => "11111111",
	2447 => "11111111",
	2448 => "11111111",
	2449 => "11111111",
	2450 => "11111111",
	2451 => "11111111",
	2452 => "11111111",
	2453 => "11111111",
	2454 => "11111111",
	2455 => "11111111",
	2456 => "11111111",
	2457 => "11111111",
	2458 => "11111111",
	2459 => "11111111",
	2460 => "11111111",
	2461 => "11111111",
	2462 => "11111111",
	2463 => "11111111",
	2464 => "11111111",
	2465 => "11111111",
	2466 => "11111111",
	2467 => "11111111",
	2468 => "11111111",
	2469 => "11111111",
	2470 => "11111111",
	2471 => "11111111",
	2472 => "11111111",
	2473 => "11111111",
	2474 => "11111111",
	2475 => "11111111",
	2476 => "11111111",
	2477 => "11111111",
	2478 => "11111111",
	2479 => "11111111",
	2480 => "11111111",
	2481 => "11111111",
	2482 => "11111111",
	2483 => "11111111",
	2484 => "11111111",
	2485 => "11111111",
	2486 => "11111111",
	2487 => "11111111",
	2488 => "11111111",
	2489 => "11111111",
	2490 => "11111111",
	2491 => "11111111",
	2492 => "11111111",
	2493 => "11111111",
	2494 => "11111111",
	2495 => "11111111",
	2496 => "11111111",
	2497 => "11111111",
	2498 => "11111111",
	2499 => "11111111",
	2500 => "11111111",
	2501 => "11111111",
	2502 => "11111111",
	2503 => "11111111",
	2504 => "11111111",
	2505 => "11111111",
	2506 => "11111111",
	2507 => "11111111",
	2508 => "11111111",
	2509 => "11111111",
	2510 => "11111111",
	2511 => "11111111",
	2512 => "11111111",
	2513 => "11111111",
	2514 => "11111111",
	2515 => "11111111",
	2516 => "11111111",
	2517 => "11111111",
	2518 => "11111111",
	2519 => "11111111",
	2520 => "11111111",
	2521 => "11111111",
	2522 => "11111111",
	2523 => "11111111",
	2524 => "11111111",
	2525 => "11111111",
	2526 => "11111111",
	2527 => "11111111",
	2528 => "11111111",
	2529 => "11111111",
	2530 => "11111111",
	2531 => "11111111",
	2532 => "11111111",
	2533 => "11111111",
	2534 => "11111111",
	2535 => "11111111",
	2536 => "11111111",
	2537 => "11111111",
	2538 => "11111111",
	2539 => "11111111",
	2540 => "11111111",
	2541 => "11111111",
	2542 => "11111111",
	2543 => "11111111",
	2544 => "11111111",
	2545 => "11111111",
	2546 => "11111111",
	2547 => "11111111",
	2548 => "11111111",
	2549 => "11111111",
	2550 => "11111111",
	2551 => "11111111",
	2560 => "11111111",
	2561 => "11111111",
	2562 => "11111111",
	2563 => "11111111",
	2564 => "11111111",
	2565 => "11111111",
	2566 => "11111111",
	2567 => "11111111",
	2568 => "11111111",
	2569 => "11111111",
	2570 => "11111111",
	2571 => "11111111",
	2572 => "11111111",
	2573 => "11111111",
	2574 => "11111111",
	2575 => "11111111",
	2576 => "11111111",
	2577 => "11111111",
	2578 => "11111111",
	2579 => "11111111",
	2580 => "11111111",
	2581 => "11111111",
	2582 => "11111111",
	2583 => "11111111",
	2584 => "11111111",
	2585 => "11111111",
	2586 => "11111111",
	2587 => "11111111",
	2588 => "11111111",
	2589 => "11111111",
	2590 => "11111111",
	2591 => "11111111",
	2592 => "11111111",
	2593 => "11111111",
	2594 => "11111111",
	2595 => "11111111",
	2596 => "11111111",
	2597 => "11111111",
	2598 => "11111111",
	2599 => "11111111",
	2600 => "11111111",
	2601 => "11111111",
	2602 => "11111111",
	2603 => "11111111",
	2604 => "11111111",
	2605 => "11111111",
	2606 => "11111111",
	2607 => "11111111",
	2608 => "11111111",
	2609 => "11111111",
	2610 => "11111111",
	2611 => "11111111",
	2612 => "11111111",
	2613 => "11111111",
	2614 => "11111111",
	2615 => "11111111",
	2616 => "11111111",
	2617 => "11111111",
	2618 => "11111111",
	2619 => "11111111",
	2620 => "11111111",
	2621 => "11111111",
	2622 => "11111111",
	2623 => "11111111",
	2624 => "11111111",
	2625 => "11111111",
	2626 => "11111111",
	2627 => "11111111",
	2628 => "11111111",
	2629 => "11111111",
	2630 => "11111111",
	2631 => "11111111",
	2632 => "11111111",
	2633 => "11111111",
	2634 => "11111111",
	2635 => "11111111",
	2636 => "11111111",
	2637 => "11111111",
	2638 => "11111111",
	2639 => "11111111",
	2640 => "11111111",
	2641 => "11111111",
	2642 => "11111111",
	2643 => "11111111",
	2644 => "11111111",
	2645 => "11111111",
	2646 => "11111111",
	2647 => "11111111",
	2648 => "11111111",
	2649 => "11111111",
	2650 => "11111111",
	2651 => "11111111",
	2652 => "11111111",
	2653 => "11111111",
	2654 => "11111111",
	2655 => "11111111",
	2656 => "11111111",
	2657 => "11111111",
	2658 => "11111111",
	2659 => "11111111",
	2660 => "11111111",
	2661 => "11111111",
	2662 => "11111111",
	2663 => "11111111",
	2664 => "11111111",
	2665 => "11111111",
	2666 => "11111111",
	2667 => "11111111",
	2668 => "11111111",
	2669 => "11111111",
	2670 => "11111111",
	2671 => "11111111",
	2672 => "11111111",
	2673 => "11111111",
	2674 => "11111111",
	2675 => "11111111",
	2676 => "11111111",
	2677 => "11111111",
	2678 => "11111111",
	2679 => "11111111",
	2688 => "11111111",
	2689 => "11111111",
	2690 => "11111111",
	2691 => "11111111",
	2692 => "11111111",
	2693 => "11111111",
	2694 => "11111111",
	2695 => "11111111",
	2696 => "11111111",
	2697 => "11111111",
	2698 => "11111111",
	2699 => "11111111",
	2700 => "11111111",
	2701 => "11111111",
	2702 => "11111111",
	2703 => "11111111",
	2704 => "11111111",
	2705 => "11111111",
	2706 => "11111111",
	2707 => "11111111",
	2708 => "11111111",
	2709 => "11111111",
	2710 => "11111111",
	2711 => "11111111",
	2712 => "11111111",
	2713 => "11111111",
	2714 => "11111111",
	2715 => "11111111",
	2716 => "11111111",
	2717 => "11111111",
	2718 => "11111111",
	2719 => "11111111",
	2720 => "11111111",
	2721 => "11111111",
	2722 => "11111111",
	2723 => "11111111",
	2724 => "11111111",
	2725 => "11111111",
	2726 => "11111111",
	2727 => "11111111",
	2728 => "11111111",
	2729 => "11111111",
	2730 => "11111111",
	2731 => "11111111",
	2732 => "11111111",
	2733 => "11111111",
	2734 => "11111111",
	2735 => "11111111",
	2736 => "11111111",
	2737 => "11111111",
	2738 => "11111111",
	2739 => "11111111",
	2740 => "11111111",
	2741 => "11111111",
	2742 => "11111111",
	2743 => "11111111",
	2744 => "11111111",
	2745 => "11111111",
	2746 => "11111111",
	2747 => "11111111",
	2748 => "11111111",
	2749 => "11111111",
	2750 => "11111111",
	2751 => "11111111",
	2752 => "11111111",
	2753 => "11111111",
	2754 => "11111111",
	2755 => "11111111",
	2756 => "11111111",
	2757 => "11111111",
	2758 => "11111111",
	2759 => "11111111",
	2760 => "11111111",
	2761 => "11111111",
	2762 => "11111111",
	2763 => "11111111",
	2764 => "11111111",
	2765 => "11111111",
	2766 => "11111111",
	2767 => "11111111",
	2768 => "11111111",
	2769 => "11111111",
	2770 => "11111111",
	2771 => "11111111",
	2772 => "11111111",
	2773 => "11111111",
	2774 => "11111111",
	2775 => "11111111",
	2776 => "11111111",
	2777 => "11111111",
	2778 => "11111111",
	2779 => "11111111",
	2780 => "11111111",
	2781 => "11111111",
	2782 => "11111111",
	2783 => "11111111",
	2784 => "11111111",
	2785 => "11111111",
	2786 => "11111111",
	2787 => "11111111",
	2788 => "11111111",
	2789 => "11111111",
	2790 => "11111111",
	2791 => "11111111",
	2792 => "11111111",
	2793 => "11111111",
	2794 => "11111111",
	2795 => "11111111",
	2796 => "11111111",
	2797 => "11111111",
	2798 => "11111111",
	2799 => "11111111",
	2800 => "11111111",
	2801 => "11111111",
	2802 => "11111111",
	2803 => "11111111",
	2804 => "11111111",
	2805 => "11111111",
	2806 => "11111111",
	2807 => "11111111",
	2816 => "11111111",
	2817 => "11111111",
	2818 => "11111111",
	2819 => "11111111",
	2820 => "11111111",
	2821 => "11111111",
	2822 => "11111111",
	2823 => "11111111",
	2824 => "11111111",
	2825 => "11111111",
	2826 => "11111111",
	2827 => "11111111",
	2828 => "11111111",
	2829 => "11111111",
	2830 => "11111111",
	2831 => "11111111",
	2832 => "11111111",
	2833 => "11111111",
	2834 => "11111111",
	2835 => "11111111",
	2836 => "11111111",
	2837 => "11111111",
	2838 => "11111111",
	2839 => "11111111",
	2840 => "11111111",
	2841 => "11111111",
	2842 => "11111111",
	2843 => "11111111",
	2844 => "11111111",
	2845 => "11111111",
	2846 => "11111111",
	2847 => "11111111",
	2848 => "11111111",
	2849 => "11111111",
	2850 => "11111111",
	2851 => "11111111",
	2852 => "11111111",
	2853 => "11111111",
	2854 => "11111111",
	2855 => "11111111",
	2856 => "11111111",
	2857 => "11111111",
	2858 => "11111111",
	2859 => "11111111",
	2860 => "11111111",
	2861 => "11111111",
	2862 => "11111111",
	2863 => "11111111",
	2864 => "11111111",
	2865 => "11111111",
	2866 => "11111111",
	2867 => "11111111",
	2868 => "11111111",
	2869 => "11111111",
	2870 => "11111111",
	2871 => "11111111",
	2872 => "11111111",
	2873 => "11111111",
	2874 => "11111111",
	2875 => "11111111",
	2876 => "11111111",
	2877 => "11111111",
	2878 => "11111111",
	2879 => "11111111",
	2880 => "11111111",
	2881 => "11111111",
	2882 => "11111111",
	2883 => "11111111",
	2884 => "11111111",
	2885 => "11111111",
	2886 => "11111111",
	2887 => "11111111",
	2888 => "11111111",
	2889 => "11111111",
	2890 => "11111111",
	2891 => "11111111",
	2892 => "11111111",
	2893 => "11111111",
	2894 => "11111111",
	2895 => "11111111",
	2896 => "11111111",
	2897 => "11111111",
	2898 => "11111111",
	2899 => "11111111",
	2900 => "11111111",
	2901 => "11111111",
	2902 => "11111111",
	2903 => "11111111",
	2904 => "11111111",
	2905 => "11111111",
	2906 => "11111111",
	2907 => "11111111",
	2908 => "11111111",
	2909 => "11111111",
	2910 => "11111111",
	2911 => "11111111",
	2912 => "11111111",
	2913 => "11111111",
	2914 => "11111111",
	2915 => "11111111",
	2916 => "11111111",
	2917 => "11111111",
	2918 => "11111111",
	2919 => "11111111",
	2920 => "11111111",
	2921 => "11111111",
	2922 => "11111111",
	2923 => "11111111",
	2924 => "11111111",
	2925 => "11111111",
	2926 => "11111111",
	2927 => "11111111",
	2928 => "11111111",
	2929 => "11111111",
	2930 => "11111111",
	2931 => "11111111",
	2932 => "11111111",
	2933 => "11111111",
	2934 => "11111111",
	2935 => "11111111",
	2944 => "11111111",
	2945 => "11111111",
	2946 => "11111111",
	2947 => "11111111",
	2948 => "11111111",
	2949 => "11111111",
	2950 => "11111111",
	2951 => "11111111",
	2952 => "11111111",
	2953 => "11111111",
	2954 => "11111111",
	2955 => "11111111",
	2956 => "11111111",
	2957 => "11111111",
	2958 => "11111111",
	2959 => "11111111",
	2960 => "11111111",
	2961 => "11111111",
	2962 => "11111111",
	2963 => "11111111",
	2964 => "11111111",
	2965 => "11111111",
	2966 => "11111111",
	2967 => "11111111",
	2968 => "11111111",
	2969 => "11111111",
	2970 => "11111111",
	2971 => "11111111",
	2972 => "11111111",
	2973 => "11111111",
	2974 => "11111111",
	2975 => "11111111",
	2976 => "11111111",
	2977 => "11111111",
	2978 => "11111111",
	2979 => "11111111",
	2980 => "11111111",
	2981 => "11111111",
	2982 => "11111111",
	2983 => "11111111",
	2984 => "11111111",
	2985 => "11111111",
	2986 => "11111111",
	2987 => "11111111",
	2988 => "11111111",
	2989 => "11111111",
	2990 => "11111111",
	2991 => "11111111",
	2992 => "11111111",
	2993 => "11111111",
	2994 => "11111111",
	2995 => "11111111",
	2996 => "11111111",
	2997 => "11111111",
	2998 => "11111111",
	2999 => "11111111",
	3000 => "11111111",
	3001 => "11111111",
	3002 => "11111111",
	3003 => "11111111",
	3004 => "11111111",
	3005 => "11111111",
	3006 => "11111111",
	3007 => "11111111",
	3008 => "11111111",
	3009 => "11111111",
	3010 => "11111111",
	3011 => "11111111",
	3012 => "11111111",
	3013 => "11111111",
	3014 => "11111111",
	3015 => "11111111",
	3016 => "11111111",
	3017 => "11111111",
	3018 => "11111111",
	3019 => "11111111",
	3020 => "11111111",
	3021 => "11111111",
	3022 => "11111111",
	3023 => "11111111",
	3024 => "11111111",
	3025 => "11111111",
	3026 => "11111111",
	3027 => "11111111",
	3028 => "11111111",
	3029 => "11111111",
	3030 => "11111111",
	3031 => "11111111",
	3032 => "11111111",
	3033 => "11111111",
	3034 => "11111111",
	3035 => "11111111",
	3036 => "11111111",
	3037 => "11111111",
	3038 => "11111111",
	3039 => "11111111",
	3040 => "11111111",
	3041 => "11111111",
	3042 => "11111111",
	3043 => "11111111",
	3044 => "11111111",
	3045 => "11111111",
	3046 => "11111111",
	3047 => "11111111",
	3048 => "11111111",
	3049 => "11111111",
	3050 => "11111111",
	3051 => "11111111",
	3052 => "11111111",
	3053 => "11111111",
	3054 => "11111111",
	3055 => "11111111",
	3056 => "11111111",
	3057 => "11111111",
	3058 => "11111111",
	3059 => "11111111",
	3060 => "11111111",
	3061 => "11111111",
	3062 => "11111111",
	3063 => "11111111",
	3072 => "11111111",
	3073 => "11111111",
	3074 => "11111111",
	3075 => "11111111",
	3076 => "11111111",
	3077 => "11111111",
	3078 => "11111111",
	3079 => "11111111",
	3080 => "11111111",
	3081 => "11111111",
	3082 => "11111111",
	3083 => "11111111",
	3084 => "11111111",
	3085 => "11111111",
	3086 => "11111111",
	3087 => "11111111",
	3088 => "11111111",
	3089 => "11111111",
	3090 => "11111111",
	3091 => "11111111",
	3092 => "11111111",
	3093 => "11111111",
	3094 => "11111111",
	3095 => "11111111",
	3096 => "11111111",
	3097 => "11111111",
	3098 => "11111111",
	3099 => "11111111",
	3100 => "11111111",
	3101 => "11111111",
	3102 => "11111111",
	3103 => "11111111",
	3104 => "11111111",
	3105 => "11111111",
	3106 => "11111111",
	3107 => "11111111",
	3108 => "11111111",
	3109 => "11111111",
	3110 => "11111111",
	3111 => "11111111",
	3112 => "11111111",
	3113 => "11111111",
	3114 => "11111111",
	3115 => "11111111",
	3116 => "11111111",
	3117 => "11111111",
	3118 => "11111111",
	3119 => "11111111",
	3120 => "11111111",
	3121 => "11111111",
	3122 => "11111111",
	3123 => "11111111",
	3124 => "11111111",
	3125 => "11111111",
	3126 => "11111111",
	3127 => "11111111",
	3128 => "11111111",
	3129 => "11111111",
	3130 => "11111111",
	3131 => "11111111",
	3132 => "11111111",
	3133 => "11111111",
	3134 => "11111111",
	3135 => "11111111",
	3136 => "11111111",
	3137 => "11111111",
	3138 => "11111111",
	3139 => "11111111",
	3140 => "11111111",
	3141 => "11111111",
	3142 => "11111111",
	3143 => "11111111",
	3144 => "11111111",
	3145 => "11111111",
	3146 => "11111111",
	3147 => "11111111",
	3148 => "11111111",
	3149 => "11111111",
	3150 => "11111111",
	3151 => "11111111",
	3152 => "11111111",
	3153 => "11111111",
	3154 => "11111111",
	3155 => "11111111",
	3156 => "11111111",
	3157 => "11111111",
	3158 => "11111111",
	3159 => "11111111",
	3160 => "11111111",
	3161 => "11111111",
	3162 => "11111111",
	3163 => "11111111",
	3164 => "11111111",
	3165 => "11111111",
	3166 => "11111111",
	3167 => "11111111",
	3168 => "11111111",
	3169 => "11111111",
	3170 => "11111111",
	3171 => "11111111",
	3172 => "11111111",
	3173 => "11111111",
	3174 => "11111111",
	3175 => "11111111",
	3176 => "11111111",
	3177 => "11111111",
	3178 => "11111111",
	3179 => "11111111",
	3180 => "11111111",
	3181 => "11111111",
	3182 => "11111111",
	3183 => "11111111",
	3184 => "11111111",
	3185 => "11111111",
	3186 => "11111111",
	3187 => "11111111",
	3188 => "11111111",
	3189 => "11111111",
	3190 => "11111111",
	3191 => "11111111",
	3200 => "11111111",
	3201 => "11111111",
	3202 => "11111111",
	3203 => "11111111",
	3204 => "11111111",
	3205 => "11111111",
	3206 => "11111111",
	3207 => "11111111",
	3208 => "11111111",
	3209 => "11111111",
	3210 => "11111111",
	3211 => "11111111",
	3212 => "11111111",
	3213 => "11111111",
	3214 => "11111111",
	3215 => "11111111",
	3216 => "11111111",
	3217 => "11111111",
	3218 => "11111111",
	3219 => "11111111",
	3220 => "11111111",
	3221 => "11111111",
	3222 => "11111111",
	3223 => "11111111",
	3224 => "11111111",
	3225 => "11111111",
	3226 => "11111111",
	3227 => "11111111",
	3228 => "11111111",
	3229 => "11111111",
	3230 => "11111111",
	3231 => "11111111",
	3232 => "11111111",
	3233 => "11111111",
	3234 => "11111111",
	3235 => "11111111",
	3236 => "11111111",
	3237 => "11111111",
	3238 => "11111111",
	3239 => "11111111",
	3240 => "11111111",
	3241 => "11111111",
	3242 => "11111111",
	3243 => "11111111",
	3244 => "11111111",
	3245 => "11111111",
	3246 => "11111111",
	3247 => "11111111",
	3248 => "11111111",
	3249 => "11111111",
	3250 => "11111111",
	3251 => "11111111",
	3252 => "11111111",
	3253 => "11111111",
	3254 => "11111111",
	3255 => "11111111",
	3256 => "11111111",
	3257 => "11111111",
	3258 => "11111111",
	3259 => "11111111",
	3260 => "11111111",
	3261 => "11111111",
	3262 => "11111111",
	3263 => "11111111",
	3264 => "11111111",
	3265 => "11111111",
	3266 => "11111111",
	3267 => "11111111",
	3268 => "11111111",
	3269 => "11111111",
	3270 => "11111111",
	3271 => "11111111",
	3272 => "11111111",
	3273 => "11111111",
	3274 => "11111111",
	3275 => "11111111",
	3276 => "11111111",
	3277 => "11111111",
	3278 => "11111111",
	3279 => "11111111",
	3280 => "11111111",
	3281 => "11111111",
	3282 => "11111111",
	3283 => "11111111",
	3284 => "11111111",
	3285 => "11111111",
	3286 => "11111111",
	3287 => "11111111",
	3288 => "11111111",
	3289 => "11111111",
	3290 => "11111111",
	3291 => "11111111",
	3292 => "11111111",
	3293 => "11111111",
	3294 => "11111111",
	3295 => "11111111",
	3296 => "11111111",
	3297 => "11111111",
	3298 => "11111111",
	3299 => "11111111",
	3300 => "11111111",
	3301 => "11111111",
	3302 => "11111111",
	3303 => "11111111",
	3304 => "11111111",
	3305 => "11111111",
	3306 => "11111111",
	3307 => "11111111",
	3308 => "11111111",
	3309 => "11111111",
	3310 => "11111111",
	3311 => "11111111",
	3312 => "11111111",
	3313 => "11111111",
	3314 => "11111111",
	3315 => "11111111",
	3316 => "11111111",
	3317 => "11111111",
	3318 => "11111111",
	3319 => "11111111",
	3328 => "11111111",
	3329 => "11111111",
	3330 => "11111111",
	3331 => "11111111",
	3332 => "11111111",
	3333 => "11111111",
	3334 => "11111111",
	3335 => "11111111",
	3336 => "11111111",
	3337 => "11111111",
	3338 => "11111111",
	3339 => "11111111",
	3340 => "11111111",
	3341 => "11111111",
	3342 => "11111111",
	3343 => "11111111",
	3344 => "11111111",
	3345 => "11111111",
	3346 => "11111111",
	3347 => "11111111",
	3348 => "11111111",
	3349 => "11111111",
	3350 => "11111111",
	3351 => "11111111",
	3352 => "11111111",
	3353 => "11111111",
	3354 => "11111111",
	3355 => "11111111",
	3356 => "11111111",
	3357 => "11111111",
	3358 => "11111111",
	3359 => "11111111",
	3360 => "11111111",
	3361 => "11111111",
	3362 => "11111111",
	3363 => "11111111",
	3364 => "11111111",
	3365 => "11111111",
	3366 => "11111111",
	3367 => "11111111",
	3368 => "11111111",
	3369 => "11111111",
	3370 => "11111111",
	3371 => "11111111",
	3372 => "11111111",
	3373 => "11111111",
	3374 => "11111111",
	3375 => "11111111",
	3376 => "11111111",
	3377 => "11111111",
	3378 => "11111111",
	3379 => "11111111",
	3380 => "11111111",
	3381 => "11111111",
	3382 => "11111111",
	3383 => "11111111",
	3384 => "11111111",
	3385 => "11111111",
	3386 => "11111111",
	3387 => "11111111",
	3388 => "11111111",
	3389 => "11111111",
	3390 => "11111111",
	3391 => "11111111",
	3392 => "11111111",
	3393 => "11111111",
	3394 => "11111111",
	3395 => "11111111",
	3396 => "11111111",
	3397 => "11111111",
	3398 => "11111111",
	3399 => "11111111",
	3400 => "11111111",
	3401 => "11111111",
	3402 => "11111111",
	3403 => "11111111",
	3404 => "11111111",
	3405 => "11111111",
	3406 => "11111111",
	3407 => "11111111",
	3408 => "11111111",
	3409 => "11111111",
	3410 => "11111111",
	3411 => "11111111",
	3412 => "11111111",
	3413 => "11111111",
	3414 => "11111111",
	3415 => "11111111",
	3416 => "11111111",
	3417 => "11111111",
	3418 => "11111111",
	3419 => "11111111",
	3420 => "11111111",
	3421 => "11111111",
	3422 => "11111111",
	3423 => "11111111",
	3424 => "11111111",
	3425 => "11111111",
	3426 => "11111111",
	3427 => "11111111",
	3428 => "11111111",
	3429 => "11111111",
	3430 => "11111111",
	3431 => "11111111",
	3432 => "11111111",
	3433 => "11111111",
	3434 => "11111111",
	3435 => "11111111",
	3436 => "11111111",
	3437 => "11111111",
	3438 => "11111111",
	3439 => "11111111",
	3440 => "11111111",
	3441 => "11111111",
	3442 => "11111111",
	3443 => "11111111",
	3444 => "11111111",
	3445 => "11111111",
	3446 => "11111111",
	3447 => "11111111",
	3456 => "11111111",
	3457 => "11111111",
	3458 => "11111111",
	3459 => "11111111",
	3460 => "11111111",
	3461 => "11111111",
	3462 => "11111111",
	3463 => "11111111",
	3464 => "11111111",
	3465 => "11111111",
	3466 => "11111111",
	3467 => "11111111",
	3468 => "11111111",
	3469 => "11111111",
	3470 => "11111111",
	3471 => "11111111",
	3472 => "11111111",
	3473 => "11111111",
	3474 => "11111111",
	3475 => "11111111",
	3476 => "11111111",
	3477 => "11111111",
	3478 => "11111111",
	3479 => "11111111",
	3480 => "11111111",
	3481 => "11111111",
	3482 => "11111111",
	3483 => "11111111",
	3484 => "11111111",
	3485 => "11111111",
	3486 => "11111111",
	3487 => "11111111",
	3488 => "11111111",
	3489 => "11111111",
	3490 => "11111111",
	3491 => "11111111",
	3492 => "11111111",
	3493 => "11111111",
	3494 => "11111111",
	3495 => "11111111",
	3496 => "11111111",
	3497 => "11111111",
	3498 => "11111111",
	3499 => "11111111",
	3500 => "11111111",
	3501 => "11111111",
	3502 => "11111111",
	3503 => "11111111",
	3504 => "11111111",
	3505 => "11111111",
	3506 => "11111111",
	3507 => "11111111",
	3508 => "11111111",
	3509 => "11111111",
	3510 => "11111111",
	3511 => "11111111",
	3512 => "11111111",
	3513 => "11111111",
	3514 => "11111111",
	3515 => "11111111",
	3516 => "11111111",
	3517 => "11111111",
	3518 => "11111111",
	3519 => "11111111",
	3520 => "11111111",
	3521 => "11111111",
	3522 => "11111111",
	3523 => "11111111",
	3524 => "11111111",
	3525 => "11111111",
	3526 => "11111111",
	3527 => "11111111",
	3528 => "11111111",
	3529 => "11111111",
	3530 => "11111111",
	3531 => "11111111",
	3532 => "11111111",
	3533 => "11111111",
	3534 => "11111111",
	3535 => "11111111",
	3536 => "11111111",
	3537 => "11111111",
	3538 => "11111111",
	3539 => "11111111",
	3540 => "11111111",
	3541 => "11111111",
	3542 => "11111111",
	3543 => "11111111",
	3544 => "11111111",
	3545 => "11111111",
	3546 => "11111111",
	3547 => "11111111",
	3548 => "11111111",
	3549 => "11111111",
	3550 => "11111111",
	3551 => "11111111",
	3552 => "11111111",
	3553 => "11111111",
	3554 => "11111111",
	3555 => "11111111",
	3556 => "11111111",
	3557 => "11111111",
	3558 => "11111111",
	3559 => "11111111",
	3560 => "11111111",
	3561 => "11111111",
	3562 => "11111111",
	3563 => "11111111",
	3564 => "11111111",
	3565 => "11111111",
	3566 => "11111111",
	3567 => "11111111",
	3568 => "11111111",
	3569 => "11111111",
	3570 => "11111111",
	3571 => "11111111",
	3572 => "11111111",
	3573 => "11111111",
	3574 => "11111111",
	3575 => "11111111",
	3584 => "11111111",
	3585 => "11111111",
	3586 => "11111111",
	3587 => "11111111",
	3588 => "11111111",
	3589 => "11111111",
	3590 => "11111111",
	3591 => "11111111",
	3592 => "11111111",
	3593 => "11111111",
	3594 => "11111111",
	3595 => "11111111",
	3596 => "11111111",
	3597 => "11111111",
	3598 => "11111111",
	3599 => "11111111",
	3600 => "11111111",
	3601 => "11111111",
	3602 => "11111111",
	3603 => "11111111",
	3604 => "11111111",
	3605 => "11111111",
	3606 => "11111111",
	3607 => "11111111",
	3608 => "11111111",
	3609 => "11111111",
	3610 => "11111111",
	3611 => "11111111",
	3612 => "11111111",
	3613 => "11111111",
	3614 => "11111111",
	3615 => "11111111",
	3616 => "11111111",
	3617 => "11111111",
	3618 => "11111111",
	3619 => "11111111",
	3620 => "11111111",
	3621 => "11111111",
	3622 => "11111111",
	3623 => "11111111",
	3624 => "11111111",
	3625 => "11111111",
	3626 => "11111111",
	3627 => "11111111",
	3628 => "11111111",
	3629 => "11111111",
	3630 => "11111111",
	3631 => "11111111",
	3632 => "11111111",
	3633 => "11111111",
	3634 => "11111111",
	3635 => "11111111",
	3636 => "11111111",
	3637 => "11111111",
	3638 => "11111111",
	3639 => "11111111",
	3640 => "11111111",
	3641 => "11111111",
	3642 => "11111111",
	3643 => "11111111",
	3644 => "11111111",
	3645 => "11111111",
	3646 => "11111111",
	3647 => "11111111",
	3648 => "11111111",
	3649 => "11111111",
	3650 => "11111111",
	3651 => "11111111",
	3652 => "11111111",
	3653 => "11111111",
	3654 => "11111111",
	3655 => "11111111",
	3656 => "11111111",
	3657 => "11111111",
	3658 => "11111111",
	3659 => "11111111",
	3660 => "11111111",
	3661 => "11111111",
	3662 => "11111111",
	3663 => "11111111",
	3664 => "11111111",
	3665 => "11111111",
	3666 => "11111111",
	3667 => "11111111",
	3668 => "11111111",
	3669 => "11111111",
	3670 => "11111111",
	3671 => "11111111",
	3672 => "11111111",
	3673 => "11111111",
	3674 => "11111111",
	3675 => "11111111",
	3676 => "11111111",
	3677 => "11111111",
	3678 => "11111111",
	3679 => "11111111",
	3680 => "11111111",
	3681 => "11111111",
	3682 => "11111111",
	3683 => "11111111",
	3684 => "11111111",
	3685 => "11111111",
	3686 => "11111111",
	3687 => "11111111",
	3688 => "11111111",
	3689 => "11111111",
	3690 => "11111111",
	3691 => "11111111",
	3692 => "11111111",
	3693 => "11111111",
	3694 => "11111111",
	3695 => "11111111",
	3696 => "11111111",
	3697 => "11111111",
	3698 => "11111111",
	3699 => "11111111",
	3700 => "11111111",
	3701 => "11111111",
	3702 => "11111111",
	3703 => "11111111",
	3712 => "11111111",
	3713 => "11111111",
	3714 => "11111111",
	3715 => "11111111",
	3716 => "11111111",
	3717 => "11111111",
	3718 => "11111111",
	3719 => "11111111",
	3720 => "11111111",
	3721 => "11111111",
	3722 => "11111111",
	3723 => "11111111",
	3724 => "11111111",
	3725 => "11111111",
	3726 => "11111111",
	3727 => "11111111",
	3728 => "11111111",
	3729 => "11111111",
	3730 => "11111111",
	3731 => "11111111",
	3732 => "11111111",
	3733 => "11111111",
	3734 => "11111111",
	3735 => "11111111",
	3736 => "11111111",
	3737 => "11111111",
	3738 => "11111111",
	3739 => "11111111",
	3740 => "11111111",
	3741 => "11111111",
	3742 => "11111111",
	3743 => "11111111",
	3744 => "11111111",
	3745 => "11111111",
	3746 => "11111111",
	3747 => "11111111",
	3748 => "11111111",
	3749 => "11111111",
	3750 => "11111111",
	3751 => "11111111",
	3752 => "11111111",
	3753 => "11111111",
	3754 => "11111111",
	3755 => "11111111",
	3756 => "11111111",
	3757 => "11111111",
	3758 => "11111111",
	3759 => "11111111",
	3760 => "11111111",
	3761 => "11111111",
	3762 => "11111111",
	3763 => "11111111",
	3764 => "11111111",
	3765 => "11111111",
	3766 => "11111111",
	3767 => "11111111",
	3768 => "11111111",
	3769 => "11111111",
	3770 => "11111111",
	3771 => "11111111",
	3772 => "11111111",
	3773 => "11111111",
	3774 => "11111111",
	3775 => "11111111",
	3776 => "11111111",
	3777 => "11111111",
	3778 => "11111111",
	3779 => "11111111",
	3780 => "11111111",
	3781 => "11111111",
	3782 => "11111111",
	3783 => "11111111",
	3784 => "11111111",
	3785 => "11111111",
	3786 => "11111111",
	3787 => "11111111",
	3788 => "11111111",
	3789 => "11111111",
	3790 => "11111111",
	3791 => "11111111",
	3792 => "11111111",
	3793 => "11111111",
	3794 => "11111111",
	3795 => "11111111",
	3796 => "11111111",
	3797 => "11111111",
	3798 => "11111111",
	3799 => "11111111",
	3800 => "11111111",
	3801 => "11111111",
	3802 => "11111111",
	3803 => "11111111",
	3804 => "11111111",
	3805 => "11111111",
	3806 => "11111111",
	3807 => "11111111",
	3808 => "11111111",
	3809 => "11111111",
	3810 => "11111111",
	3811 => "11111111",
	3812 => "11111111",
	3813 => "11111111",
	3814 => "11111111",
	3815 => "11111111",
	3816 => "11111111",
	3817 => "11111111",
	3818 => "11111111",
	3819 => "11111111",
	3820 => "11111111",
	3821 => "11111111",
	3822 => "11111111",
	3823 => "11111111",
	3824 => "11111111",
	3825 => "11111111",
	3826 => "11111111",
	3827 => "11111111",
	3828 => "11111111",
	3829 => "11111111",
	3830 => "11111111",
	3831 => "11111111",
	3840 => "11111111",
	3841 => "11111111",
	3842 => "11111111",
	3843 => "11111111",
	3844 => "11111111",
	3845 => "11111111",
	3846 => "11111111",
	3847 => "11111111",
	3848 => "11111111",
	3849 => "11111111",
	3850 => "11111111",
	3851 => "11111111",
	3852 => "11111111",
	3853 => "11111111",
	3854 => "11111111",
	3855 => "11111111",
	3856 => "11111111",
	3857 => "11111111",
	3858 => "11111111",
	3859 => "11111111",
	3860 => "11111111",
	3861 => "11111111",
	3862 => "11111111",
	3863 => "11111111",
	3864 => "11111111",
	3865 => "11111111",
	3866 => "11111111",
	3867 => "11111111",
	3868 => "11111111",
	3869 => "11111111",
	3870 => "11111111",
	3871 => "11111111",
	3872 => "11111111",
	3873 => "11111111",
	3874 => "11111111",
	3875 => "11111111",
	3876 => "11111111",
	3877 => "11111111",
	3878 => "11111111",
	3879 => "11111111",
	3880 => "11111111",
	3881 => "11111111",
	3882 => "11111111",
	3883 => "11111111",
	3884 => "11111111",
	3885 => "11111111",
	3886 => "11111111",
	3887 => "11111111",
	3888 => "11111111",
	3889 => "11111111",
	3890 => "11111111",
	3891 => "11111111",
	3892 => "11111111",
	3893 => "11111111",
	3894 => "11111111",
	3895 => "11111111",
	3896 => "11111111",
	3897 => "11111111",
	3898 => "11111111",
	3899 => "11111111",
	3900 => "11111111",
	3901 => "11111111",
	3902 => "11111111",
	3903 => "11111111",
	3904 => "11111111",
	3905 => "11111111",
	3906 => "11111111",
	3907 => "11111111",
	3908 => "11111111",
	3909 => "11111111",
	3910 => "11111111",
	3911 => "11111111",
	3912 => "11111111",
	3913 => "11111111",
	3914 => "11111111",
	3915 => "11111111",
	3916 => "11111111",
	3917 => "11111111",
	3918 => "11111111",
	3919 => "11111111",
	3920 => "11111111",
	3921 => "11111111",
	3922 => "11111111",
	3923 => "11111111",
	3924 => "11111111",
	3925 => "11111111",
	3926 => "11111111",
	3927 => "11111111",
	3928 => "11111111",
	3929 => "11111111",
	3930 => "11111111",
	3931 => "11111111",
	3932 => "11111111",
	3933 => "11111111",
	3934 => "11111111",
	3935 => "11111111",
	3936 => "11111111",
	3937 => "11111111",
	3938 => "11111111",
	3939 => "11111111",
	3940 => "11111111",
	3941 => "11111111",
	3942 => "11111111",
	3943 => "11111111",
	3944 => "11111111",
	3945 => "11111111",
	3946 => "11111111",
	3947 => "11111111",
	3948 => "11111111",
	3949 => "11111111",
	3950 => "11111111",
	3951 => "11111111",
	3952 => "11111111",
	3953 => "11111111",
	3954 => "11111111",
	3955 => "11111111",
	3956 => "11111111",
	3957 => "11111111",
	3958 => "11111111",
	3959 => "11111111",
	3968 => "11111111",
	3969 => "11111111",
	3970 => "11111111",
	3971 => "11111111",
	3972 => "11111111",
	3973 => "11111111",
	3974 => "11111111",
	3975 => "11111111",
	3976 => "11111111",
	3977 => "11111111",
	3978 => "11111111",
	3979 => "11111111",
	3980 => "11111111",
	3981 => "11111111",
	3982 => "11111111",
	3983 => "11111111",
	3984 => "11111111",
	3985 => "11111111",
	3986 => "11111111",
	3987 => "11111111",
	3988 => "11111111",
	3989 => "11111111",
	3990 => "11111111",
	3991 => "11111111",
	3992 => "11111111",
	3993 => "11111111",
	3994 => "11111111",
	3995 => "11111111",
	3996 => "11111111",
	3997 => "11111111",
	3998 => "11111111",
	3999 => "11111111",
	4000 => "11111111",
	4001 => "11111111",
	4002 => "11111111",
	4003 => "11111111",
	4004 => "11111111",
	4005 => "11111111",
	4006 => "11111111",
	4007 => "11111111",
	4008 => "11111111",
	4009 => "11111111",
	4010 => "11111111",
	4011 => "11111111",
	4012 => "11111111",
	4013 => "11111111",
	4014 => "11111111",
	4015 => "11111111",
	4016 => "11111111",
	4017 => "11111111",
	4018 => "11111111",
	4019 => "11111111",
	4020 => "11111111",
	4021 => "11111111",
	4022 => "11111111",
	4023 => "11111111",
	4024 => "11111111",
	4025 => "11111111",
	4026 => "11111111",
	4027 => "11111111",
	4028 => "11111111",
	4029 => "11111111",
	4030 => "11111111",
	4031 => "11111111",
	4032 => "11111111",
	4033 => "11111111",
	4034 => "11111111",
	4035 => "11111111",
	4036 => "11111111",
	4037 => "11111111",
	4038 => "11111111",
	4039 => "11111111",
	4040 => "11111111",
	4041 => "11111111",
	4042 => "11111111",
	4043 => "11111111",
	4044 => "11111111",
	4045 => "11111111",
	4046 => "11111111",
	4047 => "11111111",
	4048 => "11111111",
	4049 => "11111111",
	4050 => "11111111",
	4051 => "11111111",
	4052 => "11111111",
	4053 => "11111111",
	4054 => "11111111",
	4055 => "11111111",
	4056 => "11111111",
	4057 => "11111111",
	4058 => "11111111",
	4059 => "11111111",
	4060 => "11111111",
	4061 => "11111111",
	4062 => "11111111",
	4063 => "11111111",
	4064 => "11111111",
	4065 => "11111111",
	4066 => "11111111",
	4067 => "11111111",
	4068 => "11111111",
	4069 => "11111111",
	4070 => "11111111",
	4071 => "11111111",
	4072 => "11111111",
	4073 => "11111111",
	4074 => "11111111",
	4075 => "11111111",
	4076 => "11111111",
	4077 => "11111111",
	4078 => "11111111",
	4079 => "11111111",
	4080 => "11111111",
	4081 => "11111111",
	4082 => "11111111",
	4083 => "11111111",
	4084 => "11111111",
	4085 => "11111111",
	4086 => "11111111",
	4087 => "11111111",
	4096 => "11111111",
	4097 => "11111111",
	4098 => "11111111",
	4099 => "11111111",
	4100 => "11111111",
	4101 => "11111111",
	4102 => "11111111",
	4103 => "11111111",
	4104 => "11111111",
	4105 => "11111111",
	4106 => "11111111",
	4107 => "11111111",
	4108 => "11111111",
	4109 => "11111111",
	4110 => "11111111",
	4111 => "11111111",
	4112 => "11111111",
	4113 => "11111111",
	4114 => "11111111",
	4115 => "11111111",
	4116 => "11111111",
	4117 => "11111111",
	4118 => "11111111",
	4119 => "11111111",
	4120 => "11111111",
	4121 => "11111111",
	4122 => "11111111",
	4123 => "11111111",
	4124 => "11111111",
	4125 => "11111111",
	4126 => "11111111",
	4127 => "11111111",
	4128 => "11111111",
	4129 => "11111111",
	4130 => "11111111",
	4131 => "11111111",
	4132 => "11111111",
	4133 => "11111111",
	4134 => "11111111",
	4135 => "11111111",
	4136 => "11111111",
	4137 => "11111111",
	4138 => "11111111",
	4139 => "11111111",
	4140 => "11111111",
	4141 => "11111111",
	4142 => "11111111",
	4143 => "11111111",
	4144 => "11111111",
	4145 => "11111111",
	4146 => "11111111",
	4147 => "11111111",
	4148 => "11111111",
	4149 => "11111111",
	4150 => "11111111",
	4151 => "11111111",
	4152 => "11111111",
	4153 => "11111111",
	4154 => "11111111",
	4155 => "11111111",
	4156 => "11111111",
	4157 => "11111111",
	4158 => "11111111",
	4159 => "11111111",
	4160 => "11111111",
	4161 => "11111111",
	4162 => "11111111",
	4163 => "11111111",
	4164 => "11111111",
	4165 => "11111111",
	4166 => "11111111",
	4167 => "11111111",
	4168 => "11111111",
	4169 => "11111111",
	4170 => "11111111",
	4171 => "11111111",
	4172 => "11111111",
	4173 => "11111111",
	4174 => "11111111",
	4175 => "11111111",
	4176 => "11111111",
	4177 => "11111111",
	4178 => "11111111",
	4179 => "11111111",
	4180 => "11111111",
	4181 => "11111111",
	4182 => "11111111",
	4183 => "11111111",
	4184 => "11111111",
	4185 => "11111111",
	4186 => "11111111",
	4187 => "11111111",
	4188 => "11111111",
	4189 => "11111111",
	4190 => "11111111",
	4191 => "11111111",
	4192 => "11111111",
	4193 => "11111111",
	4194 => "11111111",
	4195 => "11111111",
	4196 => "11111111",
	4197 => "11111111",
	4198 => "11111111",
	4199 => "11111111",
	4200 => "11111111",
	4201 => "11111111",
	4202 => "11111111",
	4203 => "11111111",
	4204 => "11111111",
	4205 => "11111111",
	4206 => "11111111",
	4207 => "11111111",
	4208 => "11111111",
	4209 => "11111111",
	4210 => "11111111",
	4211 => "11111111",
	4212 => "11111111",
	4213 => "11111111",
	4214 => "11111111",
	4215 => "11111111",
	4224 => "11111111",
	4225 => "11111111",
	4226 => "11111111",
	4227 => "11111111",
	4228 => "11111111",
	4229 => "11111111",
	4230 => "11111111",
	4231 => "11111111",
	4232 => "11111111",
	4233 => "11111111",
	4234 => "11111111",
	4235 => "11111111",
	4236 => "11111111",
	4237 => "11111111",
	4238 => "11111111",
	4239 => "11111111",
	4240 => "11111111",
	4241 => "11111111",
	4242 => "11111111",
	4243 => "11111111",
	4244 => "11111111",
	4245 => "11111111",
	4246 => "11111111",
	4247 => "11111111",
	4248 => "11111111",
	4249 => "11111111",
	4250 => "11111111",
	4251 => "11111111",
	4252 => "11111111",
	4253 => "11111111",
	4254 => "11111111",
	4255 => "11111111",
	4256 => "11111111",
	4257 => "11111111",
	4258 => "11111111",
	4259 => "11111111",
	4260 => "11111111",
	4261 => "11111111",
	4262 => "11111111",
	4263 => "11111111",
	4264 => "11111111",
	4265 => "11111111",
	4266 => "11111111",
	4267 => "11111111",
	4268 => "11111111",
	4269 => "11111111",
	4270 => "11111111",
	4271 => "11111111",
	4272 => "11111111",
	4273 => "11111111",
	4274 => "11111111",
	4275 => "11111111",
	4276 => "11111111",
	4277 => "11111111",
	4278 => "11111111",
	4279 => "11111111",
	4280 => "11111111",
	4281 => "11111111",
	4282 => "11111111",
	4283 => "11111111",
	4284 => "11111111",
	4285 => "11111111",
	4286 => "11111111",
	4287 => "11111111",
	4288 => "11111111",
	4289 => "11111111",
	4290 => "11111111",
	4291 => "11111111",
	4292 => "11111111",
	4293 => "11111111",
	4294 => "11111111",
	4295 => "11111111",
	4296 => "11111111",
	4297 => "11111111",
	4298 => "11111111",
	4299 => "11111111",
	4300 => "11111111",
	4301 => "11111111",
	4302 => "11111111",
	4303 => "11111111",
	4304 => "11111111",
	4305 => "11111111",
	4306 => "11111111",
	4307 => "11111111",
	4308 => "11111111",
	4309 => "11111111",
	4310 => "11111111",
	4311 => "11111111",
	4312 => "11111111",
	4313 => "11111111",
	4314 => "11111111",
	4315 => "11111111",
	4316 => "11111111",
	4317 => "11111111",
	4318 => "11111111",
	4319 => "11111111",
	4320 => "11111111",
	4321 => "11111111",
	4322 => "11111111",
	4323 => "11111111",
	4324 => "11111111",
	4325 => "11111111",
	4326 => "11111111",
	4327 => "11111111",
	4328 => "11111111",
	4329 => "11111111",
	4330 => "11111111",
	4331 => "11111111",
	4332 => "11111111",
	4333 => "11111111",
	4334 => "11111111",
	4335 => "11111111",
	4336 => "11111111",
	4337 => "11111111",
	4338 => "11111111",
	4339 => "11111111",
	4340 => "11111111",
	4341 => "11111111",
	4342 => "11111111",
	4343 => "11111111",
	4352 => "11111111",
	4353 => "11111111",
	4354 => "11111111",
	4355 => "11111111",
	4356 => "11111111",
	4357 => "11111111",
	4358 => "11111111",
	4359 => "11111111",
	4360 => "11111111",
	4361 => "11111111",
	4362 => "11111111",
	4363 => "11111111",
	4364 => "11111111",
	4365 => "11111111",
	4366 => "11111111",
	4367 => "11111111",
	4368 => "11111111",
	4369 => "11111111",
	4370 => "11111111",
	4371 => "11111111",
	4372 => "11111111",
	4373 => "11111111",
	4374 => "11111111",
	4375 => "11111111",
	4376 => "11111111",
	4377 => "11111111",
	4378 => "11111111",
	4379 => "11111111",
	4380 => "11111111",
	4381 => "11111111",
	4382 => "11111111",
	4383 => "11111111",
	4384 => "11111111",
	4385 => "11111111",
	4386 => "11111111",
	4387 => "11111111",
	4388 => "11111111",
	4389 => "11111111",
	4390 => "11111111",
	4391 => "11111111",
	4392 => "11111111",
	4393 => "11111111",
	4394 => "11111111",
	4395 => "11111111",
	4396 => "11111111",
	4397 => "11111111",
	4398 => "11111111",
	4399 => "11111111",
	4400 => "11111111",
	4401 => "11111111",
	4402 => "11111111",
	4403 => "11111111",
	4404 => "11111111",
	4405 => "11111111",
	4406 => "11111111",
	4407 => "11111111",
	4408 => "11111111",
	4409 => "11111111",
	4410 => "11111111",
	4411 => "11111111",
	4412 => "11111111",
	4413 => "11111111",
	4414 => "11111111",
	4415 => "11111111",
	4416 => "11111111",
	4417 => "11111111",
	4418 => "11111111",
	4419 => "11111111",
	4420 => "11111111",
	4421 => "11111111",
	4422 => "11111111",
	4423 => "11111111",
	4424 => "11111111",
	4425 => "11111111",
	4426 => "11111111",
	4427 => "11111111",
	4428 => "11111111",
	4429 => "11111111",
	4430 => "11111111",
	4431 => "11111111",
	4432 => "11111111",
	4433 => "11111111",
	4434 => "11111111",
	4435 => "11111111",
	4436 => "11111111",
	4437 => "11111111",
	4438 => "11111111",
	4439 => "11111111",
	4440 => "11111111",
	4441 => "11111111",
	4442 => "11111111",
	4443 => "11111111",
	4444 => "11111111",
	4445 => "11111111",
	4446 => "11111111",
	4447 => "11111111",
	4448 => "11111111",
	4449 => "11111111",
	4450 => "11111111",
	4451 => "11111111",
	4452 => "11111111",
	4453 => "11111111",
	4454 => "11111111",
	4455 => "11111111",
	4456 => "11111111",
	4457 => "11111111",
	4458 => "11111111",
	4459 => "11111111",
	4460 => "11111111",
	4461 => "11111111",
	4462 => "11111111",
	4463 => "11111111",
	4464 => "11111111",
	4465 => "11111111",
	4466 => "11111111",
	4467 => "11111111",
	4468 => "11111111",
	4469 => "11111111",
	4470 => "11111111",
	4471 => "11111111",
	4480 => "11111111",
	4481 => "11111111",
	4482 => "11111111",
	4483 => "11111111",
	4484 => "11111111",
	4485 => "11111111",
	4486 => "11111111",
	4487 => "11111111",
	4488 => "11111111",
	4489 => "11111111",
	4490 => "11111111",
	4491 => "11111111",
	4492 => "11111111",
	4493 => "11111111",
	4494 => "11111111",
	4495 => "11111111",
	4496 => "11111111",
	4497 => "11111111",
	4498 => "11111111",
	4499 => "11111111",
	4500 => "11111111",
	4501 => "11111111",
	4502 => "11111111",
	4503 => "11111111",
	4504 => "11111111",
	4505 => "11111111",
	4506 => "11111111",
	4507 => "11111111",
	4508 => "11111111",
	4509 => "11111111",
	4510 => "11111111",
	4511 => "11111111",
	4512 => "11111111",
	4513 => "11111111",
	4514 => "11111111",
	4515 => "11111111",
	4516 => "11111111",
	4517 => "11111111",
	4518 => "11111111",
	4519 => "11111111",
	4520 => "11111111",
	4521 => "11111111",
	4522 => "11111111",
	4523 => "11111111",
	4524 => "11111111",
	4525 => "11111111",
	4526 => "11111111",
	4527 => "11111111",
	4528 => "11111111",
	4529 => "11111111",
	4530 => "11111111",
	4531 => "11111111",
	4532 => "11111111",
	4533 => "11111111",
	4534 => "11111111",
	4535 => "11111111",
	4536 => "11111111",
	4537 => "11111111",
	4538 => "11111111",
	4539 => "11111111",
	4540 => "11111111",
	4541 => "11111111",
	4542 => "11111111",
	4543 => "11111111",
	4544 => "11111111",
	4545 => "11111111",
	4546 => "11111111",
	4547 => "11111111",
	4548 => "11111111",
	4549 => "11111111",
	4550 => "11111111",
	4551 => "11111111",
	4552 => "11111111",
	4553 => "11111111",
	4554 => "11111111",
	4555 => "11111111",
	4556 => "11111111",
	4557 => "11111111",
	4558 => "11111111",
	4559 => "11111111",
	4560 => "11111111",
	4561 => "11111111",
	4562 => "11111111",
	4563 => "11111111",
	4564 => "11111111",
	4565 => "11111111",
	4566 => "11111111",
	4567 => "11111111",
	4568 => "11111111",
	4569 => "11111111",
	4570 => "11111111",
	4571 => "11111111",
	4572 => "11111111",
	4573 => "11111111",
	4574 => "11111111",
	4575 => "11111111",
	4576 => "11111111",
	4577 => "11111111",
	4578 => "11111111",
	4579 => "11111111",
	4580 => "11111111",
	4581 => "11111111",
	4582 => "11111111",
	4583 => "11111111",
	4584 => "11111111",
	4585 => "11111111",
	4586 => "11111111",
	4587 => "11111111",
	4588 => "11111111",
	4589 => "11111111",
	4590 => "11111111",
	4591 => "11111111",
	4592 => "11111111",
	4593 => "11111111",
	4594 => "11111111",
	4595 => "11111111",
	4596 => "11111111",
	4597 => "11111111",
	4598 => "11111111",
	4599 => "11111111",
	4608 => "11111111",
	4609 => "11111111",
	4610 => "11111111",
	4611 => "11111111",
	4612 => "11111111",
	4613 => "11111111",
	4614 => "11111111",
	4615 => "11111111",
	4616 => "11111111",
	4617 => "11111111",
	4618 => "11111111",
	4619 => "11111111",
	4620 => "11111111",
	4621 => "11111111",
	4622 => "11111111",
	4623 => "11111111",
	4624 => "11111111",
	4625 => "11111111",
	4626 => "11111111",
	4627 => "11111111",
	4628 => "11111111",
	4629 => "11111111",
	4630 => "11111111",
	4631 => "11111111",
	4632 => "11111111",
	4633 => "11111111",
	4634 => "11111111",
	4635 => "11111111",
	4636 => "11111111",
	4637 => "11111111",
	4638 => "11111111",
	4639 => "11111111",
	4640 => "11111111",
	4641 => "11111111",
	4642 => "11111111",
	4643 => "11111111",
	4644 => "11111111",
	4645 => "11111111",
	4646 => "11111111",
	4647 => "11111111",
	4648 => "11111111",
	4649 => "11111111",
	4650 => "11111111",
	4651 => "11111111",
	4652 => "11111111",
	4653 => "11111111",
	4654 => "11111111",
	4655 => "11111111",
	4656 => "11111111",
	4657 => "11111111",
	4658 => "11111111",
	4659 => "11111111",
	4660 => "11111111",
	4661 => "11111111",
	4662 => "11111111",
	4663 => "11111111",
	4664 => "11111111",
	4665 => "11111111",
	4666 => "11111111",
	4667 => "11111111",
	4668 => "11111111",
	4669 => "11111111",
	4670 => "11111111",
	4671 => "11111111",
	4672 => "11111111",
	4673 => "11111111",
	4674 => "11111111",
	4675 => "11111111",
	4676 => "11111111",
	4677 => "11111111",
	4678 => "11111111",
	4679 => "11111111",
	4680 => "11111111",
	4681 => "11111111",
	4682 => "11111111",
	4683 => "11111111",
	4684 => "11111111",
	4685 => "11111111",
	4686 => "11111111",
	4687 => "11111111",
	4688 => "11111111",
	4689 => "11111111",
	4690 => "11111111",
	4691 => "11111111",
	4692 => "11111111",
	4693 => "11111111",
	4694 => "11111111",
	4695 => "11111111",
	4696 => "11111111",
	4697 => "11111111",
	4698 => "11111111",
	4699 => "11111111",
	4700 => "11111111",
	4701 => "11111111",
	4702 => "11111111",
	4703 => "11111111",
	4704 => "11111111",
	4705 => "11111111",
	4706 => "11111111",
	4707 => "11111111",
	4708 => "11111111",
	4709 => "11111111",
	4710 => "11111111",
	4711 => "11111111",
	4712 => "11111111",
	4713 => "11111111",
	4714 => "11111111",
	4715 => "11111111",
	4716 => "11111111",
	4717 => "11111111",
	4718 => "11111111",
	4719 => "11111111",
	4720 => "11111111",
	4721 => "11111111",
	4722 => "11111111",
	4723 => "11111111",
	4724 => "11111111",
	4725 => "11111111",
	4726 => "11111111",
	4727 => "11111111",
	4736 => "11111111",
	4737 => "11111111",
	4738 => "11111111",
	4739 => "11111111",
	4740 => "11111111",
	4741 => "11111111",
	4742 => "11111111",
	4743 => "11111111",
	4744 => "11111111",
	4745 => "11111111",
	4746 => "11111111",
	4747 => "11111111",
	4748 => "11111111",
	4749 => "11111111",
	4750 => "11111111",
	4751 => "11111111",
	4752 => "11111111",
	4753 => "11111111",
	4754 => "11111111",
	4755 => "11111111",
	4756 => "11111111",
	4757 => "11111111",
	4758 => "11111111",
	4759 => "11111111",
	4760 => "11111111",
	4761 => "11111111",
	4762 => "11111111",
	4763 => "11111111",
	4764 => "11111111",
	4765 => "11111111",
	4766 => "11111111",
	4767 => "11111111",
	4768 => "11111111",
	4769 => "11111111",
	4770 => "11111111",
	4771 => "11111111",
	4772 => "11111111",
	4773 => "11111111",
	4774 => "11111111",
	4775 => "11111111",
	4776 => "11111111",
	4777 => "11111111",
	4778 => "11111111",
	4779 => "11111111",
	4780 => "11111111",
	4781 => "11111111",
	4782 => "11111111",
	4783 => "11111111",
	4784 => "11111111",
	4785 => "11111111",
	4786 => "11111111",
	4787 => "11111111",
	4788 => "11111111",
	4789 => "11111111",
	4790 => "11111111",
	4791 => "11111111",
	4792 => "11111111",
	4793 => "11111111",
	4794 => "11111111",
	4795 => "11111111",
	4796 => "11111111",
	4797 => "11111111",
	4798 => "11111111",
	4799 => "11111111",
	4800 => "11111111",
	4801 => "11111111",
	4802 => "11111111",
	4803 => "11111111",
	4804 => "11111111",
	4805 => "11111111",
	4806 => "11111111",
	4807 => "11111111",
	4808 => "11111111",
	4809 => "11111111",
	4810 => "11111111",
	4811 => "11111111",
	4812 => "11111111",
	4813 => "11111111",
	4814 => "11111111",
	4815 => "11111111",
	4816 => "11111111",
	4817 => "11111111",
	4818 => "11111111",
	4819 => "11111111",
	4820 => "11111111",
	4821 => "11111111",
	4822 => "11111111",
	4823 => "11111111",
	4824 => "11111111",
	4825 => "11111111",
	4826 => "11111111",
	4827 => "11111111",
	4828 => "11111111",
	4829 => "11111111",
	4830 => "11111111",
	4831 => "11111111",
	4832 => "11111111",
	4833 => "11111111",
	4834 => "11111111",
	4835 => "11111111",
	4836 => "11111111",
	4837 => "11111111",
	4838 => "11111111",
	4839 => "11111111",
	4840 => "11111111",
	4841 => "11111111",
	4842 => "11111111",
	4843 => "11111111",
	4844 => "11111111",
	4845 => "11111111",
	4846 => "11111111",
	4847 => "11111111",
	4848 => "11111111",
	4849 => "11111111",
	4850 => "11111111",
	4851 => "11111111",
	4852 => "11111111",
	4853 => "11111111",
	4854 => "11111111",
	4855 => "11111111",
	4864 => "11111111",
	4865 => "11111111",
	4866 => "11111111",
	4867 => "11111111",
	4868 => "11111111",
	4869 => "11111111",
	4870 => "11111111",
	4871 => "11111111",
	4872 => "11111111",
	4873 => "11111111",
	4874 => "11111111",
	4875 => "11111111",
	4876 => "11111111",
	4877 => "11111111",
	4878 => "11111111",
	4879 => "11111111",
	4880 => "11111111",
	4881 => "11111111",
	4882 => "11111111",
	4883 => "11111111",
	4884 => "11111111",
	4885 => "11111111",
	4886 => "11111111",
	4887 => "11111111",
	4888 => "11111111",
	4889 => "11111111",
	4890 => "11111111",
	4891 => "11111111",
	4892 => "11111111",
	4893 => "11111111",
	4894 => "11111111",
	4895 => "11111111",
	4896 => "11111111",
	4897 => "11111111",
	4898 => "11111111",
	4899 => "11111111",
	4900 => "11111111",
	4901 => "11111111",
	4902 => "11111111",
	4903 => "11111111",
	4904 => "11111111",
	4905 => "11111111",
	4906 => "11111111",
	4907 => "11111111",
	4908 => "11111111",
	4909 => "11111111",
	4910 => "11111111",
	4911 => "11111111",
	4912 => "11111111",
	4913 => "11111111",
	4914 => "11111111",
	4915 => "11111111",
	4916 => "11111111",
	4917 => "11111111",
	4918 => "11111111",
	4919 => "11111111",
	4920 => "11111111",
	4921 => "11111111",
	4922 => "11111111",
	4923 => "11111111",
	4924 => "11111111",
	4925 => "11111111",
	4926 => "11111111",
	4927 => "11111111",
	4928 => "11111111",
	4929 => "11111111",
	4930 => "11111111",
	4931 => "11111111",
	4932 => "11111111",
	4933 => "11111111",
	4934 => "11111111",
	4935 => "11111111",
	4936 => "11111111",
	4937 => "11111111",
	4938 => "11111111",
	4939 => "11111111",
	4940 => "11111111",
	4941 => "11111111",
	4942 => "11111111",
	4943 => "11111111",
	4944 => "11111111",
	4945 => "11111111",
	4946 => "11111111",
	4947 => "11111111",
	4948 => "11111111",
	4949 => "11111111",
	4950 => "11111111",
	4951 => "11111111",
	4952 => "11111111",
	4953 => "11111111",
	4954 => "11111111",
	4955 => "11111111",
	4956 => "11111111",
	4957 => "11111111",
	4958 => "11111111",
	4959 => "11111111",
	4960 => "11111111",
	4961 => "11111111",
	4962 => "11111111",
	4963 => "11111111",
	4964 => "11111111",
	4965 => "11111111",
	4966 => "11111111",
	4967 => "11111111",
	4968 => "11111111",
	4969 => "11111111",
	4970 => "11111111",
	4971 => "11111111",
	4972 => "11111111",
	4973 => "11111111",
	4974 => "11111111",
	4975 => "11111111",
	4976 => "11111111",
	4977 => "11111111",
	4978 => "11111111",
	4979 => "11111111",
	4980 => "11111111",
	4981 => "11111111",
	4982 => "11111111",
	4983 => "11111111",
	4992 => "11111111",
	4993 => "11111111",
	4994 => "11111111",
	4995 => "11111111",
	4996 => "11111111",
	4997 => "11111111",
	4998 => "11111111",
	4999 => "11111111",
	5000 => "11111111",
	5001 => "11111111",
	5002 => "11111111",
	5003 => "11111111",
	5004 => "11111111",
	5005 => "11111111",
	5006 => "11111111",
	5007 => "11111111",
	5008 => "11111111",
	5009 => "11111111",
	5010 => "11111111",
	5011 => "11111111",
	5012 => "11111111",
	5013 => "11111111",
	5014 => "11111111",
	5015 => "11111111",
	5016 => "11111111",
	5017 => "11111111",
	5018 => "11111111",
	5019 => "11111111",
	5020 => "11111111",
	5021 => "11111111",
	5022 => "11111111",
	5023 => "11111111",
	5024 => "11111111",
	5025 => "11111111",
	5026 => "11111111",
	5027 => "11111111",
	5028 => "11111111",
	5029 => "11111111",
	5030 => "11111111",
	5031 => "11111111",
	5032 => "11111111",
	5033 => "11111111",
	5034 => "11111111",
	5035 => "11111111",
	5036 => "11111111",
	5037 => "11111111",
	5038 => "11111111",
	5039 => "11111111",
	5040 => "11111111",
	5041 => "11111111",
	5042 => "11111111",
	5043 => "11111111",
	5044 => "11111111",
	5045 => "11111111",
	5046 => "11111111",
	5047 => "11111111",
	5048 => "11111111",
	5049 => "11111111",
	5050 => "11111111",
	5051 => "11111111",
	5052 => "11111111",
	5053 => "11111111",
	5054 => "11111111",
	5055 => "11111111",
	5056 => "11111111",
	5057 => "11111111",
	5058 => "11111111",
	5059 => "11111111",
	5060 => "11111111",
	5061 => "11111111",
	5062 => "11111111",
	5063 => "11111111",
	5064 => "11111111",
	5065 => "11111111",
	5066 => "11111111",
	5067 => "11111111",
	5068 => "11111111",
	5069 => "11111111",
	5070 => "11111111",
	5071 => "11111111",
	5072 => "11111111",
	5073 => "11111111",
	5074 => "11111111",
	5075 => "11111111",
	5076 => "11111111",
	5077 => "11111111",
	5078 => "11111111",
	5079 => "11111111",
	5080 => "11111111",
	5081 => "11111111",
	5082 => "11111111",
	5083 => "11111111",
	5084 => "11111111",
	5085 => "11111111",
	5086 => "11111111",
	5087 => "11111111",
	5088 => "11111111",
	5089 => "11111111",
	5090 => "11111111",
	5091 => "11111111",
	5092 => "11111111",
	5093 => "11111111",
	5094 => "11111111",
	5095 => "11111111",
	5096 => "11111111",
	5097 => "11111111",
	5098 => "11111111",
	5099 => "11111111",
	5100 => "11111111",
	5101 => "11111111",
	5102 => "11111111",
	5103 => "11111111",
	5104 => "11111111",
	5105 => "11111111",
	5106 => "11111111",
	5107 => "11111111",
	5108 => "11111111",
	5109 => "11111111",
	5110 => "11111111",
	5111 => "11111111",
	5120 => "11111111",
	5121 => "11111111",
	5122 => "11111111",
	5123 => "11111111",
	5124 => "11111111",
	5125 => "11111111",
	5126 => "11111111",
	5127 => "11111111",
	5128 => "11111111",
	5129 => "11111111",
	5130 => "11111111",
	5131 => "11111111",
	5132 => "11111111",
	5133 => "11111111",
	5134 => "11111111",
	5135 => "11111111",
	5136 => "11111111",
	5137 => "11111111",
	5138 => "11111111",
	5139 => "11111111",
	5140 => "11111111",
	5141 => "11111111",
	5142 => "11111111",
	5143 => "11111111",
	5144 => "11111111",
	5145 => "11111111",
	5146 => "11111111",
	5147 => "11111111",
	5148 => "11111111",
	5149 => "11111111",
	5150 => "11111111",
	5151 => "11111111",
	5152 => "11111111",
	5153 => "11111111",
	5154 => "11111111",
	5155 => "11111111",
	5156 => "11111111",
	5157 => "11111111",
	5158 => "11111111",
	5159 => "11111111",
	5160 => "11111111",
	5161 => "11111111",
	5162 => "11111111",
	5163 => "11111111",
	5164 => "11111111",
	5165 => "11111111",
	5166 => "11111111",
	5167 => "11111111",
	5168 => "11111111",
	5169 => "11111111",
	5170 => "11111111",
	5171 => "11111111",
	5172 => "11111111",
	5173 => "11111111",
	5174 => "11111111",
	5175 => "11111111",
	5176 => "11111111",
	5177 => "11111111",
	5178 => "11111111",
	5179 => "11111111",
	5180 => "11111111",
	5181 => "11111111",
	5182 => "11111111",
	5183 => "11111111",
	5184 => "11111111",
	5185 => "11111111",
	5186 => "11111111",
	5187 => "11111111",
	5188 => "11111111",
	5189 => "11111111",
	5190 => "11111111",
	5191 => "11111111",
	5192 => "11111111",
	5193 => "11111111",
	5194 => "11111111",
	5195 => "11111111",
	5196 => "11111111",
	5197 => "11111111",
	5198 => "11111111",
	5199 => "11111111",
	5200 => "11111111",
	5201 => "11111111",
	5202 => "11111111",
	5203 => "11111111",
	5204 => "11111111",
	5205 => "11111111",
	5206 => "11111111",
	5207 => "11111111",
	5208 => "11111111",
	5209 => "11111111",
	5210 => "11111111",
	5211 => "11111111",
	5212 => "11111111",
	5213 => "11111111",
	5214 => "11111111",
	5215 => "11111111",
	5216 => "11111111",
	5217 => "11111111",
	5218 => "11111111",
	5219 => "11111111",
	5220 => "11111111",
	5221 => "11111111",
	5222 => "11111111",
	5223 => "11111111",
	5224 => "11111111",
	5225 => "11111111",
	5226 => "11111111",
	5227 => "11111111",
	5228 => "11111111",
	5229 => "11111111",
	5230 => "11111111",
	5231 => "11111111",
	5232 => "11111111",
	5233 => "11111111",
	5234 => "11111111",
	5235 => "11111111",
	5236 => "11111111",
	5237 => "11111111",
	5238 => "11111111",
	5239 => "11111111",
	5248 => "11111111",
	5249 => "11111111",
	5250 => "11111111",
	5251 => "11111111",
	5252 => "11111111",
	5253 => "11111111",
	5254 => "11111111",
	5255 => "11111111",
	5256 => "11111111",
	5257 => "11111111",
	5258 => "11111111",
	5259 => "11111111",
	5260 => "11111111",
	5261 => "11111111",
	5262 => "11111111",
	5263 => "11111111",
	5264 => "11111111",
	5265 => "11111111",
	5266 => "11111111",
	5267 => "11111111",
	5268 => "11111111",
	5269 => "11111111",
	5270 => "11111111",
	5271 => "11111111",
	5272 => "11111111",
	5273 => "11111111",
	5274 => "11111111",
	5275 => "11111111",
	5276 => "11111111",
	5277 => "11111111",
	5278 => "11111111",
	5279 => "11111111",
	5280 => "11111111",
	5281 => "11111111",
	5282 => "11111111",
	5283 => "11111111",
	5284 => "11111111",
	5285 => "11111111",
	5286 => "11111111",
	5287 => "11111111",
	5288 => "11111111",
	5289 => "11111111",
	5290 => "11111111",
	5291 => "11111111",
	5292 => "11111111",
	5293 => "11111111",
	5294 => "11111111",
	5295 => "11111111",
	5296 => "11111111",
	5297 => "11111111",
	5298 => "11111111",
	5299 => "11111111",
	5300 => "11111111",
	5301 => "11111111",
	5302 => "11111111",
	5303 => "11111111",
	5304 => "11111111",
	5305 => "11111111",
	5306 => "11111111",
	5307 => "11111111",
	5308 => "11111111",
	5309 => "11111111",
	5310 => "11111111",
	5311 => "11111111",
	5312 => "11111111",
	5313 => "11111111",
	5314 => "11111111",
	5315 => "11111111",
	5316 => "11111111",
	5317 => "11111111",
	5318 => "11111111",
	5319 => "11111111",
	5320 => "11111111",
	5321 => "11111111",
	5322 => "11111111",
	5323 => "11111111",
	5324 => "11111111",
	5325 => "11111111",
	5326 => "11111111",
	5327 => "11111111",
	5328 => "11111111",
	5329 => "11111111",
	5330 => "11111111",
	5331 => "11111111",
	5332 => "11111111",
	5333 => "11111111",
	5334 => "11111111",
	5335 => "11111111",
	5336 => "11111111",
	5337 => "11111111",
	5338 => "11111111",
	5339 => "11111111",
	5340 => "11111111",
	5341 => "11111111",
	5342 => "11111111",
	5343 => "11111111",
	5344 => "11111111",
	5345 => "11111111",
	5346 => "11111111",
	5347 => "11111111",
	5348 => "11111111",
	5349 => "11111111",
	5350 => "11111111",
	5351 => "11111111",
	5352 => "11111111",
	5353 => "11111111",
	5354 => "11111111",
	5355 => "11111111",
	5356 => "11111111",
	5357 => "11111111",
	5358 => "11111111",
	5359 => "11111111",
	5360 => "11111111",
	5361 => "11111111",
	5362 => "11111111",
	5363 => "11111111",
	5364 => "11111111",
	5365 => "11111111",
	5366 => "11111111",
	5367 => "11111111",
	5376 => "11111111",
	5377 => "11111111",
	5378 => "11111111",
	5379 => "11111111",
	5380 => "11111111",
	5381 => "11111111",
	5382 => "11111111",
	5383 => "11111111",
	5384 => "11111111",
	5385 => "11111111",
	5386 => "11111111",
	5387 => "11111111",
	5388 => "11111111",
	5389 => "11111111",
	5390 => "11111111",
	5391 => "11111111",
	5392 => "11111111",
	5393 => "11111111",
	5394 => "11111111",
	5395 => "11111111",
	5396 => "11111111",
	5397 => "11111111",
	5398 => "11111111",
	5399 => "11111111",
	5400 => "11111111",
	5401 => "11111111",
	5402 => "11111111",
	5403 => "11111111",
	5404 => "11111111",
	5405 => "11111111",
	5406 => "11111111",
	5407 => "11111111",
	5408 => "11111111",
	5409 => "11111111",
	5410 => "11111111",
	5411 => "11111111",
	5412 => "11111111",
	5413 => "11111111",
	5414 => "11111111",
	5415 => "11111111",
	5416 => "11111111",
	5417 => "11111111",
	5418 => "11111111",
	5419 => "11111111",
	5420 => "11111111",
	5421 => "11111111",
	5422 => "11111111",
	5423 => "11111111",
	5424 => "11111111",
	5425 => "11111111",
	5426 => "11111111",
	5427 => "11111111",
	5428 => "11111111",
	5429 => "11111111",
	5430 => "11111111",
	5431 => "11111111",
	5432 => "11111111",
	5433 => "11111111",
	5434 => "11111111",
	5435 => "11111111",
	5436 => "11111111",
	5437 => "11111111",
	5438 => "11111111",
	5439 => "11111111",
	5440 => "11111111",
	5441 => "11111111",
	5442 => "11111111",
	5443 => "11111111",
	5444 => "11111111",
	5445 => "11111111",
	5446 => "11111111",
	5447 => "11111111",
	5448 => "11111111",
	5449 => "11111111",
	5450 => "11111111",
	5451 => "11111111",
	5452 => "11111111",
	5453 => "11111111",
	5454 => "11111111",
	5455 => "11111111",
	5456 => "11111111",
	5457 => "11111111",
	5458 => "11111111",
	5459 => "11111111",
	5460 => "11111111",
	5461 => "11111111",
	5462 => "11111111",
	5463 => "11111111",
	5464 => "11111111",
	5465 => "11111111",
	5466 => "11111111",
	5467 => "11111111",
	5468 => "11111111",
	5469 => "11111111",
	5470 => "11111111",
	5471 => "11111111",
	5472 => "11111111",
	5473 => "11111111",
	5474 => "11111111",
	5475 => "11111111",
	5476 => "11111111",
	5477 => "11111111",
	5478 => "11111111",
	5479 => "11111111",
	5480 => "11111111",
	5481 => "11111111",
	5482 => "11111111",
	5483 => "11111111",
	5484 => "11111111",
	5485 => "11111111",
	5486 => "11111111",
	5487 => "11111111",
	5488 => "11111111",
	5489 => "11111111",
	5490 => "11111111",
	5491 => "11111111",
	5492 => "11111111",
	5493 => "11111111",
	5494 => "11111111",
	5495 => "11111111",
	5504 => "11111111",
	5505 => "11111111",
	5506 => "11111111",
	5507 => "11111111",
	5508 => "11111111",
	5509 => "11111111",
	5510 => "11111111",
	5511 => "11111111",
	5512 => "11111111",
	5513 => "11111111",
	5514 => "11111111",
	5515 => "11111111",
	5516 => "11111111",
	5517 => "11111111",
	5518 => "11111111",
	5519 => "11111111",
	5520 => "11111111",
	5521 => "11111111",
	5522 => "11111111",
	5523 => "11111111",
	5524 => "11111111",
	5525 => "11111111",
	5526 => "11111111",
	5527 => "11111111",
	5528 => "11111111",
	5529 => "11111111",
	5530 => "11111111",
	5531 => "11111111",
	5532 => "11111111",
	5533 => "11111111",
	5534 => "11111111",
	5535 => "11111111",
	5536 => "11111111",
	5537 => "11111111",
	5538 => "11111111",
	5539 => "11111111",
	5540 => "11111111",
	5541 => "11111111",
	5542 => "11111111",
	5543 => "11111111",
	5544 => "11111111",
	5545 => "11111111",
	5546 => "11111111",
	5547 => "11111111",
	5548 => "11111111",
	5549 => "11111111",
	5550 => "11111111",
	5551 => "11111111",
	5552 => "11111111",
	5553 => "11111111",
	5554 => "11111111",
	5555 => "11111111",
	5556 => "11111111",
	5557 => "11111111",
	5558 => "11111111",
	5559 => "11111111",
	5560 => "11111111",
	5561 => "11111111",
	5562 => "11111111",
	5563 => "11111111",
	5564 => "11111111",
	5565 => "11111111",
	5566 => "11111111",
	5567 => "11111111",
	5568 => "11111111",
	5569 => "11111111",
	5570 => "11111111",
	5571 => "11111111",
	5572 => "11111111",
	5573 => "11111111",
	5574 => "11111111",
	5575 => "11111111",
	5576 => "11111111",
	5577 => "11111111",
	5578 => "11111111",
	5579 => "11111111",
	5580 => "11111111",
	5581 => "11111111",
	5582 => "11111111",
	5583 => "11111111",
	5584 => "11111111",
	5585 => "11111111",
	5586 => "11111111",
	5587 => "11111111",
	5588 => "11111111",
	5589 => "11111111",
	5590 => "11111111",
	5591 => "11111111",
	5592 => "11111111",
	5593 => "11111111",
	5594 => "11111111",
	5595 => "11111111",
	5596 => "11111111",
	5597 => "11111111",
	5598 => "11111111",
	5599 => "11111111",
	5600 => "11111111",
	5601 => "11111111",
	5602 => "11111111",
	5603 => "11111111",
	5604 => "11111111",
	5605 => "11111111",
	5606 => "11111111",
	5607 => "11111111",
	5608 => "11111111",
	5609 => "11111111",
	5610 => "11111111",
	5611 => "11111111",
	5612 => "11111111",
	5613 => "11111111",
	5614 => "11111111",
	5615 => "11111111",
	5616 => "11111111",
	5617 => "11111111",
	5618 => "11111111",
	5619 => "11111111",
	5620 => "11111111",
	5621 => "11111111",
	5622 => "11111111",
	5623 => "11111111",
	5632 => "11111111",
	5633 => "11111111",
	5634 => "11111111",
	5635 => "11111111",
	5636 => "11111111",
	5637 => "11111111",
	5638 => "11111111",
	5639 => "11111111",
	5640 => "11111111",
	5641 => "11111111",
	5642 => "11111111",
	5643 => "11111111",
	5644 => "11111111",
	5645 => "11111111",
	5646 => "11111111",
	5647 => "11111111",
	5648 => "11111111",
	5649 => "11111111",
	5650 => "11111111",
	5651 => "11111111",
	5652 => "11111111",
	5653 => "11111111",
	5654 => "11111111",
	5655 => "11111111",
	5656 => "11111111",
	5657 => "11111111",
	5658 => "11111111",
	5659 => "11111111",
	5660 => "11111111",
	5661 => "11111111",
	5662 => "11111111",
	5663 => "11111111",
	5664 => "11111111",
	5665 => "11111111",
	5666 => "11111111",
	5667 => "11111111",
	5668 => "11111111",
	5669 => "11111111",
	5670 => "11111111",
	5671 => "11111111",
	5672 => "11111111",
	5673 => "11111111",
	5674 => "11111111",
	5675 => "11111111",
	5676 => "11111111",
	5677 => "11111111",
	5678 => "11111111",
	5679 => "11111111",
	5680 => "11111111",
	5681 => "11111111",
	5682 => "11111111",
	5683 => "11111111",
	5684 => "11111111",
	5685 => "11111111",
	5686 => "11111111",
	5687 => "11111111",
	5688 => "11111111",
	5689 => "11111111",
	5690 => "11111111",
	5691 => "11111111",
	5692 => "11111111",
	5693 => "11111111",
	5694 => "11111111",
	5695 => "11111111",
	5696 => "11111111",
	5697 => "11111111",
	5698 => "11111111",
	5699 => "11111111",
	5700 => "11111111",
	5701 => "11111111",
	5702 => "11111111",
	5703 => "11111111",
	5704 => "11111111",
	5705 => "11111111",
	5706 => "11111111",
	5707 => "11111111",
	5708 => "11111111",
	5709 => "11111111",
	5710 => "11111111",
	5711 => "11111111",
	5712 => "11111111",
	5713 => "11111111",
	5714 => "11111111",
	5715 => "11111111",
	5716 => "11111111",
	5717 => "11111111",
	5718 => "11111111",
	5719 => "11111111",
	5720 => "11111111",
	5721 => "11111111",
	5722 => "11111111",
	5723 => "11111111",
	5724 => "11111111",
	5725 => "11111111",
	5726 => "11111111",
	5727 => "11111111",
	5728 => "11111111",
	5729 => "11111111",
	5730 => "11111111",
	5731 => "11111111",
	5732 => "11111111",
	5733 => "11111111",
	5734 => "11111111",
	5735 => "11111111",
	5736 => "11111111",
	5737 => "11111111",
	5738 => "11111111",
	5739 => "11111111",
	5740 => "11111111",
	5741 => "11111111",
	5742 => "11111111",
	5743 => "11111111",
	5744 => "11111111",
	5745 => "11111111",
	5746 => "11111111",
	5747 => "11111111",
	5748 => "11111111",
	5749 => "11111111",
	5750 => "11111111",
	5751 => "11111111",
	5760 => "11111111",
	5761 => "11111111",
	5762 => "11111111",
	5763 => "11111111",
	5764 => "11111111",
	5765 => "11111111",
	5766 => "11111111",
	5767 => "11111111",
	5768 => "11111111",
	5769 => "11111111",
	5770 => "11111111",
	5771 => "11111111",
	5772 => "11111111",
	5773 => "11111111",
	5774 => "11111111",
	5775 => "11111111",
	5776 => "11111111",
	5777 => "11111111",
	5778 => "11111111",
	5779 => "11111111",
	5780 => "11111111",
	5781 => "11111111",
	5782 => "11111111",
	5783 => "11111111",
	5784 => "11111111",
	5785 => "11111111",
	5786 => "11111111",
	5787 => "11111111",
	5788 => "11111111",
	5789 => "11111111",
	5790 => "11111111",
	5791 => "11111111",
	5792 => "11111111",
	5793 => "11111111",
	5794 => "11111111",
	5795 => "11111111",
	5796 => "11111111",
	5797 => "11111111",
	5798 => "11111111",
	5799 => "11111111",
	5800 => "11111111",
	5801 => "11111111",
	5802 => "11111111",
	5803 => "11111111",
	5804 => "11111111",
	5805 => "11111111",
	5806 => "11111111",
	5807 => "11111111",
	5808 => "11111111",
	5809 => "11111111",
	5810 => "11111111",
	5811 => "11111111",
	5812 => "11111111",
	5813 => "11111111",
	5814 => "11111111",
	5815 => "11111111",
	5816 => "11111111",
	5817 => "11111111",
	5818 => "11111111",
	5819 => "11111111",
	5820 => "11111111",
	5821 => "11111111",
	5822 => "11111111",
	5823 => "11111111",
	5824 => "11111111",
	5825 => "11111111",
	5826 => "11111111",
	5827 => "11111111",
	5828 => "11111111",
	5829 => "11111111",
	5830 => "11111111",
	5831 => "11111111",
	5832 => "11111111",
	5833 => "11111111",
	5834 => "11111111",
	5835 => "11111111",
	5836 => "11111111",
	5837 => "11111111",
	5838 => "11111111",
	5839 => "11111111",
	5840 => "11111111",
	5841 => "11111111",
	5842 => "11111111",
	5843 => "11111111",
	5844 => "11111111",
	5845 => "11111111",
	5846 => "11111111",
	5847 => "11111111",
	5848 => "11111111",
	5849 => "11111111",
	5850 => "11111111",
	5851 => "11111111",
	5852 => "11111111",
	5853 => "11111111",
	5854 => "11111111",
	5855 => "11111111",
	5856 => "11111111",
	5857 => "11111111",
	5858 => "11111111",
	5859 => "11111111",
	5860 => "11111111",
	5861 => "11111111",
	5862 => "11111111",
	5863 => "11111111",
	5864 => "11111111",
	5865 => "11111111",
	5866 => "11111111",
	5867 => "11111111",
	5868 => "11111111",
	5869 => "11111111",
	5870 => "11111111",
	5871 => "11111111",
	5872 => "11111111",
	5873 => "11111111",
	5874 => "11111111",
	5875 => "11111111",
	5876 => "11111111",
	5877 => "11111111",
	5878 => "11111111",
	5879 => "11111111",
	5888 => "11111111",
	5889 => "11111111",
	5890 => "11111111",
	5891 => "11111111",
	5892 => "11111111",
	5893 => "11111111",
	5894 => "11111111",
	5895 => "11111111",
	5896 => "11111111",
	5897 => "11111111",
	5898 => "11111111",
	5899 => "11111111",
	5900 => "11111111",
	5901 => "11111111",
	5902 => "11111111",
	5903 => "11111111",
	5904 => "11111111",
	5905 => "11111111",
	5906 => "11111111",
	5907 => "11111111",
	5908 => "11111111",
	5909 => "11111111",
	5910 => "11111111",
	5911 => "11111111",
	5912 => "11111111",
	5913 => "11111111",
	5914 => "11111111",
	5915 => "11111111",
	5916 => "11111111",
	5917 => "11111111",
	5918 => "11111111",
	5919 => "11111111",
	5920 => "11111111",
	5921 => "11111111",
	5922 => "11111111",
	5923 => "11111111",
	5924 => "11111111",
	5925 => "11111111",
	5926 => "11111111",
	5927 => "11111111",
	5928 => "11111111",
	5929 => "11111111",
	5930 => "11111111",
	5931 => "11111111",
	5932 => "11111111",
	5933 => "11111111",
	5934 => "11111111",
	5935 => "11111111",
	5936 => "11111111",
	5937 => "11111111",
	5938 => "11111111",
	5939 => "11111111",
	5940 => "11111111",
	5941 => "11111111",
	5942 => "11111111",
	5943 => "11111111",
	5944 => "11111111",
	5945 => "11111111",
	5946 => "11111111",
	5947 => "11111111",
	5948 => "11111111",
	5949 => "11111111",
	5950 => "11111111",
	5951 => "11111111",
	5952 => "11111111",
	5953 => "11111111",
	5954 => "11111111",
	5955 => "11111111",
	5956 => "11111111",
	5957 => "11111111",
	5958 => "11111111",
	5959 => "11111111",
	5960 => "11111111",
	5961 => "11111111",
	5962 => "11111111",
	5963 => "11111111",
	5964 => "11111111",
	5965 => "11111111",
	5966 => "11111111",
	5967 => "11111111",
	5968 => "11111111",
	5969 => "11111111",
	5970 => "11111111",
	5971 => "11111111",
	5972 => "11111111",
	5973 => "11111111",
	5974 => "11111111",
	5975 => "11111111",
	5976 => "11111111",
	5977 => "11111111",
	5978 => "11111111",
	5979 => "11111111",
	5980 => "11111111",
	5981 => "11111111",
	5982 => "11111111",
	5983 => "11111111",
	5984 => "11111111",
	5985 => "11111111",
	5986 => "11111111",
	5987 => "11111111",
	5988 => "11111111",
	5989 => "11111111",
	5990 => "11111111",
	5991 => "11111111",
	5992 => "11111111",
	5993 => "11111111",
	5994 => "11111111",
	5995 => "11111111",
	5996 => "11111111",
	5997 => "11111111",
	5998 => "11111111",
	5999 => "11111111",
	6000 => "11111111",
	6001 => "11111111",
	6002 => "11111111",
	6003 => "11111111",
	6004 => "11111111",
	6005 => "11111111",
	6006 => "11111111",
	6007 => "11111111",
	6016 => "11111111",
	6017 => "11111111",
	6018 => "11111111",
	6019 => "11111111",
	6020 => "11111111",
	6021 => "11111111",
	6022 => "11111111",
	6023 => "11111111",
	6024 => "11111111",
	6025 => "11111111",
	6026 => "11111111",
	6027 => "11111111",
	6028 => "11111111",
	6029 => "11111111",
	6030 => "11111111",
	6031 => "11111111",
	6032 => "11111111",
	6033 => "11111111",
	6034 => "11111111",
	6035 => "11111111",
	6036 => "11111111",
	6037 => "11111111",
	6038 => "11111111",
	6039 => "11111111",
	6040 => "11111111",
	6041 => "11111111",
	6042 => "11111111",
	6043 => "11111111",
	6044 => "11111111",
	6045 => "11111111",
	6046 => "11111111",
	6047 => "11111111",
	6048 => "11111111",
	6049 => "11111111",
	6050 => "11111111",
	6051 => "11111111",
	6052 => "11111111",
	6053 => "11111111",
	6054 => "11111111",
	6055 => "11111111",
	6056 => "11111111",
	6057 => "11111111",
	6058 => "11111111",
	6059 => "11111111",
	6060 => "11111111",
	6061 => "11111111",
	6062 => "11111111",
	6063 => "11111111",
	6064 => "11111111",
	6065 => "11111111",
	6066 => "11111111",
	6067 => "11111111",
	6068 => "11111111",
	6069 => "11111111",
	6070 => "11111111",
	6071 => "11111111",
	6072 => "11111111",
	6073 => "11111111",
	6074 => "11111111",
	6075 => "11111111",
	6076 => "11111111",
	6077 => "11111111",
	6078 => "11111111",
	6079 => "11111111",
	6080 => "11111111",
	6081 => "11111111",
	6082 => "11111111",
	6083 => "11111111",
	6084 => "11111111",
	6085 => "11111111",
	6086 => "11111111",
	6087 => "11111111",
	6088 => "11111111",
	6089 => "11111111",
	6090 => "11111111",
	6091 => "11111111",
	6092 => "11111111",
	6093 => "11111111",
	6094 => "11111111",
	6095 => "11111111",
	6096 => "11111111",
	6097 => "11111111",
	6098 => "11111111",
	6099 => "11111111",
	6100 => "11111111",
	6101 => "11111111",
	6102 => "11111111",
	6103 => "11111111",
	6104 => "11111111",
	6105 => "11111111",
	6106 => "11111111",
	6107 => "11111111",
	6108 => "11111111",
	6109 => "11111111",
	6110 => "11111111",
	6111 => "11111111",
	6112 => "11111111",
	6113 => "11111111",
	6114 => "11111111",
	6115 => "11111111",
	6116 => "11111111",
	6117 => "11111111",
	6118 => "11111111",
	6119 => "11111111",
	6120 => "11111111",
	6121 => "11111111",
	6122 => "11111111",
	6123 => "11111111",
	6124 => "11111111",
	6125 => "11111111",
	6126 => "11111111",
	6127 => "11111111",
	6128 => "11111111",
	6129 => "11111111",
	6130 => "11111111",
	6131 => "11111111",
	6132 => "11111111",
	6133 => "11111111",
	6134 => "11111111",
	6135 => "11111111",
	6144 => "11111111",
	6145 => "11111111",
	6146 => "11111111",
	6147 => "11111111",
	6148 => "11111111",
	6149 => "11111111",
	6150 => "11111111",
	6151 => "11111111",
	6152 => "11111111",
	6153 => "11111111",
	6154 => "11111111",
	6155 => "11111111",
	6156 => "11111111",
	6157 => "11111111",
	6158 => "11111111",
	6159 => "11111111",
	6160 => "11111111",
	6161 => "11111111",
	6162 => "11111111",
	6163 => "11111111",
	6164 => "11111111",
	6165 => "11111111",
	6166 => "11111111",
	6167 => "11111111",
	6168 => "11111111",
	6169 => "11111111",
	6170 => "11111111",
	6171 => "11111111",
	6172 => "11111111",
	6173 => "11111111",
	6174 => "11111111",
	6175 => "11111111",
	6176 => "11111111",
	6177 => "11111111",
	6178 => "11111111",
	6179 => "11111111",
	6180 => "11111111",
	6181 => "11111111",
	6182 => "11111111",
	6183 => "11111111",
	6184 => "11111111",
	6185 => "11111111",
	6186 => "11111111",
	6187 => "11111111",
	6188 => "11111111",
	6189 => "11111111",
	6190 => "11111111",
	6191 => "11111111",
	6192 => "11111111",
	6193 => "11111111",
	6194 => "11111111",
	6195 => "11111111",
	6196 => "11111111",
	6197 => "11111111",
	6198 => "11111111",
	6199 => "11111111",
	6200 => "11111111",
	6201 => "11111111",
	6202 => "11111111",
	6203 => "11111111",
	6204 => "11111111",
	6205 => "11111111",
	6206 => "11111111",
	6207 => "11111111",
	6208 => "11111111",
	6209 => "11111111",
	6210 => "11111111",
	6211 => "11111111",
	6212 => "11111111",
	6213 => "11111111",
	6214 => "11111111",
	6215 => "11111111",
	6216 => "11111111",
	6217 => "11111111",
	6218 => "11111111",
	6219 => "11111111",
	6220 => "11111111",
	6221 => "11111111",
	6222 => "11111111",
	6223 => "11111111",
	6224 => "11111111",
	6225 => "11111111",
	6226 => "11111111",
	6227 => "11111111",
	6228 => "11111111",
	6229 => "11111111",
	6230 => "11111111",
	6231 => "11111111",
	6232 => "11111111",
	6233 => "11111111",
	6234 => "11111111",
	6235 => "11111111",
	6236 => "11111111",
	6237 => "11111111",
	6238 => "11111111",
	6239 => "11111111",
	6240 => "11111111",
	6241 => "11111111",
	6242 => "11111111",
	6243 => "11111111",
	6244 => "11111111",
	6245 => "11111111",
	6246 => "11111111",
	6247 => "11111111",
	6248 => "11111111",
	6249 => "11111111",
	6250 => "11111111",
	6251 => "11111111",
	6252 => "11111111",
	6253 => "11111111",
	6254 => "11111111",
	6255 => "11111111",
	6256 => "11111111",
	6257 => "11111111",
	6258 => "11111111",
	6259 => "11111111",
	6260 => "11111111",
	6261 => "11111111",
	6262 => "11111111",
	6263 => "11111111",
	6272 => "11111111",
	6273 => "11111111",
	6274 => "11111111",
	6275 => "11111111",
	6276 => "11111111",
	6277 => "11111111",
	6278 => "11111111",
	6279 => "11111111",
	6280 => "11111111",
	6281 => "11111111",
	6282 => "11111111",
	6283 => "11111111",
	6284 => "11111111",
	6285 => "11111111",
	6286 => "11111111",
	6287 => "11111111",
	6288 => "11111111",
	6289 => "11111111",
	6290 => "11111111",
	6291 => "11111111",
	6292 => "11111111",
	6293 => "11111111",
	6294 => "11111111",
	6295 => "11111111",
	6296 => "11111111",
	6297 => "11111111",
	6298 => "11111111",
	6299 => "11111111",
	6300 => "11111111",
	6301 => "11111111",
	6302 => "11111111",
	6303 => "11111111",
	6304 => "11111111",
	6305 => "11111111",
	6306 => "11111111",
	6307 => "11111111",
	6308 => "11111111",
	6309 => "11111111",
	6310 => "11111111",
	6311 => "11111111",
	6312 => "11111111",
	6313 => "11111111",
	6314 => "11111111",
	6315 => "11111111",
	6316 => "11111111",
	6317 => "11111111",
	6318 => "11111111",
	6319 => "11111111",
	6320 => "11111111",
	6321 => "11111111",
	6322 => "11111111",
	6323 => "11111111",
	6324 => "11111111",
	6325 => "11111111",
	6326 => "11111111",
	6327 => "11111111",
	6328 => "11111111",
	6329 => "11111111",
	6330 => "11111111",
	6331 => "11111111",
	6332 => "11111111",
	6333 => "11111111",
	6334 => "11111111",
	6335 => "11111111",
	6336 => "11111111",
	6337 => "11111111",
	6338 => "11111111",
	6339 => "11111111",
	6340 => "11111111",
	6341 => "11111111",
	6342 => "11111111",
	6343 => "11111111",
	6344 => "11111111",
	6345 => "11111111",
	6346 => "11111111",
	6347 => "11111111",
	6348 => "11111111",
	6349 => "11111111",
	6350 => "11111111",
	6351 => "11111111",
	6352 => "11111111",
	6353 => "11111111",
	6354 => "11111111",
	6355 => "11111111",
	6356 => "11111111",
	6357 => "11111111",
	6358 => "11111111",
	6359 => "11111111",
	6360 => "11111111",
	6361 => "11111111",
	6362 => "11111111",
	6363 => "11111111",
	6364 => "11111111",
	6365 => "11111111",
	6366 => "11111111",
	6367 => "11111111",
	6368 => "11111111",
	6369 => "11111111",
	6370 => "11111111",
	6371 => "11111111",
	6372 => "11111111",
	6373 => "11111111",
	6374 => "11111111",
	6375 => "11111111",
	6376 => "11111111",
	6377 => "11111111",
	6378 => "11111111",
	6379 => "11111111",
	6380 => "11111111",
	6381 => "11111111",
	6382 => "11111111",
	6383 => "11111111",
	6384 => "11111111",
	6385 => "11111111",
	6386 => "11111111",
	6387 => "11111111",
	6388 => "11111111",
	6389 => "11111111",
	6390 => "11111111",
	6391 => "11111111",
	6400 => "11111111",
	6401 => "11111111",
	6402 => "11111111",
	6403 => "11111111",
	6404 => "11111111",
	6405 => "11111111",
	6406 => "11111111",
	6407 => "11111111",
	6408 => "11111111",
	6409 => "11111111",
	6410 => "11111111",
	6411 => "11111111",
	6412 => "11111111",
	6413 => "11111111",
	6414 => "11111111",
	6415 => "11111111",
	6416 => "11111111",
	6417 => "11111111",
	6418 => "11111111",
	6419 => "11111111",
	6420 => "11111111",
	6421 => "11111111",
	6422 => "11111111",
	6423 => "11111111",
	6424 => "11111111",
	6425 => "11111111",
	6426 => "11111111",
	6427 => "11111111",
	6428 => "11111111",
	6429 => "11111111",
	6430 => "11111111",
	6431 => "11111111",
	6432 => "11111111",
	6433 => "11111111",
	6434 => "11111111",
	6435 => "11111111",
	6436 => "11111111",
	6437 => "11111111",
	6438 => "11111111",
	6439 => "11111111",
	6440 => "11111111",
	6441 => "11111111",
	6442 => "11111111",
	6443 => "11111111",
	6444 => "11111111",
	6445 => "11111111",
	6446 => "11111111",
	6447 => "11111111",
	6448 => "11111111",
	6449 => "11111111",
	6450 => "11111111",
	6451 => "11111111",
	6452 => "11111111",
	6453 => "11111111",
	6454 => "11111111",
	6455 => "11111111",
	6456 => "11111111",
	6457 => "11111111",
	6458 => "11111111",
	6459 => "11111111",
	6460 => "11111111",
	6461 => "11111111",
	6462 => "11111111",
	6463 => "11111111",
	6464 => "11111111",
	6465 => "11111111",
	6466 => "11111111",
	6467 => "11111111",
	6468 => "11111111",
	6469 => "11111111",
	6470 => "11111111",
	6471 => "11111111",
	6472 => "11111111",
	6473 => "11111111",
	6474 => "11111111",
	6475 => "11111111",
	6476 => "11111111",
	6477 => "11111111",
	6478 => "11111111",
	6479 => "11111111",
	6480 => "11111111",
	6481 => "11111111",
	6482 => "11111111",
	6483 => "11111111",
	6484 => "11111111",
	6485 => "11111111",
	6486 => "11111111",
	6487 => "11111111",
	6488 => "11111111",
	6489 => "11111111",
	6490 => "11111111",
	6491 => "11111111",
	6492 => "11111111",
	6493 => "11111111",
	6494 => "11111111",
	6495 => "11111111",
	6496 => "11111111",
	6497 => "11111111",
	6498 => "11111111",
	6499 => "11111111",
	6500 => "11111111",
	6501 => "11111111",
	6502 => "11111111",
	6503 => "11111111",
	6504 => "11111111",
	6505 => "11111111",
	6506 => "11111111",
	6507 => "11111111",
	6508 => "11111111",
	6509 => "11111111",
	6510 => "11111111",
	6511 => "11111111",
	6512 => "11111111",
	6513 => "11111111",
	6514 => "11111111",
	6515 => "11111111",
	6516 => "11111111",
	6517 => "11111111",
	6518 => "11111111",
	6519 => "11111111",
	6528 => "11111111",
	6529 => "11111111",
	6530 => "11111111",
	6531 => "11111111",
	6532 => "11111111",
	6533 => "11111111",
	6534 => "11111111",
	6535 => "11111111",
	6536 => "11111111",
	6537 => "11111111",
	6538 => "11111111",
	6539 => "11111111",
	6540 => "11111111",
	6541 => "11111111",
	6542 => "11111111",
	6543 => "11111111",
	6544 => "11111111",
	6545 => "11111111",
	6546 => "11111111",
	6547 => "11111111",
	6548 => "11111111",
	6549 => "11111111",
	6550 => "11111111",
	6551 => "11111111",
	6552 => "11111111",
	6553 => "11111111",
	6554 => "11111111",
	6555 => "11111111",
	6556 => "11111111",
	6557 => "11111111",
	6558 => "11111111",
	6559 => "11111111",
	6560 => "11111111",
	6561 => "11111111",
	6562 => "11111111",
	6563 => "11111111",
	6564 => "11111111",
	6565 => "11111111",
	6566 => "11111111",
	6567 => "11111111",
	6568 => "11111111",
	6569 => "11111111",
	6570 => "11111111",
	6571 => "11111111",
	6572 => "11111111",
	6573 => "11111111",
	6574 => "11111111",
	6575 => "11111111",
	6576 => "11111111",
	6577 => "11111111",
	6578 => "11111111",
	6579 => "11111111",
	6580 => "11111111",
	6581 => "11111111",
	6582 => "11111111",
	6583 => "11111111",
	6584 => "11111111",
	6585 => "11111111",
	6586 => "11111111",
	6587 => "11111111",
	6588 => "11111111",
	6589 => "11111111",
	6590 => "11111111",
	6591 => "11111111",
	6592 => "11111111",
	6593 => "11111111",
	6594 => "11111111",
	6595 => "11111111",
	6596 => "11111111",
	6597 => "11111111",
	6598 => "11111111",
	6599 => "11111111",
	6600 => "11111111",
	6601 => "11111111",
	6602 => "11111111",
	6603 => "11111111",
	6604 => "11111111",
	6605 => "11111111",
	6606 => "11111111",
	6607 => "11111111",
	6608 => "11111111",
	6609 => "11111111",
	6610 => "11111111",
	6611 => "11111111",
	6612 => "11111111",
	6613 => "11111111",
	6614 => "11111111",
	6615 => "11111111",
	6616 => "11111111",
	6617 => "11111111",
	6618 => "11111111",
	6619 => "11111111",
	6620 => "11111111",
	6621 => "11111111",
	6622 => "11111111",
	6623 => "11111111",
	6624 => "11111111",
	6625 => "11111111",
	6626 => "11111111",
	6627 => "11111111",
	6628 => "11111111",
	6629 => "11111111",
	6630 => "11111111",
	6631 => "11111111",
	6632 => "11111111",
	6633 => "11111111",
	6634 => "11111111",
	6635 => "11111111",
	6636 => "11111111",
	6637 => "11111111",
	6638 => "11111111",
	6639 => "11111111",
	6640 => "11111111",
	6641 => "11111111",
	6642 => "11111111",
	6643 => "11111111",
	6644 => "11111111",
	6645 => "11111111",
	6646 => "11111111",
	6647 => "11111111",
	6656 => "11111111",
	6657 => "11111111",
	6658 => "11111111",
	6659 => "11111111",
	6660 => "11111111",
	6661 => "11111111",
	6662 => "11111111",
	6663 => "11111111",
	6664 => "11111111",
	6665 => "11111111",
	6666 => "11111111",
	6667 => "11111111",
	6668 => "11111111",
	6669 => "11111111",
	6670 => "11111111",
	6671 => "11111111",
	6672 => "11111111",
	6673 => "11111111",
	6674 => "11111111",
	6675 => "11111111",
	6676 => "11111111",
	6677 => "11111111",
	6678 => "11111111",
	6679 => "11111111",
	6680 => "11111111",
	6681 => "11111111",
	6682 => "11111111",
	6683 => "11111111",
	6684 => "11111111",
	6685 => "11111111",
	6686 => "11111111",
	6687 => "11111111",
	6688 => "11111111",
	6689 => "11111111",
	6690 => "11111111",
	6691 => "11111111",
	6692 => "11111111",
	6693 => "11111111",
	6694 => "11111111",
	6695 => "11111111",
	6696 => "11111111",
	6697 => "11111111",
	6698 => "11111111",
	6699 => "11111111",
	6700 => "11111111",
	6701 => "11111111",
	6702 => "11111111",
	6703 => "11111111",
	6704 => "11111111",
	6705 => "11111111",
	6706 => "11111111",
	6707 => "11111111",
	6708 => "11111111",
	6709 => "11111111",
	6710 => "11111111",
	6711 => "11111111",
	6712 => "11111111",
	6713 => "11111111",
	6714 => "11111111",
	6715 => "11111111",
	6716 => "11111111",
	6717 => "11111111",
	6718 => "11111111",
	6719 => "11111111",
	6720 => "11111111",
	6721 => "11111111",
	6722 => "11111111",
	6723 => "11111111",
	6724 => "11111111",
	6725 => "11111111",
	6726 => "11111111",
	6727 => "11111111",
	6728 => "11111111",
	6729 => "11111111",
	6730 => "11111111",
	6731 => "11111111",
	6732 => "11111111",
	6733 => "11111111",
	6734 => "11111111",
	6735 => "11111111",
	6736 => "11111111",
	6737 => "11111111",
	6738 => "11111111",
	6739 => "11111111",
	6740 => "11111111",
	6741 => "11111111",
	6742 => "11111111",
	6743 => "11111111",
	6744 => "11111111",
	6745 => "11111111",
	6746 => "11111111",
	6747 => "11111111",
	6748 => "11111111",
	6749 => "11111111",
	6750 => "11111111",
	6751 => "11111111",
	6752 => "11111111",
	6753 => "11111111",
	6754 => "11111111",
	6755 => "11111111",
	6756 => "11111111",
	6757 => "11111111",
	6758 => "11111111",
	6759 => "11111111",
	6760 => "11111111",
	6761 => "11111111",
	6762 => "11111111",
	6763 => "11111111",
	6764 => "11111111",
	6765 => "11111111",
	6766 => "11111111",
	6767 => "11111111",
	6768 => "11111111",
	6769 => "11111111",
	6770 => "11111111",
	6771 => "11111111",
	6772 => "11111111",
	6773 => "11111111",
	6774 => "11111111",
	6775 => "11111111",
	6784 => "11111111",
	6785 => "11111111",
	6786 => "11111111",
	6787 => "11111111",
	6788 => "11111111",
	6789 => "11111111",
	6790 => "11111111",
	6791 => "11111111",
	6792 => "11111111",
	6793 => "11111111",
	6794 => "11111111",
	6795 => "11111111",
	6796 => "11111111",
	6797 => "11111111",
	6798 => "11111111",
	6799 => "11111111",
	6800 => "11111111",
	6801 => "11111111",
	6802 => "11111111",
	6803 => "11111111",
	6804 => "11111111",
	6805 => "11111111",
	6806 => "11111111",
	6807 => "11111111",
	6808 => "11111111",
	6809 => "11111111",
	6810 => "11111111",
	6811 => "11111111",
	6812 => "11111111",
	6813 => "11111111",
	6814 => "11111111",
	6815 => "11111111",
	6816 => "11111111",
	6817 => "11111111",
	6818 => "11111111",
	6819 => "11111111",
	6820 => "11111111",
	6821 => "11111111",
	6822 => "11111111",
	6823 => "11111111",
	6824 => "11111111",
	6825 => "11111111",
	6826 => "11111111",
	6827 => "11111111",
	6828 => "11111111",
	6829 => "11111111",
	6830 => "11111111",
	6831 => "11111111",
	6832 => "11111111",
	6833 => "11111111",
	6834 => "11111111",
	6835 => "11111111",
	6836 => "11111111",
	6837 => "11111111",
	6838 => "11111111",
	6839 => "11111111",
	6840 => "11111111",
	6841 => "11111111",
	6842 => "11111111",
	6843 => "11111111",
	6844 => "11111111",
	6845 => "11111111",
	6846 => "11111111",
	6847 => "11111111",
	6848 => "11111111",
	6849 => "11111111",
	6850 => "11111111",
	6851 => "11111111",
	6852 => "11111111",
	6853 => "11111111",
	6854 => "11111111",
	6855 => "11111111",
	6856 => "11111111",
	6857 => "11111111",
	6858 => "11111111",
	6859 => "11111111",
	6860 => "11111111",
	6861 => "11111111",
	6862 => "11111111",
	6863 => "11111111",
	6864 => "11111111",
	6865 => "11111111",
	6866 => "11111111",
	6867 => "11111111",
	6868 => "11111111",
	6869 => "11111111",
	6870 => "11111111",
	6871 => "11111111",
	6872 => "11111111",
	6873 => "11111111",
	6874 => "11111111",
	6875 => "11111111",
	6876 => "11111111",
	6877 => "11111111",
	6878 => "11111111",
	6879 => "11111111",
	6880 => "11111111",
	6881 => "11111111",
	6882 => "11111111",
	6883 => "11111111",
	6884 => "11111111",
	6885 => "11111111",
	6886 => "11111111",
	6887 => "11111111",
	6888 => "11111111",
	6889 => "11111111",
	6890 => "11111111",
	6891 => "11111111",
	6892 => "11111111",
	6893 => "11111111",
	6894 => "11111111",
	6895 => "11111111",
	6896 => "11111111",
	6897 => "11111111",
	6898 => "11111111",
	6899 => "11111111",
	6900 => "11111111",
	6901 => "11111111",
	6902 => "11111111",
	6903 => "11111111",
	6912 => "11111111",
	6913 => "11111111",
	6914 => "11111111",
	6915 => "11111111",
	6916 => "11111111",
	6917 => "11111111",
	6918 => "11111111",
	6919 => "11111111",
	6920 => "11111111",
	6921 => "11111111",
	6922 => "11111111",
	6923 => "11111111",
	6924 => "11111111",
	6925 => "11111111",
	6926 => "11111111",
	6927 => "11111111",
	6928 => "11111111",
	6929 => "11111111",
	6930 => "11111111",
	6931 => "11111111",
	6932 => "11111111",
	6933 => "11111111",
	6934 => "11111111",
	6935 => "11111111",
	6936 => "11111111",
	6937 => "11111111",
	6938 => "11111111",
	6939 => "11111111",
	6940 => "11111111",
	6941 => "11111111",
	6942 => "11111111",
	6943 => "11111111",
	6944 => "11111111",
	6945 => "11111111",
	6946 => "11111111",
	6947 => "11111111",
	6948 => "11111111",
	6949 => "11111111",
	6950 => "11111111",
	6951 => "11111111",
	6952 => "11111111",
	6953 => "11111111",
	6954 => "11111111",
	6955 => "11111111",
	6956 => "11111111",
	6957 => "11111111",
	6958 => "11111111",
	6959 => "11111111",
	6960 => "11111111",
	6961 => "11111111",
	6962 => "11111111",
	6963 => "11111111",
	6964 => "11111111",
	6965 => "11111111",
	6966 => "11111111",
	6967 => "11111111",
	6968 => "11111111",
	6969 => "11111111",
	6970 => "11111111",
	6971 => "11111111",
	6972 => "11111111",
	6973 => "11111111",
	6974 => "11111111",
	6975 => "11111111",
	6976 => "11111111",
	6977 => "11111111",
	6978 => "11111111",
	6979 => "11111111",
	6980 => "11111111",
	6981 => "11111111",
	6982 => "11111111",
	6983 => "11111111",
	6984 => "11111111",
	6985 => "11111111",
	6986 => "11111111",
	6987 => "11111111",
	6988 => "11111111",
	6989 => "11111111",
	6990 => "11111111",
	6991 => "11111111",
	6992 => "11111111",
	6993 => "11111111",
	6994 => "11111111",
	6995 => "11111111",
	6996 => "11111111",
	6997 => "11111111",
	6998 => "11111111",
	6999 => "11111111",
	7000 => "11111111",
	7001 => "11111111",
	7002 => "11111111",
	7003 => "11111111",
	7004 => "11111111",
	7005 => "11111111",
	7006 => "11111111",
	7007 => "11111111",
	7008 => "11111111",
	7009 => "11111111",
	7010 => "11111111",
	7011 => "11111111",
	7012 => "11111111",
	7013 => "11111111",
	7014 => "11111111",
	7015 => "11111111",
	7016 => "11111111",
	7017 => "11111111",
	7018 => "11111111",
	7019 => "11111111",
	7020 => "11111111",
	7021 => "11111111",
	7022 => "11111111",
	7023 => "11111111",
	7024 => "11111111",
	7025 => "11111111",
	7026 => "11111111",
	7027 => "11111111",
	7028 => "11111111",
	7029 => "11111111",
	7030 => "11111111",
	7031 => "11111111",
	7040 => "11111111",
	7041 => "11111111",
	7042 => "11111111",
	7043 => "11111111",
	7044 => "11111111",
	7045 => "11111111",
	7046 => "11111111",
	7047 => "11111111",
	7048 => "11111111",
	7049 => "11111111",
	7050 => "11111111",
	7051 => "11111111",
	7052 => "11111111",
	7053 => "11111111",
	7054 => "11111111",
	7055 => "11111111",
	7056 => "11111111",
	7057 => "11111111",
	7058 => "11111111",
	7059 => "11111111",
	7060 => "11111111",
	7061 => "11111111",
	7062 => "11111111",
	7063 => "11111111",
	7064 => "11111111",
	7065 => "11111111",
	7066 => "11111111",
	7067 => "11111111",
	7068 => "11111111",
	7069 => "11111111",
	7070 => "11111111",
	7071 => "11111111",
	7072 => "11111111",
	7073 => "11111111",
	7074 => "11111111",
	7075 => "11111111",
	7076 => "11111111",
	7077 => "11111111",
	7078 => "11111111",
	7079 => "11111111",
	7080 => "11111111",
	7081 => "11111111",
	7082 => "11111111",
	7083 => "11111111",
	7084 => "11111111",
	7085 => "11111111",
	7086 => "11111111",
	7087 => "11111111",
	7088 => "11111111",
	7089 => "11111111",
	7090 => "11111111",
	7091 => "11111111",
	7092 => "11111111",
	7093 => "11111111",
	7094 => "11111111",
	7095 => "11111111",
	7096 => "11111111",
	7097 => "11111111",
	7098 => "11111111",
	7099 => "11111111",
	7100 => "11111111",
	7101 => "11111111",
	7102 => "11111111",
	7103 => "11111111",
	7104 => "11111111",
	7105 => "11111111",
	7106 => "11111111",
	7107 => "11111111",
	7108 => "11111111",
	7109 => "11111111",
	7110 => "11111111",
	7111 => "11111111",
	7112 => "11111111",
	7113 => "11111111",
	7114 => "11111111",
	7115 => "11111111",
	7116 => "11111111",
	7117 => "11111111",
	7118 => "11111111",
	7119 => "11111111",
	7120 => "11111111",
	7121 => "11111111",
	7122 => "11111111",
	7123 => "11111111",
	7124 => "11111111",
	7125 => "11111111",
	7126 => "11111111",
	7127 => "11111111",
	7128 => "11111111",
	7129 => "11111111",
	7130 => "11111111",
	7131 => "11111111",
	7132 => "11111111",
	7133 => "11111111",
	7134 => "11111111",
	7135 => "11111111",
	7136 => "11111111",
	7137 => "11111111",
	7138 => "11111111",
	7139 => "11111111",
	7140 => "11111111",
	7141 => "11111111",
	7142 => "11111111",
	7143 => "11111111",
	7144 => "11111111",
	7145 => "11111111",
	7146 => "11111111",
	7147 => "11111111",
	7148 => "11111111",
	7149 => "11111111",
	7150 => "11111111",
	7151 => "11111111",
	7152 => "11111111",
	7153 => "11111111",
	7154 => "11111111",
	7155 => "11111111",
	7156 => "11111111",
	7157 => "11111111",
	7158 => "11111111",
	7159 => "11111111",
	7168 => "11111111",
	7169 => "11111111",
	7170 => "11111111",
	7171 => "11111111",
	7172 => "11111111",
	7173 => "11111111",
	7174 => "11111111",
	7175 => "11111111",
	7176 => "11111111",
	7177 => "11111111",
	7178 => "11111111",
	7179 => "11111111",
	7180 => "11111111",
	7181 => "11111111",
	7182 => "11111111",
	7183 => "11111111",
	7184 => "11111111",
	7185 => "11111111",
	7186 => "11111111",
	7187 => "11111111",
	7188 => "11111111",
	7189 => "11111111",
	7190 => "11111111",
	7191 => "11111111",
	7192 => "11111111",
	7193 => "11111111",
	7194 => "11111111",
	7195 => "11111111",
	7196 => "11111111",
	7197 => "11111111",
	7198 => "11111111",
	7199 => "11111111",
	7200 => "11111111",
	7201 => "11111111",
	7202 => "11111111",
	7203 => "11111111",
	7204 => "11111111",
	7205 => "11111111",
	7206 => "11111111",
	7207 => "11111111",
	7208 => "11111111",
	7209 => "11111111",
	7210 => "11111111",
	7211 => "11111111",
	7212 => "11111111",
	7213 => "11111111",
	7214 => "11111111",
	7215 => "11111111",
	7216 => "11111111",
	7217 => "11111111",
	7218 => "11111111",
	7219 => "11111111",
	7220 => "11111111",
	7221 => "11111111",
	7222 => "11111111",
	7223 => "11111111",
	7224 => "11111111",
	7225 => "11111111",
	7226 => "11111111",
	7227 => "11111111",
	7228 => "11111111",
	7229 => "11111111",
	7230 => "11111111",
	7231 => "11111111",
	7232 => "11111111",
	7233 => "11111111",
	7234 => "11111111",
	7235 => "11111111",
	7236 => "11111111",
	7237 => "11111111",
	7238 => "11111111",
	7239 => "11111111",
	7240 => "11111111",
	7241 => "11111111",
	7242 => "11111111",
	7243 => "11111111",
	7244 => "11111111",
	7245 => "11111111",
	7246 => "11111111",
	7247 => "11111111",
	7248 => "11111111",
	7249 => "11111111",
	7250 => "11111111",
	7251 => "11111111",
	7252 => "11111111",
	7253 => "11111111",
	7254 => "11111111",
	7255 => "11111111",
	7256 => "11111111",
	7257 => "11111111",
	7258 => "11111111",
	7259 => "11111111",
	7260 => "11111111",
	7261 => "11111111",
	7262 => "11111111",
	7263 => "11111111",
	7264 => "11111111",
	7265 => "11111111",
	7266 => "11111111",
	7267 => "11111111",
	7268 => "11111111",
	7269 => "11111111",
	7270 => "11111111",
	7271 => "11111111",
	7272 => "11111111",
	7273 => "11111111",
	7274 => "11111111",
	7275 => "11111111",
	7276 => "11111111",
	7277 => "11111111",
	7278 => "11111111",
	7279 => "11111111",
	7280 => "11111111",
	7281 => "11111111",
	7282 => "11111111",
	7283 => "11111111",
	7284 => "11111111",
	7285 => "11111111",
	7286 => "11111111",
	7287 => "11111111",
	7296 => "11111111",
	7297 => "11111111",
	7298 => "11111111",
	7299 => "11111111",
	7300 => "11111111",
	7301 => "11111111",
	7302 => "11111111",
	7303 => "11111111",
	7304 => "11111111",
	7305 => "11111111",
	7306 => "11111111",
	7307 => "11111111",
	7308 => "11111111",
	7309 => "11111111",
	7310 => "11111111",
	7311 => "11111111",
	7312 => "11111111",
	7313 => "11111111",
	7314 => "11111111",
	7315 => "11111111",
	7316 => "11111111",
	7317 => "11111111",
	7318 => "11111111",
	7319 => "11111111",
	7320 => "11111111",
	7321 => "11111111",
	7322 => "11111111",
	7323 => "11111111",
	7324 => "11111111",
	7325 => "11111111",
	7326 => "11111111",
	7327 => "11111111",
	7328 => "11111111",
	7329 => "11111111",
	7330 => "11111111",
	7331 => "11111111",
	7332 => "11111111",
	7333 => "11111111",
	7334 => "11111111",
	7335 => "11111111",
	7336 => "11111111",
	7337 => "11111111",
	7338 => "11111111",
	7339 => "11111111",
	7340 => "11111111",
	7341 => "11111111",
	7342 => "11111111",
	7343 => "11111111",
	7344 => "11111111",
	7345 => "11111111",
	7346 => "11111111",
	7347 => "11111111",
	7348 => "11111111",
	7349 => "11111111",
	7350 => "11111111",
	7351 => "11111111",
	7352 => "11111111",
	7353 => "11111111",
	7354 => "11111111",
	7355 => "11111111",
	7356 => "11111111",
	7357 => "11111111",
	7358 => "11111111",
	7359 => "11111111",
	7360 => "11111111",
	7361 => "11111111",
	7362 => "11111111",
	7363 => "11111111",
	7364 => "11111111",
	7365 => "11111111",
	7366 => "11111111",
	7367 => "11111111",
	7368 => "11111111",
	7369 => "11111111",
	7370 => "11111111",
	7371 => "11111111",
	7372 => "11111111",
	7373 => "11111111",
	7374 => "11111111",
	7375 => "11111111",
	7376 => "11111111",
	7377 => "11111111",
	7378 => "11111111",
	7379 => "11111111",
	7380 => "11111111",
	7381 => "11111111",
	7382 => "11111111",
	7383 => "11111111",
	7384 => "11111111",
	7385 => "11111111",
	7386 => "11111111",
	7387 => "11111111",
	7388 => "11111111",
	7389 => "11111111",
	7390 => "11111111",
	7391 => "11111111",
	7392 => "11111111",
	7393 => "11111111",
	7394 => "11111111",
	7395 => "11111111",
	7396 => "11111111",
	7397 => "11111111",
	7398 => "11111111",
	7399 => "11111111",
	7400 => "11111111",
	7401 => "11111111",
	7402 => "11111111",
	7403 => "11111111",
	7404 => "11111111",
	7405 => "11111111",
	7406 => "11111111",
	7407 => "11111111",
	7408 => "11111111",
	7409 => "11111111",
	7410 => "11111111",
	7411 => "11111111",
	7412 => "11111111",
	7413 => "11111111",
	7414 => "11111111",
	7415 => "11111111",
	7424 => "11111111",
	7425 => "11111111",
	7426 => "11111111",
	7427 => "11111111",
	7428 => "11111111",
	7429 => "11111111",
	7430 => "11111111",
	7431 => "11111111",
	7432 => "11111111",
	7433 => "11111111",
	7434 => "11111111",
	7435 => "11111111",
	7436 => "11111111",
	7437 => "11111111",
	7438 => "11111111",
	7439 => "11111111",
	7440 => "11111111",
	7441 => "11111111",
	7442 => "11111111",
	7443 => "11111111",
	7444 => "11111111",
	7445 => "11111111",
	7446 => "11111111",
	7447 => "11111111",
	7448 => "11111111",
	7449 => "11111111",
	7450 => "11111111",
	7451 => "11111111",
	7452 => "11111111",
	7453 => "11111111",
	7454 => "11111111",
	7455 => "11111111",
	7456 => "11111111",
	7457 => "11111111",
	7458 => "11111111",
	7459 => "11111111",
	7460 => "11111111",
	7461 => "11111111",
	7462 => "11111111",
	7463 => "11111111",
	7464 => "11111111",
	7465 => "11111111",
	7466 => "11111111",
	7467 => "11111111",
	7468 => "11111111",
	7469 => "11111111",
	7470 => "11111111",
	7471 => "11111111",
	7472 => "11111111",
	7473 => "11111111",
	7474 => "11111111",
	7475 => "11111111",
	7476 => "11111111",
	7477 => "11111111",
	7478 => "11111111",
	7479 => "11111111",
	7480 => "11111111",
	7481 => "11111111",
	7482 => "11111111",
	7483 => "11111111",
	7484 => "11111111",
	7485 => "11111111",
	7486 => "11111111",
	7487 => "11111111",
	7488 => "11111111",
	7489 => "11111111",
	7490 => "11111111",
	7491 => "11111111",
	7492 => "11111111",
	7493 => "11111111",
	7494 => "11111111",
	7495 => "11111111",
	7496 => "11111111",
	7497 => "11111111",
	7498 => "11111111",
	7499 => "11111111",
	7500 => "11111111",
	7501 => "11111111",
	7502 => "11111111",
	7503 => "11111111",
	7504 => "11111111",
	7505 => "11111111",
	7506 => "11111111",
	7507 => "11111111",
	7508 => "11111111",
	7509 => "11111111",
	7510 => "11111111",
	7511 => "11111111",
	7512 => "11111111",
	7513 => "11111111",
	7514 => "11111111",
	7515 => "11111111",
	7516 => "11111111",
	7517 => "11111111",
	7518 => "11111111",
	7519 => "11111111",
	7520 => "11111111",
	7521 => "11111111",
	7522 => "11111111",
	7523 => "11111111",
	7524 => "11111111",
	7525 => "11111111",
	7526 => "11111111",
	7527 => "11111111",
	7528 => "11111111",
	7529 => "11111111",
	7530 => "11111111",
	7531 => "11111111",
	7532 => "11111111",
	7533 => "11111111",
	7534 => "11111111",
	7535 => "11111111",
	7536 => "11111111",
	7537 => "11111111",
	7538 => "11111111",
	7539 => "11111111",
	7540 => "11111111",
	7541 => "11111111",
	7542 => "11111111",
	7543 => "11111111",
	7552 => "11111111",
	7553 => "11111111",
	7554 => "11111111",
	7555 => "11111111",
	7556 => "11111111",
	7557 => "11111111",
	7558 => "11111111",
	7559 => "11111111",
	7560 => "11111111",
	7561 => "11111111",
	7562 => "11111111",
	7563 => "11111111",
	7564 => "11111111",
	7565 => "11111111",
	7566 => "11111111",
	7567 => "11111111",
	7568 => "11111111",
	7569 => "11111111",
	7570 => "11111111",
	7571 => "11111111",
	7572 => "11111111",
	7573 => "11111111",
	7574 => "11111111",
	7575 => "11111111",
	7576 => "11111111",
	7577 => "11111111",
	7578 => "11111111",
	7579 => "11111111",
	7580 => "11111111",
	7581 => "11111111",
	7582 => "11111111",
	7583 => "11111111",
	7584 => "11111111",
	7585 => "11111111",
	7586 => "11111111",
	7587 => "11111111",
	7588 => "11111111",
	7589 => "11111111",
	7590 => "11111111",
	7591 => "11111111",
	7592 => "11111111",
	7593 => "11111111",
	7594 => "11111111",
	7595 => "11111111",
	7596 => "11111111",
	7597 => "11111111",
	7598 => "11111111",
	7599 => "11111111",
	7600 => "11111111",
	7601 => "11111111",
	7602 => "11111111",
	7603 => "11111111",
	7604 => "11111111",
	7605 => "11111111",
	7606 => "11111111",
	7607 => "11111111",
	7608 => "11111111",
	7609 => "11111111",
	7610 => "11111111",
	7611 => "11111111",
	7612 => "11111111",
	7613 => "11111111",
	7614 => "11111111",
	7615 => "11111111",
	7616 => "11111111",
	7617 => "11111111",
	7618 => "11111111",
	7619 => "11111111",
	7620 => "11111111",
	7621 => "11111111",
	7622 => "11111111",
	7623 => "11111111",
	7624 => "11111111",
	7625 => "11111111",
	7626 => "11111111",
	7627 => "11111111",
	7628 => "11111111",
	7629 => "11111111",
	7630 => "11111111",
	7631 => "11111111",
	7632 => "11111111",
	7633 => "11111111",
	7634 => "11111111",
	7635 => "11111111",
	7636 => "11111111",
	7637 => "11111111",
	7638 => "11111111",
	7639 => "11111111",
	7640 => "11111111",
	7641 => "11111111",
	7642 => "11111111",
	7643 => "11111111",
	7644 => "11111111",
	7645 => "11111111",
	7646 => "11111111",
	7647 => "11111111",
	7648 => "11111111",
	7649 => "11111111",
	7650 => "11111111",
	7651 => "11111111",
	7652 => "11111111",
	7653 => "11111111",
	7654 => "11111111",
	7655 => "11111111",
	7656 => "11111111",
	7657 => "11111111",
	7658 => "11111111",
	7659 => "11111111",
	7660 => "11111111",
	7661 => "11111111",
	7662 => "11111111",
	7663 => "11111111",
	7664 => "11111111",
	7665 => "11111111",
	7666 => "11111111",
	7667 => "11111111",
	7668 => "11111111",
	7669 => "11111111",
	7670 => "11111111",
	7671 => "11111111",
	7680 => "11111111",
	7681 => "11111111",
	7682 => "11111111",
	7683 => "11111111",
	7684 => "11111111",
	7685 => "11111111",
	7686 => "11111111",
	7687 => "11111111",
	7688 => "11111111",
	7689 => "11111111",
	7690 => "11111111",
	7691 => "11111111",
	7692 => "11111111",
	7693 => "11111111",
	7694 => "11111111",
	7695 => "11111111",
	7696 => "11111111",
	7697 => "11111111",
	7698 => "11111111",
	7699 => "11111111",
	7700 => "11111111",
	7701 => "11111111",
	7702 => "11111111",
	7703 => "11111111",
	7704 => "11111111",
	7705 => "11111111",
	7706 => "11111111",
	7707 => "11111111",
	7708 => "11111111",
	7709 => "11111111",
	7710 => "11111111",
	7711 => "11111111",
	7712 => "11111111",
	7713 => "11111111",
	7714 => "11111111",
	7715 => "11111111",
	7716 => "11111111",
	7717 => "11111111",
	7718 => "11111111",
	7719 => "11111111",
	7720 => "11111111",
	7721 => "11111111",
	7722 => "11111111",
	7723 => "11111111",
	7724 => "11111111",
	7725 => "11111111",
	7726 => "11111111",
	7727 => "11111111",
	7728 => "11111111",
	7729 => "11111111",
	7730 => "11111111",
	7731 => "11111111",
	7732 => "11111111",
	7733 => "11111111",
	7734 => "11111111",
	7735 => "11111111",
	7736 => "11111111",
	7737 => "11111111",
	7738 => "11111111",
	7739 => "11111111",
	7740 => "11111111",
	7741 => "11111111",
	7742 => "11111111",
	7743 => "11111111",
	7744 => "11111111",
	7745 => "11111111",
	7746 => "11111111",
	7747 => "11111111",
	7748 => "11111111",
	7749 => "11111111",
	7750 => "11111111",
	7751 => "11111111",
	7752 => "11111111",
	7753 => "11111111",
	7754 => "11111111",
	7755 => "11111111",
	7756 => "11111111",
	7757 => "11111111",
	7758 => "11111111",
	7759 => "11111111",
	7760 => "11111111",
	7761 => "11111111",
	7762 => "11111111",
	7763 => "11111111",
	7764 => "11111111",
	7765 => "11111111",
	7766 => "11111111",
	7767 => "11111111",
	7768 => "11111111",
	7769 => "11111111",
	7770 => "11111111",
	7771 => "11111111",
	7772 => "11111111",
	7773 => "11111111",
	7774 => "11111111",
	7775 => "11111111",
	7776 => "11111111",
	7777 => "11111111",
	7778 => "11111111",
	7779 => "11111111",
	7780 => "11111111",
	7781 => "11111111",
	7782 => "11111111",
	7783 => "11111111",
	7784 => "11111111",
	7785 => "11111111",
	7786 => "11111111",
	7787 => "11111111",
	7788 => "11111111",
	7789 => "11111111",
	7790 => "11111111",
	7791 => "11111111",
	7792 => "11111111",
	7793 => "11111111",
	7794 => "11111111",
	7795 => "11111111",
	7796 => "11111111",
	7797 => "11111111",
	7798 => "11111111",
	7799 => "11111111",
	7808 => "11111111",
	7809 => "11111111",
	7810 => "11111111",
	7811 => "11111111",
	7812 => "11111111",
	7813 => "11111111",
	7814 => "11111111",
	7815 => "11111111",
	7816 => "11111111",
	7817 => "11111111",
	7818 => "11111111",
	7819 => "11111111",
	7820 => "11111111",
	7821 => "11111111",
	7822 => "11111111",
	7823 => "11111111",
	7824 => "11111111",
	7825 => "11111111",
	7826 => "11111111",
	7827 => "11111111",
	7828 => "11111111",
	7829 => "11111111",
	7830 => "11111111",
	7831 => "11111111",
	7832 => "11111111",
	7833 => "11111111",
	7834 => "11111111",
	7835 => "11111111",
	7836 => "11111111",
	7837 => "11111111",
	7838 => "11111111",
	7839 => "11111111",
	7840 => "11111111",
	7841 => "11111111",
	7842 => "11111111",
	7843 => "11111111",
	7844 => "11111111",
	7845 => "11111111",
	7846 => "11111111",
	7847 => "11111111",
	7848 => "11111111",
	7849 => "11111111",
	7850 => "11111111",
	7851 => "11111111",
	7852 => "11111111",
	7853 => "11111111",
	7854 => "11111111",
	7855 => "11111111",
	7856 => "11111111",
	7857 => "11111111",
	7858 => "11111111",
	7859 => "11111111",
	7860 => "11111111",
	7861 => "11111111",
	7862 => "11111111",
	7863 => "11111111",
	7864 => "11111111",
	7865 => "11111111",
	7866 => "11111111",
	7867 => "11111111",
	7868 => "11111111",
	7869 => "11111111",
	7870 => "11111111",
	7871 => "11111111",
	7872 => "11111111",
	7873 => "11111111",
	7874 => "11111111",
	7875 => "11111111",
	7876 => "11111111",
	7877 => "11111111",
	7878 => "11111111",
	7879 => "11111111",
	7880 => "11111111",
	7881 => "11111111",
	7882 => "11111111",
	7883 => "11111111",
	7884 => "11111111",
	7885 => "11111111",
	7886 => "11111111",
	7887 => "11111111",
	7888 => "11111111",
	7889 => "11111111",
	7890 => "11111111",
	7891 => "11111111",
	7892 => "11111111",
	7893 => "11111111",
	7894 => "11111111",
	7895 => "11111111",
	7896 => "11111111",
	7897 => "11111111",
	7898 => "11111111",
	7899 => "11111111",
	7900 => "11111111",
	7901 => "11111111",
	7902 => "11111111",
	7903 => "11111111",
	7904 => "11111111",
	7905 => "11111111",
	7906 => "11111111",
	7907 => "11111111",
	7908 => "11111111",
	7909 => "11111111",
	7910 => "11111111",
	7911 => "11111111",
	7912 => "11111111",
	7913 => "11111111",
	7914 => "11111111",
	7915 => "11111111",
	7916 => "11111111",
	7917 => "11111111",
	7918 => "11111111",
	7919 => "11111111",
	7920 => "11111111",
	7921 => "11111111",
	7922 => "11111111",
	7923 => "11111111",
	7924 => "11111111",
	7925 => "11111111",
	7926 => "11111111",
	7927 => "11111111",
	7936 => "11111111",
	7937 => "11111111",
	7938 => "11111111",
	7939 => "11111111",
	7940 => "11111111",
	7941 => "11111111",
	7942 => "11111111",
	7943 => "11111111",
	7944 => "11111111",
	7945 => "11111111",
	7946 => "11111111",
	7947 => "11111111",
	7948 => "11111111",
	7949 => "11111111",
	7950 => "11111111",
	7951 => "11111111",
	7952 => "11111111",
	7953 => "11111111",
	7954 => "11111111",
	7955 => "11111111",
	7956 => "11111111",
	7957 => "11111111",
	7958 => "11111111",
	7959 => "11111111",
	7960 => "11111111",
	7961 => "11111111",
	7962 => "11111111",
	7963 => "11111111",
	7964 => "11111111",
	7965 => "11111111",
	7966 => "11111111",
	7967 => "11111111",
	7968 => "11111111",
	7969 => "11111111",
	7970 => "11111111",
	7971 => "11111111",
	7972 => "11111111",
	7973 => "11111111",
	7974 => "11111111",
	7975 => "11111111",
	7976 => "11111111",
	7977 => "11111111",
	7978 => "11111111",
	7979 => "11111111",
	7980 => "11111111",
	7981 => "11111111",
	7982 => "11111111",
	7983 => "11111111",
	7984 => "11111111",
	7985 => "11111111",
	7986 => "11111111",
	7987 => "11111111",
	7988 => "11111111",
	7989 => "11111111",
	7990 => "11111111",
	7991 => "11111111",
	7992 => "11111111",
	7993 => "11111111",
	7994 => "11111111",
	7995 => "11111111",
	7996 => "11111111",
	7997 => "11111111",
	7998 => "11111111",
	7999 => "11111111",
	8000 => "11111111",
	8001 => "11111111",
	8002 => "11111111",
	8003 => "11111111",
	8004 => "11111111",
	8005 => "11111111",
	8006 => "11111111",
	8007 => "11111111",
	8008 => "11111111",
	8009 => "11111111",
	8010 => "11111111",
	8011 => "11111111",
	8012 => "11111111",
	8013 => "11111111",
	8014 => "11111111",
	8015 => "11111111",
	8016 => "11111111",
	8017 => "11111111",
	8018 => "11111111",
	8019 => "11111111",
	8020 => "11111111",
	8021 => "11111111",
	8022 => "11111111",
	8023 => "11111111",
	8024 => "11111111",
	8025 => "11111111",
	8026 => "11111111",
	8027 => "11111111",
	8028 => "11111111",
	8029 => "11111111",
	8030 => "11111111",
	8031 => "11111111",
	8032 => "11111111",
	8033 => "11111111",
	8034 => "11111111",
	8035 => "11111111",
	8036 => "11111111",
	8037 => "11111111",
	8038 => "11111111",
	8039 => "11111111",
	8040 => "11111111",
	8041 => "11111111",
	8042 => "11111111",
	8043 => "11111111",
	8044 => "11111111",
	8045 => "11111111",
	8046 => "11111111",
	8047 => "11111111",
	8048 => "11111111",
	8049 => "11111111",
	8050 => "11111111",
	8051 => "11111111",
	8052 => "11111111",
	8053 => "11111111",
	8054 => "11111111",
	8055 => "11111111",
	8064 => "11111111",
	8065 => "11111111",
	8066 => "11111111",
	8067 => "11111111",
	8068 => "11111111",
	8069 => "11111111",
	8070 => "11111111",
	8071 => "11111111",
	8072 => "11111111",
	8073 => "11111111",
	8074 => "11111111",
	8075 => "11111111",
	8076 => "11111111",
	8077 => "11111111",
	8078 => "11111111",
	8079 => "11111111",
	8080 => "11111111",
	8081 => "11111111",
	8082 => "11111111",
	8083 => "11111111",
	8084 => "11111111",
	8085 => "11111111",
	8086 => "11111111",
	8087 => "11111111",
	8088 => "11111111",
	8089 => "11111111",
	8090 => "11111111",
	8091 => "11111111",
	8092 => "11111111",
	8093 => "11111111",
	8094 => "11111111",
	8095 => "11111111",
	8096 => "11111111",
	8097 => "11111111",
	8098 => "11111111",
	8099 => "11111111",
	8100 => "11111111",
	8101 => "11111111",
	8102 => "11111111",
	8103 => "11111111",
	8104 => "11111111",
	8105 => "11111111",
	8106 => "11111111",
	8107 => "11111111",
	8108 => "11111111",
	8109 => "11111111",
	8110 => "11111111",
	8111 => "11111111",
	8112 => "11111111",
	8113 => "11111111",
	8114 => "11111111",
	8115 => "11111111",
	8116 => "11111111",
	8117 => "11111111",
	8118 => "11111111",
	8119 => "11111111",
	8120 => "11111111",
	8121 => "11111111",
	8122 => "11111111",
	8123 => "11111111",
	8124 => "11111111",
	8125 => "11111111",
	8126 => "11111111",
	8127 => "11111111",
	8128 => "11111111",
	8129 => "11111111",
	8130 => "11111111",
	8131 => "11111111",
	8132 => "11111111",
	8133 => "11111111",
	8134 => "11111111",
	8135 => "11111111",
	8136 => "11111111",
	8137 => "11111111",
	8138 => "11111111",
	8139 => "11111111",
	8140 => "11111111",
	8141 => "11111111",
	8142 => "11111111",
	8143 => "11111111",
	8144 => "11111111",
	8145 => "11111111",
	8146 => "11111111",
	8147 => "11111111",
	8148 => "11111111",
	8149 => "11111111",
	8150 => "11111111",
	8151 => "11111111",
	8152 => "11111111",
	8153 => "11111111",
	8154 => "11111111",
	8155 => "11111111",
	8156 => "11111111",
	8157 => "11111111",
	8158 => "11111111",
	8159 => "11111111",
	8160 => "11111111",
	8161 => "11111111",
	8162 => "11111111",
	8163 => "11111111",
	8164 => "11111111",
	8165 => "11111111",
	8166 => "11111111",
	8167 => "11111111",
	8168 => "11111111",
	8169 => "11111111",
	8170 => "11111111",
	8171 => "11111111",
	8172 => "11111111",
	8173 => "11111111",
	8174 => "11111111",
	8175 => "11111111",
	8176 => "11111111",
	8177 => "11111111",
	8178 => "11111111",
	8179 => "11111111",
	8180 => "11111111",
	8181 => "11111111",
	8182 => "11111111",
	8183 => "11111111",
	8192 => "11111111",
	8193 => "11111111",
	8194 => "11111111",
	8195 => "11111111",
	8196 => "11111111",
	8197 => "11111111",
	8198 => "11111111",
	8199 => "11111111",
	8200 => "11111111",
	8201 => "11111111",
	8202 => "11111111",
	8203 => "11111111",
	8204 => "11111111",
	8205 => "11111111",
	8206 => "11111111",
	8207 => "11111111",
	8208 => "11111111",
	8209 => "11111111",
	8210 => "11111111",
	8211 => "11111111",
	8212 => "11111111",
	8213 => "11111111",
	8214 => "11111111",
	8215 => "11111111",
	8216 => "11111111",
	8217 => "11111111",
	8218 => "11111111",
	8219 => "11111111",
	8220 => "11111111",
	8221 => "11111111",
	8222 => "11111111",
	8223 => "11111111",
	8224 => "11111111",
	8225 => "11111111",
	8226 => "11111111",
	8227 => "11111111",
	8228 => "11111111",
	8229 => "11111111",
	8230 => "11111111",
	8231 => "11111111",
	8232 => "11111111",
	8233 => "11111111",
	8234 => "11111111",
	8235 => "11111111",
	8236 => "11111111",
	8237 => "11111111",
	8238 => "11111111",
	8239 => "11111111",
	8240 => "11111111",
	8241 => "11111111",
	8242 => "11111111",
	8243 => "11111111",
	8244 => "11111111",
	8245 => "11111111",
	8246 => "11111111",
	8247 => "11111111",
	8248 => "11111111",
	8249 => "11111111",
	8250 => "11111111",
	8251 => "11111111",
	8252 => "11111111",
	8253 => "11111111",
	8254 => "11111111",
	8255 => "11111111",
	8256 => "11111111",
	8257 => "11111111",
	8258 => "11111111",
	8259 => "11111111",
	8260 => "11111111",
	8261 => "11111111",
	8262 => "11111111",
	8263 => "11111111",
	8264 => "11111111",
	8265 => "11111111",
	8266 => "11111111",
	8267 => "11111111",
	8268 => "11111111",
	8269 => "11111111",
	8270 => "11111111",
	8271 => "11111111",
	8272 => "11111111",
	8273 => "11111111",
	8274 => "11111111",
	8275 => "11111111",
	8276 => "11111111",
	8277 => "11111111",
	8278 => "11111111",
	8279 => "11111111",
	8280 => "11111111",
	8281 => "11111111",
	8282 => "11111111",
	8283 => "11111111",
	8284 => "11111111",
	8285 => "11111111",
	8286 => "11111111",
	8287 => "11111111",
	8288 => "11111111",
	8289 => "11111111",
	8290 => "11111111",
	8291 => "11111111",
	8292 => "11111111",
	8293 => "11111111",
	8294 => "11111111",
	8295 => "11111111",
	8296 => "11111111",
	8297 => "11111111",
	8298 => "11111111",
	8299 => "11111111",
	8300 => "11111111",
	8301 => "11111111",
	8302 => "11111111",
	8303 => "11111111",
	8304 => "11111111",
	8305 => "11111111",
	8306 => "11111111",
	8307 => "11111111",
	8308 => "11111111",
	8309 => "11111111",
	8310 => "11111111",
	8311 => "11111111",
	8320 => "11111111",
	8321 => "11111111",
	8322 => "11111111",
	8323 => "11111111",
	8324 => "11111111",
	8325 => "11111111",
	8326 => "11111111",
	8327 => "11111111",
	8328 => "11111111",
	8329 => "11111111",
	8330 => "11111111",
	8331 => "11111111",
	8332 => "11111111",
	8333 => "11111111",
	8334 => "11111111",
	8335 => "11111111",
	8336 => "11111111",
	8337 => "11111111",
	8338 => "11111111",
	8339 => "11111111",
	8340 => "11111111",
	8341 => "11111111",
	8342 => "11111111",
	8343 => "11111111",
	8344 => "11111111",
	8345 => "11111111",
	8346 => "11111111",
	8347 => "11111111",
	8348 => "11111111",
	8349 => "11111111",
	8350 => "11111111",
	8351 => "11111111",
	8352 => "11111111",
	8353 => "11111111",
	8354 => "11111111",
	8355 => "11111111",
	8356 => "11111111",
	8357 => "11111111",
	8358 => "11111111",
	8359 => "11111111",
	8360 => "11111111",
	8361 => "11111111",
	8362 => "11111111",
	8363 => "11111111",
	8364 => "11111111",
	8365 => "11111111",
	8366 => "11111111",
	8367 => "11111111",
	8368 => "11111111",
	8369 => "11111111",
	8370 => "11111111",
	8371 => "11111111",
	8372 => "11111111",
	8373 => "11111111",
	8374 => "11111111",
	8375 => "11111111",
	8376 => "11111111",
	8377 => "11111111",
	8378 => "11111111",
	8379 => "11111111",
	8380 => "11111111",
	8381 => "11111111",
	8382 => "11111111",
	8383 => "11111111",
	8384 => "11111111",
	8385 => "11111111",
	8386 => "11111111",
	8387 => "11111111",
	8388 => "11111111",
	8389 => "11111111",
	8390 => "11111111",
	8391 => "11111111",
	8392 => "11111111",
	8393 => "11111111",
	8394 => "11111111",
	8395 => "11111111",
	8396 => "11111111",
	8397 => "11111111",
	8398 => "11111111",
	8399 => "11111111",
	8400 => "11111111",
	8401 => "11111111",
	8402 => "11111111",
	8403 => "11111111",
	8404 => "11111111",
	8405 => "11111111",
	8406 => "11111111",
	8407 => "11111111",
	8408 => "11111111",
	8409 => "11111111",
	8410 => "11111111",
	8411 => "11111111",
	8412 => "11111111",
	8413 => "11111111",
	8414 => "11111111",
	8415 => "11111111",
	8416 => "11111111",
	8417 => "11111111",
	8418 => "11111111",
	8419 => "11111111",
	8420 => "11111111",
	8421 => "11111111",
	8422 => "11111111",
	8423 => "11111111",
	8424 => "11111111",
	8425 => "11111111",
	8426 => "11111111",
	8427 => "11111111",
	8428 => "11111111",
	8429 => "11111111",
	8430 => "11111111",
	8431 => "11111111",
	8432 => "11111111",
	8433 => "11111111",
	8434 => "11111111",
	8435 => "11111111",
	8436 => "11111111",
	8437 => "11111111",
	8438 => "11111111",
	8439 => "11111111",
	8448 => "11111111",
	8449 => "11111111",
	8450 => "11111111",
	8451 => "11111111",
	8452 => "11111111",
	8453 => "11111111",
	8454 => "11111111",
	8455 => "11111111",
	8456 => "11111111",
	8457 => "11111111",
	8458 => "11111111",
	8459 => "11111111",
	8460 => "11111111",
	8461 => "11111111",
	8462 => "11111111",
	8463 => "11111111",
	8464 => "11111111",
	8465 => "11111111",
	8466 => "11111111",
	8467 => "11111111",
	8468 => "11111111",
	8469 => "11111111",
	8470 => "11111111",
	8471 => "11111111",
	8472 => "11111111",
	8473 => "11111111",
	8474 => "11111111",
	8475 => "11111111",
	8476 => "11111111",
	8477 => "11111111",
	8478 => "11111111",
	8479 => "11111111",
	8480 => "11111111",
	8481 => "11111111",
	8482 => "11111111",
	8483 => "11111111",
	8484 => "11111111",
	8485 => "11111111",
	8486 => "11111111",
	8487 => "11111111",
	8488 => "11111111",
	8489 => "11111111",
	8490 => "11111111",
	8491 => "11111111",
	8492 => "11111111",
	8493 => "11111111",
	8494 => "11111111",
	8495 => "11111111",
	8496 => "11111111",
	8497 => "11111111",
	8498 => "11111111",
	8499 => "11111111",
	8500 => "11111111",
	8501 => "11111111",
	8502 => "11111111",
	8503 => "11111111",
	8504 => "11111111",
	8505 => "11111111",
	8506 => "11111111",
	8507 => "11111111",
	8508 => "11111111",
	8509 => "11111111",
	8510 => "11111111",
	8511 => "11111111",
	8512 => "11111111",
	8513 => "11111111",
	8514 => "11111111",
	8515 => "11111111",
	8516 => "11111111",
	8517 => "11111111",
	8518 => "11111111",
	8519 => "11111111",
	8520 => "11111111",
	8521 => "11111111",
	8522 => "11111111",
	8523 => "11111111",
	8524 => "11111111",
	8525 => "11111111",
	8526 => "11111111",
	8527 => "11111111",
	8528 => "11111111",
	8529 => "11111111",
	8530 => "11111111",
	8531 => "11111111",
	8532 => "11111111",
	8533 => "11111111",
	8534 => "11111111",
	8535 => "11111111",
	8536 => "11111111",
	8537 => "11111111",
	8538 => "11111111",
	8539 => "11111111",
	8540 => "11111111",
	8541 => "11111111",
	8542 => "11111111",
	8543 => "11111111",
	8544 => "11111111",
	8545 => "11111111",
	8546 => "11111111",
	8547 => "11111111",
	8548 => "11111111",
	8549 => "11111111",
	8550 => "11111111",
	8551 => "11111111",
	8552 => "11111111",
	8553 => "11111111",
	8554 => "11111111",
	8555 => "11111111",
	8556 => "11111111",
	8557 => "11111111",
	8558 => "11111111",
	8559 => "11111111",
	8560 => "11111111",
	8561 => "11111111",
	8562 => "11111111",
	8563 => "11111111",
	8564 => "11111111",
	8565 => "11111111",
	8566 => "11111111",
	8567 => "11111111",
	8576 => "11111111",
	8577 => "11111111",
	8578 => "11111111",
	8579 => "11111111",
	8580 => "11111111",
	8581 => "11111111",
	8582 => "11111111",
	8583 => "11111111",
	8584 => "11111111",
	8585 => "11111111",
	8586 => "11111111",
	8587 => "11111111",
	8588 => "11111111",
	8589 => "11111111",
	8590 => "11111111",
	8591 => "11111111",
	8592 => "11111111",
	8593 => "11111111",
	8594 => "11111111",
	8595 => "11111111",
	8596 => "11111111",
	8597 => "11111111",
	8598 => "11111111",
	8599 => "11111111",
	8600 => "11111111",
	8601 => "11111111",
	8602 => "11111111",
	8603 => "11111111",
	8604 => "11111111",
	8605 => "11111111",
	8606 => "11111111",
	8607 => "11111111",
	8608 => "11111111",
	8609 => "11111111",
	8610 => "11111111",
	8611 => "11111111",
	8612 => "11111111",
	8613 => "11111111",
	8614 => "11111111",
	8615 => "11111111",
	8616 => "11111111",
	8617 => "11111111",
	8618 => "11111111",
	8619 => "11111111",
	8620 => "11111111",
	8621 => "11111111",
	8622 => "11111111",
	8623 => "11111111",
	8624 => "11111111",
	8625 => "11111111",
	8626 => "11111111",
	8627 => "11111111",
	8628 => "11111111",
	8629 => "11111111",
	8630 => "11111111",
	8631 => "11111111",
	8632 => "11111111",
	8633 => "11111111",
	8634 => "11111111",
	8635 => "11111111",
	8636 => "11111111",
	8637 => "11111111",
	8638 => "11111111",
	8639 => "11111111",
	8640 => "11111111",
	8641 => "11111111",
	8642 => "11111111",
	8643 => "11111111",
	8644 => "11111111",
	8645 => "11111111",
	8646 => "11111111",
	8647 => "11111111",
	8648 => "11111111",
	8649 => "11111111",
	8650 => "11111111",
	8651 => "11111111",
	8652 => "11111111",
	8653 => "11111111",
	8654 => "11111111",
	8655 => "11111111",
	8656 => "11111111",
	8657 => "11111111",
	8658 => "11111111",
	8659 => "11111111",
	8660 => "11111111",
	8661 => "11111111",
	8662 => "11111111",
	8663 => "11111111",
	8664 => "11111111",
	8665 => "11111111",
	8666 => "11111111",
	8667 => "11111111",
	8668 => "11111111",
	8669 => "11111111",
	8670 => "11111111",
	8671 => "11111111",
	8672 => "11111111",
	8673 => "11111111",
	8674 => "11111111",
	8675 => "11111111",
	8676 => "11111111",
	8677 => "11111111",
	8678 => "11111111",
	8679 => "11111111",
	8680 => "11111111",
	8681 => "11111111",
	8682 => "11111111",
	8683 => "11111111",
	8684 => "11111111",
	8685 => "11111111",
	8686 => "11111111",
	8687 => "11111111",
	8688 => "11111111",
	8689 => "11111111",
	8690 => "11111111",
	8691 => "11111111",
	8692 => "11111111",
	8693 => "11111111",
	8694 => "11111111",
	8695 => "11111111",
	8704 => "11111111",
	8705 => "11111111",
	8706 => "11111111",
	8707 => "11111111",
	8708 => "11111111",
	8709 => "11111111",
	8710 => "11111111",
	8711 => "11111111",
	8712 => "11111111",
	8713 => "11111111",
	8714 => "11111111",
	8715 => "11111111",
	8716 => "11111111",
	8717 => "11111111",
	8718 => "11111111",
	8719 => "11111111",
	8720 => "11111111",
	8721 => "11111111",
	8722 => "11111111",
	8723 => "11111111",
	8724 => "11111111",
	8725 => "11111111",
	8726 => "11111111",
	8727 => "11111111",
	8728 => "11111111",
	8729 => "11111111",
	8730 => "11111111",
	8731 => "11111111",
	8732 => "11111111",
	8733 => "11111111",
	8734 => "11111111",
	8735 => "11111111",
	8736 => "11111111",
	8737 => "11111111",
	8738 => "11111111",
	8739 => "11111111",
	8740 => "11111111",
	8741 => "11111111",
	8742 => "11111111",
	8743 => "11111111",
	8744 => "11111111",
	8745 => "11111111",
	8746 => "11111111",
	8747 => "11111111",
	8748 => "11111111",
	8749 => "11111111",
	8750 => "11111111",
	8751 => "11111111",
	8752 => "11111111",
	8753 => "11111111",
	8754 => "11111111",
	8755 => "11111111",
	8756 => "11111111",
	8757 => "11111111",
	8758 => "11111111",
	8759 => "11111111",
	8760 => "11111111",
	8761 => "11111111",
	8762 => "11111111",
	8763 => "11111111",
	8764 => "11111111",
	8765 => "11111111",
	8766 => "11111111",
	8767 => "11111111",
	8768 => "11111111",
	8769 => "11111111",
	8770 => "11111111",
	8771 => "11111111",
	8772 => "11111111",
	8773 => "11111111",
	8774 => "11111111",
	8775 => "11111111",
	8776 => "11111111",
	8777 => "11111111",
	8778 => "11111111",
	8779 => "11111111",
	8780 => "11111111",
	8781 => "11111111",
	8782 => "11111111",
	8783 => "11111111",
	8784 => "11111111",
	8785 => "11111111",
	8786 => "11111111",
	8787 => "11111111",
	8788 => "11111111",
	8789 => "11111111",
	8790 => "11111111",
	8791 => "11111111",
	8792 => "11111111",
	8793 => "11111111",
	8794 => "11111111",
	8795 => "11111111",
	8796 => "11111111",
	8797 => "11111111",
	8798 => "11111111",
	8799 => "11111111",
	8800 => "11111111",
	8801 => "11111111",
	8802 => "11111111",
	8803 => "11111111",
	8804 => "11111111",
	8805 => "11111111",
	8806 => "11111111",
	8807 => "11111111",
	8808 => "11111111",
	8809 => "11111111",
	8810 => "11111111",
	8811 => "11111111",
	8812 => "11111111",
	8813 => "11111111",
	8814 => "11111111",
	8815 => "11111111",
	8816 => "11111111",
	8817 => "11111111",
	8818 => "11111111",
	8819 => "11111111",
	8820 => "11111111",
	8821 => "11111111",
	8822 => "11111111",
	8823 => "11111111",
	8832 => "11111111",
	8833 => "11111111",
	8834 => "11111111",
	8835 => "11111111",
	8836 => "11111111",
	8837 => "11111111",
	8838 => "11111111",
	8839 => "11111111",
	8840 => "11111111",
	8841 => "11111111",
	8842 => "11111111",
	8843 => "11111111",
	8844 => "11111111",
	8845 => "11111111",
	8846 => "11111111",
	8847 => "11111111",
	8848 => "11111111",
	8849 => "11111111",
	8850 => "11111111",
	8851 => "11111111",
	8852 => "11111111",
	8853 => "11111111",
	8854 => "11111111",
	8855 => "11111111",
	8856 => "11111111",
	8857 => "11111111",
	8858 => "11111111",
	8859 => "11111111",
	8860 => "11111111",
	8861 => "11111111",
	8862 => "11111111",
	8863 => "11111111",
	8864 => "11111111",
	8865 => "11111111",
	8866 => "11111111",
	8867 => "11111111",
	8868 => "11111111",
	8869 => "11111111",
	8870 => "11111111",
	8871 => "11111111",
	8872 => "11111111",
	8873 => "11111111",
	8874 => "11111111",
	8875 => "11111111",
	8876 => "11111111",
	8877 => "11111111",
	8878 => "11111111",
	8879 => "11111111",
	8880 => "11111111",
	8881 => "11111111",
	8882 => "11111111",
	8883 => "11111111",
	8884 => "11111111",
	8885 => "11111111",
	8886 => "11111111",
	8887 => "11111111",
	8888 => "11111111",
	8889 => "11111111",
	8890 => "11111111",
	8891 => "11111111",
	8892 => "11111111",
	8893 => "11111111",
	8894 => "11111111",
	8895 => "11111111",
	8896 => "11111111",
	8897 => "11111111",
	8898 => "11111111",
	8899 => "11111111",
	8900 => "11111111",
	8901 => "11111111",
	8902 => "11111111",
	8903 => "11111111",
	8904 => "11111111",
	8905 => "11111111",
	8906 => "11111111",
	8907 => "11111111",
	8908 => "11111111",
	8909 => "11111111",
	8910 => "11111111",
	8911 => "11111111",
	8912 => "11111111",
	8913 => "11111111",
	8914 => "11111111",
	8915 => "11111111",
	8916 => "11111111",
	8917 => "11111111",
	8918 => "11111111",
	8919 => "11111111",
	8920 => "11111111",
	8921 => "11111111",
	8922 => "11111111",
	8923 => "11111111",
	8924 => "11111111",
	8925 => "11111111",
	8926 => "11111111",
	8927 => "11111111",
	8928 => "11111111",
	8929 => "11111111",
	8930 => "11111111",
	8931 => "11111111",
	8932 => "11111111",
	8933 => "11111111",
	8934 => "11111111",
	8935 => "11111111",
	8936 => "11111111",
	8937 => "11111111",
	8938 => "11111111",
	8939 => "11111111",
	8940 => "11111111",
	8941 => "11111111",
	8942 => "11111111",
	8943 => "11111111",
	8944 => "11111111",
	8945 => "11111111",
	8946 => "11111111",
	8947 => "11111111",
	8948 => "11111111",
	8949 => "11111111",
	8950 => "11111111",
	8951 => "11111111",
	8960 => "11111111",
	8961 => "11111111",
	8962 => "11111111",
	8963 => "11111111",
	8964 => "11111111",
	8965 => "11111111",
	8966 => "11111111",
	8967 => "11111111",
	8968 => "11111111",
	8969 => "11111111",
	8970 => "11111111",
	8971 => "11111111",
	8972 => "11111111",
	8973 => "11111111",
	8974 => "11111111",
	8975 => "11111111",
	8976 => "11111111",
	8977 => "11111111",
	8978 => "11111111",
	8979 => "11111111",
	8980 => "11111111",
	8981 => "11111111",
	8982 => "11111111",
	8983 => "11111111",
	8984 => "11111111",
	8985 => "11111111",
	8986 => "11111111",
	8987 => "11111111",
	8988 => "11111111",
	8989 => "11111111",
	8990 => "11111111",
	8991 => "11111111",
	8992 => "11111111",
	8993 => "11111111",
	8994 => "11111111",
	8995 => "11111111",
	8996 => "11111111",
	8997 => "11111111",
	8998 => "11111111",
	8999 => "11111111",
	9000 => "11111111",
	9001 => "11111111",
	9002 => "11111111",
	9003 => "11111111",
	9004 => "11111111",
	9005 => "11111111",
	9006 => "11111111",
	9007 => "11111111",
	9008 => "11111111",
	9009 => "11111111",
	9010 => "11111111",
	9011 => "11111111",
	9012 => "11111111",
	9013 => "11111111",
	9014 => "11111111",
	9015 => "11111111",
	9016 => "11111111",
	9017 => "11111111",
	9018 => "11111111",
	9019 => "11111111",
	9020 => "11111111",
	9021 => "11111111",
	9022 => "11111111",
	9023 => "11111111",
	9024 => "11111111",
	9025 => "11111111",
	9026 => "11111111",
	9027 => "11111111",
	9028 => "11111111",
	9029 => "11111111",
	9030 => "11111111",
	9031 => "11111111",
	9032 => "11111111",
	9033 => "11111111",
	9034 => "11111111",
	9035 => "11111111",
	9036 => "11111111",
	9037 => "11111111",
	9038 => "11111111",
	9039 => "11111111",
	9040 => "11111111",
	9041 => "11111111",
	9042 => "11111111",
	9043 => "11111111",
	9044 => "11111111",
	9045 => "11111111",
	9046 => "11111111",
	9047 => "11111111",
	9048 => "11111111",
	9049 => "11111111",
	9050 => "11111111",
	9051 => "11111111",
	9052 => "11111111",
	9053 => "11111111",
	9054 => "11111111",
	9055 => "11111111",
	9056 => "11111111",
	9057 => "11111111",
	9058 => "11111111",
	9059 => "11111111",
	9060 => "11111111",
	9061 => "11111111",
	9062 => "11111111",
	9063 => "11111111",
	9064 => "11111111",
	9065 => "11111111",
	9066 => "11111111",
	9067 => "11111111",
	9068 => "11111111",
	9069 => "11111111",
	9070 => "11111111",
	9071 => "11111111",
	9072 => "11111111",
	9073 => "11111111",
	9074 => "11111111",
	9075 => "11111111",
	9076 => "11111111",
	9077 => "11111111",
	9078 => "11111111",
	9079 => "11111111",
	9088 => "11111111",
	9089 => "11111111",
	9090 => "11111111",
	9091 => "11111111",
	9092 => "11111111",
	9093 => "11111111",
	9094 => "11111111",
	9095 => "11111111",
	9096 => "11111111",
	9097 => "11111111",
	9098 => "11111111",
	9099 => "11111111",
	9100 => "11111111",
	9101 => "11111111",
	9102 => "11111111",
	9103 => "11111111",
	9104 => "11111111",
	9105 => "11111111",
	9106 => "11111111",
	9107 => "11111111",
	9108 => "11111111",
	9109 => "11111111",
	9110 => "11111111",
	9111 => "11111111",
	9112 => "11111111",
	9113 => "11111111",
	9114 => "11111111",
	9115 => "11111111",
	9116 => "11111111",
	9117 => "11111111",
	9118 => "11111111",
	9119 => "11111111",
	9120 => "11111111",
	9121 => "11111111",
	9122 => "11111111",
	9123 => "11111111",
	9124 => "11111111",
	9125 => "11111111",
	9126 => "11111111",
	9127 => "11111111",
	9128 => "11111111",
	9129 => "11111111",
	9130 => "11111111",
	9131 => "11111111",
	9132 => "11111111",
	9133 => "11111111",
	9134 => "11111111",
	9135 => "11111111",
	9136 => "11111111",
	9137 => "11111111",
	9138 => "11111111",
	9139 => "11111111",
	9140 => "11111111",
	9141 => "11111111",
	9142 => "11111111",
	9143 => "11111111",
	9144 => "11111111",
	9145 => "11111111",
	9146 => "11111111",
	9147 => "11111111",
	9148 => "11111111",
	9149 => "11111111",
	9150 => "11111111",
	9151 => "11111111",
	9152 => "11111111",
	9153 => "11111111",
	9154 => "11111111",
	9155 => "11111111",
	9156 => "11111111",
	9157 => "11111111",
	9158 => "11111111",
	9159 => "11111111",
	9160 => "11111111",
	9161 => "11111111",
	9162 => "11111111",
	9163 => "11111111",
	9164 => "11111111",
	9165 => "11111111",
	9166 => "11111111",
	9167 => "11111111",
	9168 => "11111111",
	9169 => "11111111",
	9170 => "11111111",
	9171 => "11111111",
	9172 => "11111111",
	9173 => "11111111",
	9174 => "11111111",
	9175 => "11111111",
	9176 => "11111111",
	9177 => "11111111",
	9178 => "11111111",
	9179 => "11111111",
	9180 => "11111111",
	9181 => "11111111",
	9182 => "11111111",
	9183 => "11111111",
	9184 => "11111111",
	9185 => "11111111",
	9186 => "11111111",
	9187 => "11111111",
	9188 => "11111111",
	9189 => "11111111",
	9190 => "11111111",
	9191 => "11111111",
	9192 => "11111111",
	9193 => "11111111",
	9194 => "11111111",
	9195 => "11111111",
	9196 => "11111111",
	9197 => "11111111",
	9198 => "11111111",
	9199 => "11111111",
	9200 => "11111111",
	9201 => "11111111",
	9202 => "11111111",
	9203 => "11111111",
	9204 => "11111111",
	9205 => "11111111",
	9206 => "11111111",
	9207 => "11111111",
	9216 => "11111111",
	9217 => "11111111",
	9218 => "11111111",
	9219 => "11111111",
	9220 => "11111111",
	9221 => "11111111",
	9222 => "11111111",
	9223 => "11111111",
	9224 => "11111111",
	9225 => "11111111",
	9226 => "11111111",
	9227 => "11111111",
	9228 => "11111111",
	9229 => "11111111",
	9230 => "11111111",
	9231 => "11111111",
	9232 => "11111111",
	9233 => "11111111",
	9234 => "11111111",
	9235 => "11111111",
	9236 => "11111111",
	9237 => "11111111",
	9238 => "11111111",
	9239 => "11111111",
	9240 => "11111111",
	9241 => "11111111",
	9242 => "11111111",
	9243 => "11111111",
	9244 => "11111111",
	9245 => "11111111",
	9246 => "11111111",
	9247 => "11111111",
	9248 => "11111111",
	9249 => "11111111",
	9250 => "11111111",
	9251 => "11111111",
	9252 => "11111111",
	9253 => "11111111",
	9254 => "11111111",
	9255 => "11111111",
	9256 => "11111111",
	9257 => "11111111",
	9258 => "11111111",
	9259 => "11111111",
	9260 => "11111111",
	9261 => "11111111",
	9262 => "11111111",
	9263 => "11111111",
	9264 => "11111111",
	9265 => "11111111",
	9266 => "11111111",
	9267 => "11111111",
	9268 => "11111111",
	9269 => "11111111",
	9270 => "11111111",
	9271 => "11111111",
	9272 => "11111111",
	9273 => "11111111",
	9274 => "11111111",
	9275 => "11111111",
	9276 => "11111111",
	9277 => "11111111",
	9278 => "11111111",
	9279 => "11111111",
	9280 => "11111111",
	9281 => "11111111",
	9282 => "11111111",
	9283 => "11111111",
	9284 => "11111111",
	9285 => "11111111",
	9286 => "11111111",
	9287 => "11111111",
	9288 => "11111111",
	9289 => "11111111",
	9290 => "11111111",
	9291 => "11111111",
	9292 => "11111111",
	9293 => "11111111",
	9294 => "11111111",
	9295 => "11111111",
	9296 => "11111111",
	9297 => "11111111",
	9298 => "11111111",
	9299 => "11111111",
	9300 => "11111111",
	9301 => "11111111",
	9302 => "11111111",
	9303 => "11111111",
	9304 => "11111111",
	9305 => "11111111",
	9306 => "11111111",
	9307 => "11111111",
	9308 => "11111111",
	9309 => "11111111",
	9310 => "11111111",
	9311 => "11111111",
	9312 => "11111111",
	9313 => "11111111",
	9314 => "11111111",
	9315 => "11111111",
	9316 => "11111111",
	9317 => "11111111",
	9318 => "11111111",
	9319 => "11111111",
	9320 => "11111111",
	9321 => "11111111",
	9322 => "11111111",
	9323 => "11111111",
	9324 => "11111111",
	9325 => "11111111",
	9326 => "11111111",
	9327 => "11111111",
	9328 => "11111111",
	9329 => "11111111",
	9330 => "11111111",
	9331 => "11111111",
	9332 => "11111111",
	9333 => "11111111",
	9334 => "11111111",
	9335 => "11111111",
	9344 => "11111111",
	9345 => "11111111",
	9346 => "11111111",
	9347 => "11111111",
	9348 => "11111111",
	9349 => "11111111",
	9350 => "11111111",
	9351 => "11111111",
	9352 => "11111111",
	9353 => "11111111",
	9354 => "11111111",
	9355 => "11111111",
	9356 => "11111111",
	9357 => "11111111",
	9358 => "11111111",
	9359 => "11111111",
	9360 => "11111111",
	9361 => "11111111",
	9362 => "11111111",
	9363 => "11111111",
	9364 => "11111111",
	9365 => "11111111",
	9366 => "11111111",
	9367 => "11111111",
	9368 => "11111111",
	9369 => "11111111",
	9370 => "11111111",
	9371 => "11111111",
	9372 => "11111111",
	9373 => "11111111",
	9374 => "11111111",
	9375 => "11111111",
	9376 => "11111111",
	9377 => "11111111",
	9378 => "11111111",
	9379 => "11111111",
	9380 => "11111111",
	9381 => "11111111",
	9382 => "11111111",
	9383 => "11111111",
	9384 => "11111111",
	9385 => "11111111",
	9386 => "11111111",
	9387 => "11111111",
	9388 => "11111111",
	9389 => "11111111",
	9390 => "11111111",
	9391 => "11111111",
	9392 => "11111111",
	9393 => "11111111",
	9394 => "11111111",
	9395 => "11111111",
	9396 => "11111111",
	9397 => "11111111",
	9398 => "11111111",
	9399 => "11111111",
	9400 => "11111111",
	9401 => "11111111",
	9402 => "11111111",
	9403 => "11111111",
	9404 => "11111111",
	9405 => "11111111",
	9406 => "11111111",
	9407 => "11111111",
	9408 => "11111111",
	9409 => "11111111",
	9410 => "11111111",
	9411 => "11111111",
	9412 => "11111111",
	9413 => "11111111",
	9414 => "11111111",
	9415 => "11111111",
	9416 => "11111111",
	9417 => "11111111",
	9418 => "11111111",
	9419 => "11111111",
	9420 => "11111111",
	9421 => "11111111",
	9422 => "11111111",
	9423 => "11111111",
	9424 => "11111111",
	9425 => "11111111",
	9426 => "11111111",
	9427 => "11111111",
	9428 => "11111111",
	9429 => "11111111",
	9430 => "11111111",
	9431 => "11111111",
	9432 => "11111111",
	9433 => "11111111",
	9434 => "11111111",
	9435 => "11111111",
	9436 => "11111111",
	9437 => "11111111",
	9438 => "11111111",
	9439 => "11111111",
	9440 => "11111111",
	9441 => "11111111",
	9442 => "11111111",
	9443 => "11111111",
	9444 => "11111111",
	9445 => "11111111",
	9446 => "11111111",
	9447 => "11111111",
	9448 => "11111111",
	9449 => "11111111",
	9450 => "11111111",
	9451 => "11111111",
	9452 => "11111111",
	9453 => "11111111",
	9454 => "11111111",
	9455 => "11111111",
	9456 => "11111111",
	9457 => "11111111",
	9458 => "11111111",
	9459 => "11111111",
	9460 => "11111111",
	9461 => "11111111",
	9462 => "11111111",
	9463 => "11111111",
	9472 => "11111111",
	9473 => "11111111",
	9474 => "11111111",
	9475 => "11111111",
	9476 => "11111111",
	9477 => "11111111",
	9478 => "11111111",
	9479 => "11111111",
	9480 => "11111111",
	9481 => "11111111",
	9482 => "11111111",
	9483 => "11111111",
	9484 => "11111111",
	9485 => "11111111",
	9486 => "11111111",
	9487 => "11111111",
	9488 => "11111111",
	9489 => "11111111",
	9490 => "11111111",
	9491 => "11111111",
	9492 => "11111111",
	9493 => "11111111",
	9494 => "11111111",
	9495 => "11111111",
	9496 => "11111111",
	9497 => "11111111",
	9498 => "11111111",
	9499 => "11111111",
	9500 => "11111111",
	9501 => "11111111",
	9502 => "11111111",
	9503 => "11111111",
	9504 => "11111111",
	9505 => "11111111",
	9506 => "11111111",
	9507 => "11111111",
	9508 => "11111111",
	9509 => "11111111",
	9510 => "11111111",
	9511 => "11111111",
	9512 => "11111111",
	9513 => "11111111",
	9514 => "11111111",
	9515 => "11111111",
	9516 => "11111111",
	9517 => "11111111",
	9518 => "11111111",
	9519 => "11111111",
	9520 => "11111111",
	9521 => "11111111",
	9522 => "11111111",
	9523 => "11111111",
	9524 => "11111111",
	9525 => "11111111",
	9526 => "11111111",
	9527 => "11111111",
	9528 => "11111111",
	9529 => "11111111",
	9530 => "11111111",
	9531 => "11111111",
	9532 => "11111111",
	9533 => "11111111",
	9534 => "11111111",
	9535 => "11111111",
	9536 => "11111111",
	9537 => "11111111",
	9538 => "11111111",
	9539 => "11111111",
	9540 => "11111111",
	9541 => "11111111",
	9542 => "11111111",
	9543 => "11111111",
	9544 => "11111111",
	9545 => "11111111",
	9546 => "11111111",
	9547 => "11111111",
	9548 => "11111111",
	9549 => "11111111",
	9550 => "11111111",
	9551 => "11111111",
	9552 => "11111111",
	9553 => "11111111",
	9554 => "11111111",
	9555 => "11111111",
	9556 => "11111111",
	9557 => "11111111",
	9558 => "11111111",
	9559 => "11111111",
	9560 => "11111111",
	9561 => "11111111",
	9562 => "11111111",
	9563 => "11111111",
	9564 => "11111111",
	9565 => "11111111",
	9566 => "11111111",
	9567 => "11111111",
	9568 => "11111111",
	9569 => "11111111",
	9570 => "11111111",
	9571 => "11111111",
	9572 => "11111111",
	9573 => "11111111",
	9574 => "11111111",
	9575 => "11111111",
	9576 => "11111111",
	9577 => "11111111",
	9578 => "11111111",
	9579 => "11111111",
	9580 => "11111111",
	9581 => "11111111",
	9582 => "11111111",
	9583 => "11111111",
	9584 => "11111111",
	9585 => "11111111",
	9586 => "11111111",
	9587 => "11111111",
	9588 => "11111111",
	9589 => "11111111",
	9590 => "11111111",
	9591 => "11111111",
	9600 => "11111111",
	9601 => "11111111",
	9602 => "11111111",
	9603 => "11111111",
	9604 => "11111111",
	9605 => "11111111",
	9606 => "11111111",
	9607 => "11111111",
	9608 => "11111111",
	9609 => "11111111",
	9610 => "11111111",
	9611 => "11111111",
	9612 => "11111111",
	9613 => "11111111",
	9614 => "11111111",
	9615 => "11111111",
	9616 => "11111111",
	9617 => "11111111",
	9618 => "11111111",
	9619 => "11111111",
	9620 => "11111111",
	9621 => "11111111",
	9622 => "11111111",
	9623 => "11111111",
	9624 => "11111111",
	9625 => "11111111",
	9626 => "11111111",
	9627 => "11111111",
	9628 => "11111111",
	9629 => "11111111",
	9630 => "11111111",
	9631 => "11111111",
	9632 => "11111111",
	9633 => "11111111",
	9634 => "11111111",
	9635 => "11111111",
	9636 => "11111111",
	9637 => "11111111",
	9638 => "11111111",
	9639 => "11111111",
	9640 => "11111111",
	9641 => "11111111",
	9642 => "11111111",
	9643 => "11111111",
	9644 => "11111111",
	9645 => "11111111",
	9646 => "11111111",
	9647 => "11111111",
	9648 => "11111111",
	9649 => "11111111",
	9650 => "11111111",
	9651 => "11111111",
	9652 => "11111111",
	9653 => "11111111",
	9654 => "11111111",
	9655 => "11111111",
	9656 => "11111111",
	9657 => "11111111",
	9658 => "11111111",
	9659 => "11111111",
	9660 => "11111111",
	9661 => "11111111",
	9662 => "11111111",
	9663 => "11111111",
	9664 => "11111111",
	9665 => "11111111",
	9666 => "11111111",
	9667 => "11111111",
	9668 => "11111111",
	9669 => "11111111",
	9670 => "11111111",
	9671 => "11111111",
	9672 => "11111111",
	9673 => "11111111",
	9674 => "11111111",
	9675 => "11111111",
	9676 => "11111111",
	9677 => "11111111",
	9678 => "11111111",
	9679 => "11111111",
	9680 => "11111111",
	9681 => "11111111",
	9682 => "11111111",
	9683 => "11111111",
	9684 => "11111111",
	9685 => "11111111",
	9686 => "11111111",
	9687 => "11111111",
	9688 => "11111111",
	9689 => "11111111",
	9690 => "11111111",
	9691 => "11111111",
	9692 => "11111111",
	9693 => "11111111",
	9694 => "11111111",
	9695 => "11111111",
	9696 => "11111111",
	9697 => "11111111",
	9698 => "11111111",
	9699 => "11111111",
	9700 => "11111111",
	9701 => "11111111",
	9702 => "11111111",
	9703 => "11111111",
	9704 => "11111111",
	9705 => "11111111",
	9706 => "11111111",
	9707 => "11111111",
	9708 => "11111111",
	9709 => "11111111",
	9710 => "11111111",
	9711 => "11111111",
	9712 => "11111111",
	9713 => "11111111",
	9714 => "11111111",
	9715 => "11111111",
	9716 => "11111111",
	9717 => "11111111",
	9718 => "11111111",
	9719 => "11111111",
	9728 => "11111111",
	9729 => "11111111",
	9730 => "11111111",
	9731 => "11111111",
	9732 => "11111111",
	9733 => "11111111",
	9734 => "11111111",
	9735 => "11111111",
	9736 => "11111111",
	9737 => "11111111",
	9738 => "11111111",
	9739 => "11111111",
	9740 => "11111111",
	9741 => "11111111",
	9742 => "11111111",
	9743 => "11111111",
	9744 => "11111111",
	9745 => "11111111",
	9746 => "11111111",
	9747 => "11111111",
	9748 => "11111111",
	9749 => "11111111",
	9750 => "11111111",
	9751 => "11111111",
	9752 => "11111111",
	9753 => "11111111",
	9754 => "11111111",
	9755 => "11111111",
	9756 => "11111111",
	9757 => "11111111",
	9758 => "11111111",
	9759 => "11111111",
	9760 => "11111111",
	9761 => "11111111",
	9762 => "11111111",
	9763 => "11111111",
	9764 => "11111111",
	9765 => "11111111",
	9766 => "11111111",
	9767 => "11111111",
	9768 => "11111111",
	9769 => "11111111",
	9770 => "11111111",
	9771 => "11111111",
	9772 => "11111111",
	9773 => "11111111",
	9774 => "11111111",
	9775 => "11111111",
	9776 => "11111111",
	9777 => "11111111",
	9778 => "11111111",
	9779 => "11111111",
	9780 => "11111111",
	9781 => "11111111",
	9782 => "11111111",
	9783 => "11111111",
	9784 => "11111111",
	9785 => "11111111",
	9786 => "11111111",
	9787 => "11111111",
	9788 => "11111111",
	9789 => "11111111",
	9790 => "11111111",
	9791 => "11111111",
	9792 => "11111111",
	9793 => "11111111",
	9794 => "11111111",
	9795 => "11111111",
	9796 => "11111111",
	9797 => "11111111",
	9798 => "11111111",
	9799 => "11111111",
	9800 => "11111111",
	9801 => "11111111",
	9802 => "11111111",
	9803 => "11111111",
	9804 => "11111111",
	9805 => "11111111",
	9806 => "11111111",
	9807 => "11111111",
	9808 => "11111111",
	9809 => "11111111",
	9810 => "11111111",
	9811 => "11111111",
	9812 => "11111111",
	9813 => "11111111",
	9814 => "11111111",
	9815 => "11111111",
	9816 => "11111111",
	9817 => "11111111",
	9818 => "11111111",
	9819 => "11111111",
	9820 => "11111111",
	9821 => "11111111",
	9822 => "11111111",
	9823 => "11111111",
	9824 => "11111111",
	9825 => "11111111",
	9826 => "11111111",
	9827 => "11111111",
	9828 => "11111111",
	9829 => "11111111",
	9830 => "11111111",
	9831 => "11111111",
	9832 => "11111111",
	9833 => "11111111",
	9834 => "11111111",
	9835 => "11111111",
	9836 => "11111111",
	9837 => "11111111",
	9838 => "11111111",
	9839 => "11111111",
	9840 => "11111111",
	9841 => "11111111",
	9842 => "11111111",
	9843 => "11111111",
	9844 => "11111111",
	9845 => "11111111",
	9846 => "11111111",
	9847 => "11111111",
	9856 => "11111111",
	9857 => "11111111",
	9858 => "11111111",
	9859 => "11111111",
	9860 => "11111111",
	9861 => "11111111",
	9862 => "11111111",
	9863 => "11111111",
	9864 => "11111111",
	9865 => "11111111",
	9866 => "11111111",
	9867 => "11111111",
	9868 => "11111111",
	9869 => "11111111",
	9870 => "11111111",
	9871 => "11111111",
	9872 => "11111111",
	9873 => "11111111",
	9874 => "11111111",
	9875 => "11111111",
	9876 => "11111111",
	9877 => "11111111",
	9878 => "11111111",
	9879 => "11111111",
	9880 => "11111111",
	9881 => "11111111",
	9882 => "11111111",
	9883 => "11111111",
	9884 => "11111111",
	9885 => "11111111",
	9886 => "11111111",
	9887 => "11111111",
	9888 => "11111111",
	9889 => "11111111",
	9890 => "11111111",
	9891 => "11111111",
	9892 => "11111111",
	9893 => "11111111",
	9894 => "11111111",
	9895 => "11111111",
	9896 => "11111111",
	9897 => "11111111",
	9898 => "11111111",
	9899 => "11111111",
	9900 => "11111111",
	9901 => "11111111",
	9902 => "11111111",
	9903 => "11111111",
	9904 => "11111111",
	9905 => "11111111",
	9906 => "11111111",
	9907 => "11111111",
	9908 => "11111111",
	9909 => "11111111",
	9910 => "11111111",
	9911 => "11111111",
	9912 => "11111111",
	9913 => "11111111",
	9914 => "11111111",
	9915 => "11111111",
	9916 => "11111111",
	9917 => "11111111",
	9918 => "11111111",
	9919 => "11111111",
	9920 => "11111111",
	9921 => "11111111",
	9922 => "11111111",
	9923 => "11111111",
	9924 => "11111111",
	9925 => "11111111",
	9926 => "11111111",
	9927 => "11111111",
	9928 => "11111111",
	9929 => "11111111",
	9930 => "11111111",
	9931 => "11111111",
	9932 => "11111111",
	9933 => "11111111",
	9934 => "11111111",
	9935 => "11111111",
	9936 => "11111111",
	9937 => "11111111",
	9938 => "11111111",
	9939 => "11111111",
	9940 => "11111111",
	9941 => "11111111",
	9942 => "11111111",
	9943 => "11111111",
	9944 => "11111111",
	9945 => "11111111",
	9946 => "11111111",
	9947 => "11111111",
	9948 => "11111111",
	9949 => "11111111",
	9950 => "11111111",
	9951 => "11111111",
	9952 => "11111111",
	9953 => "11111111",
	9954 => "11111111",
	9955 => "11111111",
	9956 => "11111111",
	9957 => "11111111",
	9958 => "11111111",
	9959 => "11111111",
	9960 => "11111111",
	9961 => "11111111",
	9962 => "11111111",
	9963 => "11111111",
	9964 => "11111111",
	9965 => "11111111",
	9966 => "11111111",
	9967 => "11111111",
	9968 => "11111111",
	9969 => "11111111",
	9970 => "11111111",
	9971 => "11111111",
	9972 => "11111111",
	9973 => "11111111",
	9974 => "11111111",
	9975 => "11111111",
	9984 => "11111111",
	9985 => "11111111",
	9986 => "11111111",
	9987 => "11111111",
	9988 => "11111111",
	9989 => "11111111",
	9990 => "11111111",
	9991 => "11111111",
	9992 => "11111111",
	9993 => "11111111",
	9994 => "11111111",
	9995 => "11111111",
	9996 => "11111111",
	9997 => "11111111",
	9998 => "11111111",
	9999 => "11111111",
	10000 => "11111111",
	10001 => "11111111",
	10002 => "11111111",
	10003 => "11111111",
	10004 => "11111111",
	10005 => "11111111",
	10006 => "11111111",
	10007 => "11111111",
	10008 => "11111111",
	10009 => "11111111",
	10010 => "11111111",
	10011 => "11111111",
	10012 => "11111111",
	10013 => "11111111",
	10014 => "11111111",
	10015 => "11111111",
	10016 => "11111111",
	10017 => "11111111",
	10018 => "11111111",
	10019 => "11111111",
	10020 => "11111111",
	10021 => "11111111",
	10022 => "11111111",
	10023 => "11111111",
	10024 => "11111111",
	10025 => "11111111",
	10026 => "11111111",
	10027 => "11111111",
	10028 => "11111111",
	10029 => "11111111",
	10030 => "11111111",
	10031 => "11111111",
	10032 => "11111111",
	10033 => "11111111",
	10034 => "11111111",
	10035 => "11111111",
	10036 => "11111111",
	10037 => "11111111",
	10038 => "11111111",
	10039 => "11111111",
	10040 => "11111111",
	10041 => "11111111",
	10042 => "11111111",
	10043 => "11111111",
	10044 => "11111111",
	10045 => "11111111",
	10046 => "11111111",
	10047 => "11111111",
	10048 => "11111111",
	10049 => "11111111",
	10050 => "11111111",
	10051 => "11111111",
	10052 => "11111111",
	10053 => "11111111",
	10054 => "11111111",
	10055 => "11111111",
	10056 => "11111111",
	10057 => "11111111",
	10058 => "11111111",
	10059 => "11111111",
	10060 => "11111111",
	10061 => "11111111",
	10062 => "11111111",
	10063 => "11111111",
	10064 => "11111111",
	10065 => "11111111",
	10066 => "11111111",
	10067 => "11111111",
	10068 => "11111111",
	10069 => "11111111",
	10070 => "11111111",
	10071 => "11111111",
	10072 => "11111111",
	10073 => "11111111",
	10074 => "11111111",
	10075 => "11111111",
	10076 => "11111111",
	10077 => "11111111",
	10078 => "11111111",
	10079 => "11111111",
	10080 => "11111111",
	10081 => "11111111",
	10082 => "11111111",
	10083 => "11111111",
	10084 => "11111111",
	10085 => "11111111",
	10086 => "11111111",
	10087 => "11111111",
	10088 => "11111111",
	10089 => "11111111",
	10090 => "11111111",
	10091 => "11111111",
	10092 => "11111111",
	10093 => "11111111",
	10094 => "11111111",
	10095 => "11111111",
	10096 => "11111111",
	10097 => "11111111",
	10098 => "11111111",
	10099 => "11111111",
	10100 => "11111111",
	10101 => "11111111",
	10102 => "11111111",
	10103 => "11111111",
	10112 => "11111111",
	10113 => "11111111",
	10114 => "11111111",
	10115 => "11111111",
	10116 => "11111111",
	10117 => "11111111",
	10118 => "11111111",
	10119 => "11111111",
	10120 => "11111111",
	10121 => "11111111",
	10122 => "11111111",
	10123 => "11111111",
	10124 => "11111111",
	10125 => "11111111",
	10126 => "11111111",
	10127 => "11111111",
	10128 => "11111111",
	10129 => "11111111",
	10130 => "11111111",
	10131 => "11111111",
	10132 => "11111111",
	10133 => "11111111",
	10134 => "11111111",
	10135 => "11111111",
	10136 => "11111111",
	10137 => "11111111",
	10138 => "11111111",
	10139 => "11111111",
	10140 => "11111111",
	10141 => "11111111",
	10142 => "11111111",
	10143 => "11111111",
	10144 => "11111111",
	10145 => "11111111",
	10146 => "11111111",
	10147 => "11111111",
	10148 => "11111111",
	10149 => "11111111",
	10150 => "11111111",
	10151 => "11111111",
	10152 => "11111111",
	10153 => "11111111",
	10154 => "11111111",
	10155 => "11111111",
	10156 => "11111111",
	10157 => "11111111",
	10158 => "11111111",
	10159 => "11111111",
	10160 => "11111111",
	10161 => "11111111",
	10162 => "11111111",
	10163 => "11111111",
	10164 => "11111111",
	10165 => "11111111",
	10166 => "11111111",
	10167 => "11111111",
	10168 => "11111111",
	10169 => "11111111",
	10170 => "11111111",
	10171 => "11111111",
	10172 => "11111111",
	10173 => "11111111",
	10174 => "11111111",
	10175 => "11111111",
	10176 => "11111111",
	10177 => "11111111",
	10178 => "11111111",
	10179 => "11111111",
	10180 => "11111111",
	10181 => "11111111",
	10182 => "11111111",
	10183 => "11111111",
	10184 => "11111111",
	10185 => "11111111",
	10186 => "11111111",
	10187 => "11111111",
	10188 => "11111111",
	10189 => "11111111",
	10190 => "11111111",
	10191 => "11111111",
	10192 => "11111111",
	10193 => "11111111",
	10194 => "11111111",
	10195 => "11111111",
	10196 => "11111111",
	10197 => "11111111",
	10198 => "11111111",
	10199 => "11111111",
	10200 => "11111111",
	10201 => "11111111",
	10202 => "11111111",
	10203 => "11111111",
	10204 => "11111111",
	10205 => "11111111",
	10206 => "11111111",
	10207 => "11111111",
	10208 => "11111111",
	10209 => "11111111",
	10210 => "11111111",
	10211 => "11111111",
	10212 => "11111111",
	10213 => "11111111",
	10214 => "11111111",
	10215 => "11111111",
	10216 => "11111111",
	10217 => "11111111",
	10218 => "11111111",
	10219 => "11111111",
	10220 => "11111111",
	10221 => "11111111",
	10222 => "11111111",
	10223 => "11111111",
	10224 => "11111111",
	10225 => "11111111",
	10226 => "11111111",
	10227 => "11111111",
	10228 => "11111111",
	10229 => "11111111",
	10230 => "11111111",
	10231 => "11111111",
	10240 => "11111111",
	10241 => "11111111",
	10242 => "11111111",
	10243 => "11111111",
	10244 => "11111111",
	10245 => "11111111",
	10246 => "11111111",
	10247 => "11111111",
	10248 => "11111111",
	10249 => "11111111",
	10250 => "11111111",
	10251 => "11111111",
	10252 => "11111111",
	10253 => "11111111",
	10254 => "11111111",
	10255 => "11111111",
	10256 => "11111111",
	10257 => "11111111",
	10258 => "11111111",
	10259 => "11111111",
	10260 => "11111111",
	10261 => "11111111",
	10262 => "11111111",
	10263 => "11111111",
	10264 => "11111111",
	10265 => "11111111",
	10266 => "11111111",
	10267 => "11111111",
	10268 => "11111111",
	10269 => "11111111",
	10270 => "11111111",
	10271 => "11111111",
	10272 => "11111111",
	10273 => "11111111",
	10274 => "11111111",
	10275 => "11111111",
	10276 => "11111111",
	10277 => "11111111",
	10278 => "11111111",
	10279 => "11111111",
	10280 => "11111111",
	10281 => "11111111",
	10282 => "11111111",
	10283 => "11111111",
	10284 => "11111111",
	10285 => "11111111",
	10286 => "11111111",
	10287 => "11111111",
	10288 => "11111111",
	10289 => "11111111",
	10290 => "11111111",
	10291 => "11111111",
	10292 => "11111111",
	10293 => "11111111",
	10294 => "11111111",
	10295 => "11111111",
	10296 => "11111111",
	10297 => "11111111",
	10298 => "11111111",
	10299 => "11111111",
	10300 => "11111111",
	10301 => "11111111",
	10302 => "11111111",
	10303 => "11111111",
	10304 => "11111111",
	10305 => "11111111",
	10306 => "11111111",
	10307 => "11111111",
	10308 => "11111111",
	10309 => "11111111",
	10310 => "11111111",
	10311 => "11111111",
	10312 => "11111111",
	10313 => "11111111",
	10314 => "11111111",
	10315 => "11111111",
	10316 => "11111111",
	10317 => "11111111",
	10318 => "11111111",
	10319 => "11111111",
	10320 => "11111111",
	10321 => "11111111",
	10322 => "11111111",
	10323 => "11111111",
	10324 => "11111111",
	10325 => "11111111",
	10326 => "11111111",
	10327 => "11111111",
	10328 => "11111111",
	10329 => "11111111",
	10330 => "11111111",
	10331 => "11111111",
	10332 => "11111111",
	10333 => "11111111",
	10334 => "11111111",
	10335 => "11111111",
	10336 => "11111111",
	10337 => "11111111",
	10338 => "11111111",
	10339 => "11111111",
	10340 => "11111111",
	10341 => "11111111",
	10342 => "11111111",
	10343 => "11111111",
	10344 => "11111111",
	10345 => "11111111",
	10346 => "11111111",
	10347 => "11111111",
	10348 => "11111111",
	10349 => "11111111",
	10350 => "11111111",
	10351 => "11111111",
	10352 => "11111111",
	10353 => "11111111",
	10354 => "11111111",
	10355 => "11111111",
	10356 => "11111111",
	10357 => "11111111",
	10358 => "11111111",
	10359 => "11111111",
	10368 => "11111111",
	10369 => "11111111",
	10370 => "11111111",
	10371 => "11111111",
	10372 => "11111111",
	10373 => "11111111",
	10374 => "11111111",
	10375 => "11111111",
	10376 => "11111111",
	10377 => "11111111",
	10378 => "11111111",
	10379 => "11111111",
	10380 => "11111111",
	10381 => "11111111",
	10382 => "11111111",
	10383 => "11111111",
	10384 => "11111111",
	10385 => "11111111",
	10386 => "11111111",
	10387 => "11111111",
	10388 => "11111111",
	10389 => "11111111",
	10390 => "11111111",
	10391 => "11111111",
	10392 => "11111111",
	10393 => "11111111",
	10394 => "11111111",
	10395 => "11111111",
	10396 => "11111111",
	10397 => "11111111",
	10398 => "11111111",
	10399 => "11111111",
	10400 => "11111111",
	10401 => "11111111",
	10402 => "11111111",
	10403 => "11111111",
	10404 => "11111111",
	10405 => "11111111",
	10406 => "11111111",
	10407 => "11111111",
	10408 => "11111111",
	10409 => "11111111",
	10410 => "11111111",
	10411 => "11111111",
	10412 => "11111111",
	10413 => "11111111",
	10414 => "11111111",
	10415 => "11111111",
	10416 => "11111111",
	10417 => "11111111",
	10418 => "11111111",
	10419 => "11111111",
	10420 => "11111111",
	10421 => "11111111",
	10422 => "11111111",
	10423 => "11111111",
	10424 => "11111111",
	10425 => "11111111",
	10426 => "11111111",
	10427 => "11111111",
	10428 => "11111111",
	10429 => "11111111",
	10430 => "11111111",
	10431 => "11111111",
	10432 => "11111111",
	10433 => "11111111",
	10434 => "11111111",
	10435 => "11111111",
	10436 => "11111111",
	10437 => "11111111",
	10438 => "11111111",
	10439 => "11111111",
	10440 => "11111111",
	10441 => "11111111",
	10442 => "11111111",
	10443 => "11111111",
	10444 => "11111111",
	10445 => "11111111",
	10446 => "11111111",
	10447 => "11111111",
	10448 => "11111111",
	10449 => "11111111",
	10450 => "11111111",
	10451 => "11111111",
	10452 => "11111111",
	10453 => "11111111",
	10454 => "11111111",
	10455 => "11111111",
	10456 => "11111111",
	10457 => "11111111",
	10458 => "11111111",
	10459 => "11111111",
	10460 => "11111111",
	10461 => "11111111",
	10462 => "11111111",
	10463 => "11111111",
	10464 => "11111111",
	10465 => "11111111",
	10466 => "11111111",
	10467 => "11111111",
	10468 => "11111111",
	10469 => "11111111",
	10470 => "11111111",
	10471 => "11111111",
	10472 => "11111111",
	10473 => "11111111",
	10474 => "11111111",
	10475 => "11111111",
	10476 => "11111111",
	10477 => "11111111",
	10478 => "11111111",
	10479 => "11111111",
	10480 => "11111111",
	10481 => "11111111",
	10482 => "11111111",
	10483 => "11111111",
	10484 => "11111111",
	10485 => "11111111",
	10486 => "11111111",
	10487 => "11111111",
	10496 => "11111111",
	10497 => "11111111",
	10498 => "11111111",
	10499 => "11111111",
	10500 => "11111111",
	10501 => "11111111",
	10502 => "11111111",
	10503 => "11111111",
	10504 => "11111111",
	10505 => "11111111",
	10506 => "11111111",
	10507 => "11111111",
	10508 => "11111111",
	10509 => "11111111",
	10510 => "11111111",
	10511 => "11111111",
	10512 => "11111111",
	10513 => "11111111",
	10514 => "11111111",
	10515 => "11111111",
	10516 => "11111111",
	10517 => "11111111",
	10518 => "11111111",
	10519 => "11111111",
	10520 => "11111111",
	10521 => "11111111",
	10522 => "11111111",
	10523 => "11111111",
	10524 => "11111111",
	10525 => "11111111",
	10526 => "11111111",
	10527 => "11111111",
	10528 => "11111111",
	10529 => "11111111",
	10530 => "11111111",
	10531 => "11111111",
	10532 => "11111111",
	10533 => "11111111",
	10534 => "11111111",
	10535 => "11111111",
	10536 => "11111111",
	10537 => "11111111",
	10538 => "11111111",
	10539 => "11111111",
	10540 => "11111111",
	10541 => "11111111",
	10542 => "11111111",
	10543 => "11111111",
	10544 => "11111111",
	10545 => "11111111",
	10546 => "11111111",
	10547 => "11111111",
	10548 => "11111111",
	10549 => "11111111",
	10550 => "11111111",
	10551 => "11111111",
	10552 => "11111111",
	10553 => "11111111",
	10554 => "11111111",
	10555 => "11111111",
	10556 => "11111111",
	10557 => "11111111",
	10558 => "11111111",
	10559 => "11111111",
	10560 => "11111111",
	10561 => "11111111",
	10562 => "11111111",
	10563 => "11111111",
	10564 => "11111111",
	10565 => "11111111",
	10566 => "11111111",
	10567 => "11111111",
	10568 => "11111111",
	10569 => "11111111",
	10570 => "11111111",
	10571 => "11111111",
	10572 => "11111111",
	10573 => "11111111",
	10574 => "11111111",
	10575 => "11111111",
	10576 => "11111111",
	10577 => "11111111",
	10578 => "11111111",
	10579 => "11111111",
	10580 => "11111111",
	10581 => "11111111",
	10582 => "11111111",
	10583 => "11111111",
	10584 => "11111111",
	10585 => "11111111",
	10586 => "11111111",
	10587 => "11111111",
	10588 => "11111111",
	10589 => "11111111",
	10590 => "11111111",
	10591 => "11111111",
	10592 => "11111111",
	10593 => "11111111",
	10594 => "11111111",
	10595 => "11111111",
	10596 => "11111111",
	10597 => "11111111",
	10598 => "11111111",
	10599 => "11111111",
	10600 => "11111111",
	10601 => "11111111",
	10602 => "11111111",
	10603 => "11111111",
	10604 => "11111111",
	10605 => "11111111",
	10606 => "11111111",
	10607 => "11111111",
	10608 => "11111111",
	10609 => "11111111",
	10610 => "11111111",
	10611 => "11111111",
	10612 => "11111111",
	10613 => "11111111",
	10614 => "11111111",
	10615 => "11111111",
	10624 => "11111111",
	10625 => "11111111",
	10626 => "11111111",
	10627 => "11111111",
	10628 => "11111111",
	10629 => "11111111",
	10630 => "11111111",
	10631 => "11111111",
	10632 => "11111111",
	10633 => "11111111",
	10634 => "11111111",
	10635 => "11111111",
	10636 => "11111111",
	10637 => "11111111",
	10638 => "11111111",
	10639 => "11111111",
	10640 => "11111111",
	10641 => "11111111",
	10642 => "11111111",
	10643 => "11111111",
	10644 => "11111111",
	10645 => "11111111",
	10646 => "11111111",
	10647 => "11111111",
	10648 => "11111111",
	10649 => "11111111",
	10650 => "11111111",
	10651 => "11111111",
	10652 => "11111111",
	10653 => "11111111",
	10654 => "11111111",
	10655 => "11111111",
	10656 => "11111111",
	10657 => "11111111",
	10658 => "11111111",
	10659 => "11111111",
	10660 => "11111111",
	10661 => "11111111",
	10662 => "11111111",
	10663 => "11111111",
	10664 => "11111111",
	10665 => "11111111",
	10666 => "11111111",
	10667 => "11111111",
	10668 => "11111111",
	10669 => "11111111",
	10670 => "11111111",
	10671 => "11111111",
	10672 => "11111111",
	10673 => "11111111",
	10674 => "11111111",
	10675 => "11111111",
	10676 => "11111111",
	10677 => "11111111",
	10678 => "11111111",
	10679 => "11111111",
	10680 => "11111111",
	10681 => "11111111",
	10682 => "11111111",
	10683 => "11111111",
	10684 => "11111111",
	10685 => "11111111",
	10686 => "11111111",
	10687 => "11111111",
	10688 => "11111111",
	10689 => "11111111",
	10690 => "11111111",
	10691 => "11111111",
	10692 => "11111111",
	10693 => "11111111",
	10694 => "11111111",
	10695 => "11111111",
	10696 => "11111111",
	10697 => "11111111",
	10698 => "11111111",
	10699 => "11111111",
	10700 => "11111111",
	10701 => "11111111",
	10702 => "11111111",
	10703 => "11111111",
	10704 => "11111111",
	10705 => "11111111",
	10706 => "11111111",
	10707 => "11111111",
	10708 => "11111111",
	10709 => "11111111",
	10710 => "11111111",
	10711 => "11111111",
	10712 => "11111111",
	10713 => "11111111",
	10714 => "11111111",
	10715 => "11111111",
	10716 => "11111111",
	10717 => "11111111",
	10718 => "11111111",
	10719 => "11111111",
	10720 => "11111111",
	10721 => "11111111",
	10722 => "11111111",
	10723 => "11111111",
	10724 => "11111111",
	10725 => "11111111",
	10726 => "11111111",
	10727 => "11111111",
	10728 => "11111111",
	10729 => "11111111",
	10730 => "11111111",
	10731 => "11111111",
	10732 => "11111111",
	10733 => "11111111",
	10734 => "11111111",
	10735 => "11111111",
	10736 => "11111111",
	10737 => "11111111",
	10738 => "11111111",
	10739 => "11111111",
	10740 => "11111111",
	10741 => "11111111",
	10742 => "11111111",
	10743 => "11111111",
	10752 => "11111111",
	10753 => "11111111",
	10754 => "11111111",
	10755 => "11111111",
	10756 => "11111111",
	10757 => "11111111",
	10758 => "11111111",
	10759 => "11111111",
	10760 => "11111111",
	10761 => "11111111",
	10762 => "11111111",
	10763 => "11111111",
	10764 => "11111111",
	10765 => "11111111",
	10766 => "11111111",
	10767 => "11111111",
	10768 => "11111111",
	10769 => "11111111",
	10770 => "11111111",
	10771 => "11111111",
	10772 => "11111111",
	10773 => "11111111",
	10774 => "11111111",
	10775 => "11111111",
	10776 => "11111111",
	10777 => "11111111",
	10778 => "11111111",
	10779 => "11111111",
	10780 => "11111111",
	10781 => "11111111",
	10782 => "11111111",
	10783 => "11111111",
	10784 => "11111111",
	10785 => "11111111",
	10786 => "11111111",
	10787 => "11111111",
	10788 => "11111111",
	10789 => "11111111",
	10790 => "11111111",
	10791 => "11111111",
	10792 => "11111111",
	10793 => "11111111",
	10794 => "11111111",
	10795 => "11111111",
	10796 => "11111111",
	10797 => "11111111",
	10798 => "11111111",
	10799 => "11111111",
	10800 => "11111111",
	10801 => "11111111",
	10802 => "11111111",
	10803 => "11111111",
	10804 => "11111111",
	10805 => "11111111",
	10806 => "11111111",
	10807 => "11111111",
	10808 => "11111111",
	10809 => "11111111",
	10810 => "11111111",
	10811 => "11111111",
	10812 => "11111111",
	10813 => "11111111",
	10814 => "11111111",
	10815 => "11111111",
	10816 => "11111111",
	10817 => "11111111",
	10818 => "11111111",
	10819 => "11111111",
	10820 => "11111111",
	10821 => "11111111",
	10822 => "11111111",
	10823 => "11111111",
	10824 => "11111111",
	10825 => "11111111",
	10826 => "11111111",
	10827 => "11111111",
	10828 => "11111111",
	10829 => "11111111",
	10830 => "11111111",
	10831 => "11111111",
	10832 => "11111111",
	10833 => "11111111",
	10834 => "11111111",
	10835 => "11111111",
	10836 => "11111111",
	10837 => "11111111",
	10838 => "11111111",
	10839 => "11111111",
	10840 => "11111111",
	10841 => "11111111",
	10842 => "11111111",
	10843 => "11111111",
	10844 => "11111111",
	10845 => "11111111",
	10846 => "11111111",
	10847 => "11111111",
	10848 => "11111111",
	10849 => "11111111",
	10850 => "11111111",
	10851 => "11111111",
	10852 => "11111111",
	10853 => "11111111",
	10854 => "11111111",
	10855 => "11111111",
	10856 => "11111111",
	10857 => "11111111",
	10858 => "11111111",
	10859 => "11111111",
	10860 => "11111111",
	10861 => "11111111",
	10862 => "11111111",
	10863 => "11111111",
	10864 => "11111111",
	10865 => "11111111",
	10866 => "11111111",
	10867 => "11111111",
	10868 => "11111111",
	10869 => "11111111",
	10870 => "11111111",
	10871 => "11111111",
	10880 => "11111111",
	10881 => "11111111",
	10882 => "11111111",
	10883 => "11111111",
	10884 => "11111111",
	10885 => "11111111",
	10886 => "11111111",
	10887 => "11111111",
	10888 => "11111111",
	10889 => "11111111",
	10890 => "11111111",
	10891 => "11111111",
	10892 => "11111111",
	10893 => "11111111",
	10894 => "11111111",
	10895 => "11111111",
	10896 => "11111111",
	10897 => "11111111",
	10898 => "11111111",
	10899 => "11111111",
	10900 => "11111111",
	10901 => "11111111",
	10902 => "11111111",
	10903 => "11111111",
	10904 => "11111111",
	10905 => "11111111",
	10906 => "11111111",
	10907 => "11111111",
	10908 => "11111111",
	10909 => "11111111",
	10910 => "11111111",
	10911 => "11111111",
	10912 => "11111111",
	10913 => "11111111",
	10914 => "11111111",
	10915 => "11111111",
	10916 => "11111111",
	10917 => "11111111",
	10918 => "11111111",
	10919 => "11111111",
	10920 => "11111111",
	10921 => "11111111",
	10922 => "11111111",
	10923 => "11111111",
	10924 => "11111111",
	10925 => "11111111",
	10926 => "11111111",
	10927 => "11111111",
	10928 => "11111111",
	10929 => "11111111",
	10930 => "11111111",
	10931 => "11111111",
	10932 => "11111111",
	10933 => "11111111",
	10934 => "11111111",
	10935 => "11111111",
	10936 => "11111111",
	10937 => "11111111",
	10938 => "11111111",
	10939 => "11111111",
	10940 => "11111111",
	10941 => "11111111",
	10942 => "11111111",
	10943 => "11111111",
	10944 => "11111111",
	10945 => "11111111",
	10946 => "11111111",
	10947 => "11111111",
	10948 => "11111111",
	10949 => "11111111",
	10950 => "11111111",
	10951 => "11111111",
	10952 => "11111111",
	10953 => "11111111",
	10954 => "11111111",
	10955 => "11111111",
	10956 => "11111111",
	10957 => "11111111",
	10958 => "11111111",
	10959 => "11111111",
	10960 => "11111111",
	10961 => "11111111",
	10962 => "11111111",
	10963 => "11111111",
	10964 => "11111111",
	10965 => "11111111",
	10966 => "11111111",
	10967 => "11111111",
	10968 => "11111111",
	10969 => "11111111",
	10970 => "11111111",
	10971 => "11111111",
	10972 => "11111111",
	10973 => "11111111",
	10974 => "11111111",
	10975 => "11111111",
	10976 => "11111111",
	10977 => "11111111",
	10978 => "11111111",
	10979 => "11111111",
	10980 => "11111111",
	10981 => "11111111",
	10982 => "11111111",
	10983 => "11111111",
	10984 => "11111111",
	10985 => "11111111",
	10986 => "11111111",
	10987 => "11111111",
	10988 => "11111111",
	10989 => "11111111",
	10990 => "11111111",
	10991 => "11111111",
	10992 => "11111111",
	10993 => "11111111",
	10994 => "11111111",
	10995 => "11111111",
	10996 => "11111111",
	10997 => "11111111",
	10998 => "11111111",
	10999 => "11111111",
	11008 => "11111111",
	11009 => "11111111",
	11010 => "11111111",
	11011 => "11111111",
	11012 => "11111111",
	11013 => "11111111",
	11014 => "11111111",
	11015 => "11111111",
	11016 => "11111111",
	11017 => "11111111",
	11018 => "11111111",
	11019 => "11111111",
	11020 => "11111111",
	11021 => "11111111",
	11022 => "11111111",
	11023 => "11111111",
	11024 => "11111111",
	11025 => "11111111",
	11026 => "11111111",
	11027 => "11111111",
	11028 => "11111111",
	11029 => "11111111",
	11030 => "11111111",
	11031 => "11111111",
	11032 => "11111111",
	11033 => "11111111",
	11034 => "11111111",
	11035 => "11111111",
	11036 => "11111111",
	11037 => "11111111",
	11038 => "11111111",
	11039 => "11111111",
	11040 => "11111111",
	11041 => "11111111",
	11042 => "11111111",
	11043 => "11111111",
	11044 => "11111111",
	11045 => "11111111",
	11046 => "11111111",
	11047 => "11111111",
	11048 => "11111111",
	11049 => "11111111",
	11050 => "11111111",
	11051 => "11111111",
	11052 => "11111111",
	11053 => "11111111",
	11054 => "11111111",
	11055 => "11111111",
	11056 => "11111111",
	11057 => "11111111",
	11058 => "11111111",
	11059 => "11111111",
	11060 => "11111111",
	11061 => "11111111",
	11062 => "11111111",
	11063 => "11111111",
	11064 => "11111111",
	11065 => "11111111",
	11066 => "11111111",
	11067 => "11111111",
	11068 => "11111111",
	11069 => "11111111",
	11070 => "11111111",
	11071 => "11111111",
	11072 => "11111111",
	11073 => "11111111",
	11074 => "11111111",
	11075 => "11111111",
	11076 => "11111111",
	11077 => "11111111",
	11078 => "11111111",
	11079 => "11111111",
	11080 => "11111111",
	11081 => "11111111",
	11082 => "11111111",
	11083 => "11111111",
	11084 => "11111111",
	11085 => "11111111",
	11086 => "11111111",
	11087 => "11111111",
	11088 => "11111111",
	11089 => "11111111",
	11090 => "11111111",
	11091 => "11111111",
	11092 => "11111111",
	11093 => "11111111",
	11094 => "11111111",
	11095 => "11111111",
	11096 => "11111111",
	11097 => "11111111",
	11098 => "11111111",
	11099 => "11111111",
	11100 => "11111111",
	11101 => "11111111",
	11102 => "11111111",
	11103 => "11111111",
	11104 => "11111111",
	11105 => "11111111",
	11106 => "11111111",
	11107 => "11111111",
	11108 => "11111111",
	11109 => "11111111",
	11110 => "11111111",
	11111 => "11111111",
	11112 => "11111111",
	11113 => "11111111",
	11114 => "11111111",
	11115 => "11111111",
	11116 => "11111111",
	11117 => "11111111",
	11118 => "11111111",
	11119 => "11111111",
	11120 => "11111111",
	11121 => "11111111",
	11122 => "11111111",
	11123 => "11111111",
	11124 => "11111111",
	11125 => "11111111",
	11126 => "11111111",
	11127 => "11111111",
	11136 => "11111111",
	11137 => "11111111",
	11138 => "11111111",
	11139 => "11111111",
	11140 => "11111111",
	11141 => "11111111",
	11142 => "11111111",
	11143 => "11111111",
	11144 => "11111111",
	11145 => "11111111",
	11146 => "11111111",
	11147 => "11111111",
	11148 => "11111111",
	11149 => "11111111",
	11150 => "11111111",
	11151 => "11111111",
	11152 => "11111111",
	11153 => "11111111",
	11154 => "11111111",
	11155 => "11111111",
	11156 => "11111111",
	11157 => "11111111",
	11158 => "11111111",
	11159 => "11111111",
	11160 => "11111111",
	11161 => "11111111",
	11162 => "11111111",
	11163 => "11111111",
	11164 => "11111111",
	11165 => "11111111",
	11166 => "11111111",
	11167 => "11111111",
	11168 => "11111111",
	11169 => "11111111",
	11170 => "11111111",
	11171 => "11111111",
	11172 => "11111111",
	11173 => "11111111",
	11174 => "11111111",
	11175 => "11111111",
	11176 => "11111111",
	11177 => "11111111",
	11178 => "11111111",
	11179 => "11111111",
	11180 => "11111111",
	11181 => "11111111",
	11182 => "11111111",
	11183 => "11111111",
	11184 => "11111111",
	11185 => "11111111",
	11186 => "11111111",
	11187 => "11111111",
	11188 => "11111111",
	11189 => "11111111",
	11190 => "11111111",
	11191 => "11111111",
	11192 => "11111111",
	11193 => "11111111",
	11194 => "11111111",
	11195 => "11111111",
	11196 => "11111111",
	11197 => "11111111",
	11198 => "11111111",
	11199 => "11111111",
	11200 => "11111111",
	11201 => "11111111",
	11202 => "11111111",
	11203 => "11111111",
	11204 => "11111111",
	11205 => "11111111",
	11206 => "11111111",
	11207 => "11111111",
	11208 => "11111111",
	11209 => "11111111",
	11210 => "11111111",
	11211 => "11111111",
	11212 => "11111111",
	11213 => "11111111",
	11214 => "11111111",
	11215 => "11111111",
	11216 => "11111111",
	11217 => "11111111",
	11218 => "11111111",
	11219 => "11111111",
	11220 => "11111111",
	11221 => "11111111",
	11222 => "11111111",
	11223 => "11111111",
	11224 => "11111111",
	11225 => "11111111",
	11226 => "11111111",
	11227 => "11111111",
	11228 => "11111111",
	11229 => "11111111",
	11230 => "11111111",
	11231 => "11111111",
	11232 => "11111111",
	11233 => "11111111",
	11234 => "11111111",
	11235 => "11111111",
	11236 => "11111111",
	11237 => "11111111",
	11238 => "11111111",
	11239 => "11111111",
	11240 => "11111111",
	11241 => "11111111",
	11242 => "11111111",
	11243 => "11111111",
	11244 => "11111111",
	11245 => "11111111",
	11246 => "11111111",
	11247 => "11111111",
	11248 => "11111111",
	11249 => "11111111",
	11250 => "11111111",
	11251 => "11111111",
	11252 => "11111111",
	11253 => "11111111",
	11254 => "11111111",
	11255 => "11111111",
	11264 => "11111111",
	11265 => "11111111",
	11266 => "11111111",
	11267 => "11111111",
	11268 => "11111111",
	11269 => "11111111",
	11270 => "11111111",
	11271 => "11111111",
	11272 => "11111111",
	11273 => "11111111",
	11274 => "11111111",
	11275 => "11111111",
	11276 => "11111111",
	11277 => "11111111",
	11278 => "11111111",
	11279 => "11111111",
	11280 => "11111111",
	11281 => "11111111",
	11282 => "11111111",
	11283 => "11111111",
	11284 => "11111111",
	11285 => "11111111",
	11286 => "11111111",
	11287 => "11111111",
	11288 => "11111111",
	11289 => "11111111",
	11290 => "11111111",
	11291 => "11111111",
	11292 => "11111111",
	11293 => "11111111",
	11294 => "11111111",
	11295 => "11111111",
	11296 => "11111111",
	11297 => "11111111",
	11298 => "11111111",
	11299 => "11111111",
	11300 => "11111111",
	11301 => "11111111",
	11302 => "11111111",
	11303 => "11111111",
	11304 => "11111111",
	11305 => "11111111",
	11306 => "11111111",
	11307 => "11111111",
	11308 => "11111111",
	11309 => "11111111",
	11310 => "11111111",
	11311 => "11111111",
	11312 => "11111111",
	11313 => "11111111",
	11314 => "11111111",
	11315 => "11111111",
	11316 => "11111111",
	11317 => "11111111",
	11318 => "11111111",
	11319 => "11111111",
	11320 => "11111111",
	11321 => "11111111",
	11322 => "11111111",
	11323 => "11111111",
	11324 => "11111111",
	11325 => "11111111",
	11326 => "11111111",
	11327 => "11111111",
	11328 => "11111111",
	11329 => "11111111",
	11330 => "11111111",
	11331 => "11111111",
	11332 => "11111111",
	11333 => "11111111",
	11334 => "11111111",
	11335 => "11111111",
	11336 => "11111111",
	11337 => "11111111",
	11338 => "11111111",
	11339 => "11111111",
	11340 => "11111111",
	11341 => "11111111",
	11342 => "11111111",
	11343 => "11111111",
	11344 => "11111111",
	11345 => "11111111",
	11346 => "11111111",
	11347 => "11111111",
	11348 => "11111111",
	11349 => "11111111",
	11350 => "11111111",
	11351 => "11111111",
	11352 => "11111111",
	11353 => "11111111",
	11354 => "11111111",
	11355 => "11111111",
	11356 => "11111111",
	11357 => "11111111",
	11358 => "11111111",
	11359 => "11111111",
	11360 => "11111111",
	11361 => "11111111",
	11362 => "11111111",
	11363 => "11111111",
	11364 => "11111111",
	11365 => "11111111",
	11366 => "11111111",
	11367 => "11111111",
	11368 => "11111111",
	11369 => "11111111",
	11370 => "11111111",
	11371 => "11111111",
	11372 => "11111111",
	11373 => "11111111",
	11374 => "11111111",
	11375 => "11111111",
	11376 => "11111111",
	11377 => "11111111",
	11378 => "11111111",
	11379 => "11111111",
	11380 => "11111111",
	11381 => "11111111",
	11382 => "11111111",
	11383 => "11111111",
	11392 => "11111111",
	11393 => "11111111",
	11394 => "11111111",
	11395 => "11111111",
	11396 => "11111111",
	11397 => "11111111",
	11398 => "11111111",
	11399 => "11111111",
	11400 => "11111111",
	11401 => "11111111",
	11402 => "11111111",
	11403 => "11111111",
	11404 => "11111111",
	11405 => "11111111",
	11406 => "11111111",
	11407 => "11111111",
	11408 => "11111111",
	11409 => "11111111",
	11410 => "11111111",
	11411 => "11111111",
	11412 => "11111111",
	11413 => "11111111",
	11414 => "11111111",
	11415 => "11111111",
	11416 => "11111111",
	11417 => "11111111",
	11418 => "11111111",
	11419 => "11111111",
	11420 => "11111111",
	11421 => "11111111",
	11422 => "11111111",
	11423 => "11111111",
	11424 => "11111111",
	11425 => "11111111",
	11426 => "11111111",
	11427 => "11111111",
	11428 => "11111111",
	11429 => "11111111",
	11430 => "11111111",
	11431 => "11111111",
	11432 => "11111111",
	11433 => "11111111",
	11434 => "11111111",
	11435 => "11111111",
	11436 => "11111111",
	11437 => "11111111",
	11438 => "11111111",
	11439 => "11111111",
	11440 => "11111111",
	11441 => "11111111",
	11442 => "11111111",
	11443 => "11111111",
	11444 => "11111111",
	11445 => "11111111",
	11446 => "11111111",
	11447 => "11111111",
	11448 => "11111111",
	11449 => "11111111",
	11450 => "11111111",
	11451 => "11111111",
	11452 => "11111111",
	11453 => "11111111",
	11454 => "11111111",
	11455 => "11111111",
	11456 => "11111111",
	11457 => "11111111",
	11458 => "11111111",
	11459 => "11111111",
	11460 => "11111111",
	11461 => "11111111",
	11462 => "11111111",
	11463 => "11111111",
	11464 => "11111111",
	11465 => "11111111",
	11466 => "11111111",
	11467 => "11111111",
	11468 => "11111111",
	11469 => "11111111",
	11470 => "11111111",
	11471 => "11111111",
	11472 => "11111111",
	11473 => "11111111",
	11474 => "11111111",
	11475 => "11111111",
	11476 => "11111111",
	11477 => "11111111",
	11478 => "11111111",
	11479 => "11111111",
	11480 => "11111111",
	11481 => "11111111",
	11482 => "11111111",
	11483 => "11111111",
	11484 => "11111111",
	11485 => "11111111",
	11486 => "11111111",
	11487 => "11111111",
	11488 => "11111111",
	11489 => "11111111",
	11490 => "11111111",
	11491 => "11111111",
	11492 => "11111111",
	11493 => "11111111",
	11494 => "11111111",
	11495 => "11111111",
	11496 => "11111111",
	11497 => "11111111",
	11498 => "11111111",
	11499 => "11111111",
	11500 => "11111111",
	11501 => "11111111",
	11502 => "11111111",
	11503 => "11111111",
	11504 => "11111111",
	11505 => "11111111",
	11506 => "11111111",
	11507 => "11111111",
	11508 => "11111111",
	11509 => "11111111",
	11510 => "11111111",
	11511 => "11111111",
	11520 => "11111111",
	11521 => "11111111",
	11522 => "11111111",
	11523 => "11111111",
	11524 => "11111111",
	11525 => "11111111",
	11526 => "11111111",
	11527 => "11111111",
	11528 => "11111111",
	11529 => "11111111",
	11530 => "11111111",
	11531 => "11111111",
	11532 => "11111111",
	11533 => "11111111",
	11534 => "11111111",
	11535 => "11111111",
	11536 => "11111111",
	11537 => "11111111",
	11538 => "11111111",
	11539 => "11111111",
	11540 => "11111111",
	11541 => "11111111",
	11542 => "11111111",
	11543 => "11111111",
	11544 => "11111111",
	11545 => "11111111",
	11546 => "11111111",
	11547 => "11111111",
	11548 => "11111111",
	11549 => "11111111",
	11550 => "11111111",
	11551 => "11111111",
	11552 => "11111111",
	11553 => "11111111",
	11554 => "11111111",
	11555 => "11111111",
	11556 => "11111111",
	11557 => "11111111",
	11558 => "11111111",
	11559 => "11111111",
	11560 => "11111111",
	11561 => "11111111",
	11562 => "11111111",
	11563 => "11111111",
	11564 => "11111111",
	11565 => "11111111",
	11566 => "11111111",
	11567 => "11111111",
	11568 => "11111111",
	11569 => "11111111",
	11570 => "11111111",
	11571 => "11111111",
	11572 => "11111111",
	11573 => "11111111",
	11574 => "11111111",
	11575 => "11111111",
	11576 => "11111111",
	11577 => "11111111",
	11578 => "11111111",
	11579 => "11111111",
	11580 => "11111111",
	11581 => "11111111",
	11582 => "11111111",
	11583 => "11111111",
	11584 => "11111111",
	11585 => "11111111",
	11586 => "11111111",
	11587 => "11111111",
	11588 => "11111111",
	11589 => "11111111",
	11590 => "11111111",
	11591 => "11111111",
	11592 => "11111111",
	11593 => "11111111",
	11594 => "11111111",
	11595 => "11111111",
	11596 => "11111111",
	11597 => "11111111",
	11598 => "11111111",
	11599 => "11111111",
	11600 => "11111111",
	11601 => "11111111",
	11602 => "11111111",
	11603 => "11111111",
	11604 => "11111111",
	11605 => "11111111",
	11606 => "11111111",
	11607 => "11111111",
	11608 => "11111111",
	11609 => "11111111",
	11610 => "11111111",
	11611 => "11111111",
	11612 => "11111111",
	11613 => "11111111",
	11614 => "11111111",
	11615 => "11111111",
	11616 => "11111111",
	11617 => "11111111",
	11618 => "11111111",
	11619 => "11111111",
	11620 => "11111111",
	11621 => "11111111",
	11622 => "11111111",
	11623 => "11111111",
	11624 => "11111111",
	11625 => "11111111",
	11626 => "11111111",
	11627 => "11111111",
	11628 => "11111111",
	11629 => "11111111",
	11630 => "11111111",
	11631 => "11111111",
	11632 => "11111111",
	11633 => "11111111",
	11634 => "11111111",
	11635 => "11111111",
	11636 => "11111111",
	11637 => "11111111",
	11638 => "11111111",
	11639 => "11111111",
	11648 => "11111111",
	11649 => "11111111",
	11650 => "11111111",
	11651 => "11111111",
	11652 => "11111111",
	11653 => "11111111",
	11654 => "11111111",
	11655 => "11111111",
	11656 => "11111111",
	11657 => "11111111",
	11658 => "11111111",
	11659 => "11111111",
	11660 => "11111111",
	11661 => "11111111",
	11662 => "11111111",
	11663 => "11111111",
	11664 => "11111111",
	11665 => "11111111",
	11666 => "11111111",
	11667 => "11111111",
	11668 => "11111111",
	11669 => "11111111",
	11670 => "11111111",
	11671 => "11111111",
	11672 => "11111111",
	11673 => "11111111",
	11674 => "11111111",
	11675 => "11111111",
	11676 => "11111111",
	11677 => "11111111",
	11678 => "11111111",
	11679 => "11111111",
	11680 => "11111111",
	11681 => "11111111",
	11682 => "11111111",
	11683 => "11111111",
	11684 => "11111111",
	11685 => "11111111",
	11686 => "11111111",
	11687 => "11111111",
	11688 => "11111111",
	11689 => "11111111",
	11690 => "11111111",
	11691 => "11111111",
	11692 => "11111111",
	11693 => "11111111",
	11694 => "11111111",
	11695 => "11111111",
	11696 => "11111111",
	11697 => "11111111",
	11698 => "11111111",
	11699 => "11111111",
	11700 => "11111111",
	11701 => "11111111",
	11702 => "11111111",
	11703 => "11111111",
	11704 => "11111111",
	11705 => "11111111",
	11706 => "11111111",
	11707 => "11111111",
	11708 => "11111111",
	11709 => "11111111",
	11710 => "11111111",
	11711 => "11111111",
	11712 => "11111111",
	11713 => "11111111",
	11714 => "11111111",
	11715 => "11111111",
	11716 => "11111111",
	11717 => "11111111",
	11718 => "11111111",
	11719 => "11111111",
	11720 => "11111111",
	11721 => "11111111",
	11722 => "11111111",
	11723 => "11111111",
	11724 => "11111111",
	11725 => "11111111",
	11726 => "11111111",
	11727 => "11111111",
	11728 => "11111111",
	11729 => "11111111",
	11730 => "11111111",
	11731 => "11111111",
	11732 => "11111111",
	11733 => "11111111",
	11734 => "11111111",
	11735 => "11111111",
	11736 => "11111111",
	11737 => "11111111",
	11738 => "11111111",
	11739 => "11111111",
	11740 => "11111111",
	11741 => "11111111",
	11742 => "11111111",
	11743 => "11111111",
	11744 => "11111111",
	11745 => "11111111",
	11746 => "11111111",
	11747 => "11111111",
	11748 => "11111111",
	11749 => "11111111",
	11750 => "11111111",
	11751 => "11111111",
	11752 => "11111111",
	11753 => "11111111",
	11754 => "11111111",
	11755 => "11111111",
	11756 => "11111111",
	11757 => "11111111",
	11758 => "11111111",
	11759 => "11111111",
	11760 => "11111111",
	11761 => "11111111",
	11762 => "11111111",
	11763 => "11111111",
	11764 => "11111111",
	11765 => "11111111",
	11766 => "11111111",
	11767 => "11111111",
	11776 => "11111111",
	11777 => "11111111",
	11778 => "11111111",
	11779 => "11111111",
	11780 => "11111111",
	11781 => "11111111",
	11782 => "11111111",
	11783 => "11111111",
	11784 => "11111111",
	11785 => "11111111",
	11786 => "11111111",
	11787 => "11111111",
	11788 => "11111111",
	11789 => "11111111",
	11790 => "11111111",
	11791 => "11111111",
	11792 => "11111111",
	11793 => "11111111",
	11794 => "11111111",
	11795 => "11111111",
	11796 => "11111111",
	11797 => "11111111",
	11798 => "11111111",
	11799 => "11111111",
	11800 => "11111111",
	11801 => "11111111",
	11802 => "11111111",
	11803 => "11111111",
	11804 => "11111111",
	11805 => "11111111",
	11806 => "11111111",
	11807 => "11111111",
	11808 => "11111111",
	11809 => "11111111",
	11810 => "11111111",
	11811 => "11111111",
	11812 => "11111111",
	11813 => "11111111",
	11814 => "11111111",
	11815 => "11111111",
	11816 => "11111111",
	11817 => "11111111",
	11818 => "11111111",
	11819 => "11111111",
	11820 => "11111111",
	11821 => "11111111",
	11822 => "11111111",
	11823 => "11111111",
	11824 => "11111111",
	11825 => "11111111",
	11826 => "11111111",
	11827 => "11111111",
	11828 => "11111111",
	11829 => "11111111",
	11830 => "11111111",
	11831 => "11111111",
	11832 => "11111111",
	11833 => "11111111",
	11834 => "11111111",
	11835 => "11111111",
	11836 => "11111111",
	11837 => "11111111",
	11838 => "11111111",
	11839 => "11111111",
	11840 => "11111111",
	11841 => "11111111",
	11842 => "11111111",
	11843 => "11111111",
	11844 => "11111111",
	11845 => "11111111",
	11846 => "11111111",
	11847 => "11111111",
	11848 => "11111111",
	11849 => "11111111",
	11850 => "11111111",
	11851 => "11111111",
	11852 => "11111111",
	11853 => "11111111",
	11854 => "11111111",
	11855 => "11111111",
	11856 => "11111111",
	11857 => "11111111",
	11858 => "11111111",
	11859 => "11111111",
	11860 => "11111111",
	11861 => "11111111",
	11862 => "11111111",
	11863 => "11111111",
	11864 => "11111111",
	11865 => "11111111",
	11866 => "11111111",
	11867 => "11111111",
	11868 => "11111111",
	11869 => "11111111",
	11870 => "11111111",
	11871 => "11111111",
	11872 => "11111111",
	11873 => "11111111",
	11874 => "11111111",
	11875 => "11111111",
	11876 => "11111111",
	11877 => "11111111",
	11878 => "11111111",
	11879 => "11111111",
	11880 => "11111111",
	11881 => "11111111",
	11882 => "11111111",
	11883 => "11111111",
	11884 => "11111111",
	11885 => "11111111",
	11886 => "11111111",
	11887 => "11111111",
	11888 => "11111111",
	11889 => "11111111",
	11890 => "11111111",
	11891 => "11111111",
	11892 => "11111111",
	11893 => "11111111",
	11894 => "11111111",
	11895 => "11111111",
	11904 => "11111111",
	11905 => "11111111",
	11906 => "11111111",
	11907 => "11111111",
	11908 => "11111111",
	11909 => "11111111",
	11910 => "11111111",
	11911 => "11111111",
	11912 => "11111111",
	11913 => "11111111",
	11914 => "11111111",
	11915 => "11111111",
	11916 => "11111111",
	11917 => "11111111",
	11918 => "11111111",
	11919 => "11111111",
	11920 => "11111111",
	11921 => "11111111",
	11922 => "11111111",
	11923 => "11111111",
	11924 => "11111111",
	11925 => "11111111",
	11926 => "11111111",
	11927 => "11111111",
	11928 => "11111111",
	11929 => "11111111",
	11930 => "11111111",
	11931 => "11111111",
	11932 => "11111111",
	11933 => "11111111",
	11934 => "11111111",
	11935 => "11111111",
	11936 => "11111111",
	11937 => "11111111",
	11938 => "11111111",
	11939 => "11111111",
	11940 => "11111111",
	11941 => "11111111",
	11942 => "11111111",
	11943 => "11111111",
	11944 => "11111111",
	11945 => "11111111",
	11946 => "11111111",
	11947 => "11111111",
	11948 => "11111111",
	11949 => "11111111",
	11950 => "11111111",
	11951 => "11111111",
	11952 => "11111111",
	11953 => "11111111",
	11954 => "11111111",
	11955 => "11111111",
	11956 => "11111111",
	11957 => "11111111",
	11958 => "11111111",
	11959 => "11111111",
	11960 => "11111111",
	11961 => "11111111",
	11962 => "11111111",
	11963 => "11111111",
	11964 => "11111111",
	11965 => "11111111",
	11966 => "11111111",
	11967 => "11111111",
	11968 => "11111111",
	11969 => "11111111",
	11970 => "11111111",
	11971 => "11111111",
	11972 => "11111111",
	11973 => "11111111",
	11974 => "11111111",
	11975 => "11111111",
	11976 => "11111111",
	11977 => "11111111",
	11978 => "11111111",
	11979 => "11111111",
	11980 => "11111111",
	11981 => "11111111",
	11982 => "11111111",
	11983 => "11111111",
	11984 => "11111111",
	11985 => "11111111",
	11986 => "11111111",
	11987 => "11111111",
	11988 => "11111111",
	11989 => "11111111",
	11990 => "11111111",
	11991 => "11111111",
	11992 => "11111111",
	11993 => "11111111",
	11994 => "11111111",
	11995 => "11111111",
	11996 => "11111111",
	11997 => "11111111",
	11998 => "11111111",
	11999 => "11111111",
	12000 => "11111111",
	12001 => "11111111",
	12002 => "11111111",
	12003 => "11111111",
	12004 => "11111111",
	12005 => "11111111",
	12006 => "11111111",
	12007 => "11111111",
	12008 => "11111111",
	12009 => "11111111",
	12010 => "11111111",
	12011 => "11111111",
	12012 => "11111111",
	12013 => "11111111",
	12014 => "11111111",
	12015 => "11111111",
	12016 => "11111111",
	12017 => "11111111",
	12018 => "11111111",
	12019 => "11111111",
	12020 => "11111111",
	12021 => "11111111",
	12022 => "11111111",
	12023 => "11111111",
	12032 => "11111111",
	12033 => "11111111",
	12034 => "11111111",
	12035 => "11111111",
	12036 => "11111111",
	12037 => "11111111",
	12038 => "11111111",
	12039 => "11111111",
	12040 => "11111111",
	12041 => "11111111",
	12042 => "11111111",
	12043 => "11111111",
	12044 => "11111111",
	12045 => "11111111",
	12046 => "11111111",
	12047 => "11111111",
	12048 => "11111111",
	12049 => "11111111",
	12050 => "11111111",
	12051 => "11111111",
	12052 => "11111111",
	12053 => "11111111",
	12054 => "11111111",
	12055 => "11111111",
	12056 => "11111111",
	12057 => "11111111",
	12058 => "11111111",
	12059 => "11111111",
	12060 => "11111111",
	12061 => "11111111",
	12062 => "11111111",
	12063 => "11111111",
	12064 => "11111111",
	12065 => "11111111",
	12066 => "11111111",
	12067 => "11111111",
	12068 => "11111111",
	12069 => "11111111",
	12070 => "11111111",
	12071 => "11111111",
	12072 => "11111111",
	12073 => "11111111",
	12074 => "11111111",
	12075 => "11111111",
	12076 => "11111111",
	12077 => "11111111",
	12078 => "11111111",
	12079 => "11111111",
	12080 => "11111111",
	12081 => "11111111",
	12082 => "11111111",
	12083 => "11111111",
	12084 => "11111111",
	12085 => "11111111",
	12086 => "11111111",
	12087 => "11111111",
	12088 => "11111111",
	12089 => "11111111",
	12090 => "11111111",
	12091 => "11111111",
	12092 => "11111111",
	12093 => "11111111",
	12094 => "11111111",
	12095 => "11111111",
	12096 => "11111111",
	12097 => "11111111",
	12098 => "11111111",
	12099 => "11111111",
	12100 => "11111111",
	12101 => "11111111",
	12102 => "11111111",
	12103 => "11111111",
	12104 => "11111111",
	12105 => "11111111",
	12106 => "11111111",
	12107 => "11111111",
	12108 => "11111111",
	12109 => "11111111",
	12110 => "11111111",
	12111 => "11111111",
	12112 => "11111111",
	12113 => "11111111",
	12114 => "11111111",
	12115 => "11111111",
	12116 => "11111111",
	12117 => "11111111",
	12118 => "11111111",
	12119 => "11111111",
	12120 => "11111111",
	12121 => "11111111",
	12122 => "11111111",
	12123 => "11111111",
	12124 => "11111111",
	12125 => "11111111",
	12126 => "11111111",
	12127 => "11111111",
	12128 => "11111111",
	12129 => "11111111",
	12130 => "11111111",
	12131 => "11111111",
	12132 => "11111111",
	12133 => "11111111",
	12134 => "11111111",
	12135 => "11111111",
	12136 => "11111111",
	12137 => "11111111",
	12138 => "11111111",
	12139 => "11111111",
	12140 => "11111111",
	12141 => "11111111",
	12142 => "11111111",
	12143 => "11111111",
	12144 => "11111111",
	12145 => "11111111",
	12146 => "11111111",
	12147 => "11111111",
	12148 => "11111111",
	12149 => "11111111",
	12150 => "11111111",
	12151 => "11111111",
	12160 => "11111111",
	12161 => "11111111",
	12162 => "11111111",
	12163 => "11111111",
	12164 => "11111111",
	12165 => "11111111",
	12166 => "11111111",
	12167 => "11111111",
	12168 => "11111111",
	12169 => "11111111",
	12170 => "11111111",
	12171 => "11111111",
	12172 => "11111111",
	12173 => "11111111",
	12174 => "11111111",
	12175 => "11111111",
	12176 => "11111111",
	12177 => "11111111",
	12178 => "11111111",
	12179 => "11111111",
	12180 => "11111111",
	12181 => "11111111",
	12182 => "11111111",
	12183 => "11111111",
	12184 => "11111111",
	12185 => "11111111",
	12186 => "11111111",
	12187 => "11111111",
	12188 => "11111111",
	12189 => "11111111",
	12190 => "11111111",
	12191 => "11111111",
	12192 => "11111111",
	12193 => "11111111",
	12194 => "11111111",
	12195 => "11111111",
	12196 => "11111111",
	12197 => "11111111",
	12198 => "11111111",
	12199 => "11111111",
	12200 => "11111111",
	12201 => "11111111",
	12202 => "11111111",
	12203 => "11111111",
	12204 => "11111111",
	12205 => "11111111",
	12206 => "11111111",
	12207 => "11111111",
	12208 => "11111111",
	12209 => "11111111",
	12210 => "11111111",
	12211 => "11111111",
	12212 => "11111111",
	12213 => "11111111",
	12214 => "11111111",
	12215 => "11111111",
	12216 => "11111111",
	12217 => "11111111",
	12218 => "11111111",
	12219 => "11111111",
	12220 => "11111111",
	12221 => "11111111",
	12222 => "11111111",
	12223 => "11111111",
	12224 => "11111111",
	12225 => "11111111",
	12226 => "11111111",
	12227 => "11111111",
	12228 => "11111111",
	12229 => "11111111",
	12230 => "11111111",
	12231 => "11111111",
	12232 => "11111111",
	12233 => "11111111",
	12234 => "11111111",
	12235 => "11111111",
	12236 => "11111111",
	12237 => "11111111",
	12238 => "11111111",
	12239 => "11111111",
	12240 => "11111111",
	12241 => "11111111",
	12242 => "11111111",
	12243 => "11111111",
	12244 => "11111111",
	12245 => "11111111",
	12246 => "11111111",
	12247 => "11111111",
	12248 => "11111111",
	12249 => "11111111",
	12250 => "11111111",
	12251 => "11111111",
	12252 => "11111111",
	12253 => "11111111",
	12254 => "11111111",
	12255 => "11111111",
	12256 => "11111111",
	12257 => "11111111",
	12258 => "11111111",
	12259 => "11111111",
	12260 => "11111111",
	12261 => "11111111",
	12262 => "11111111",
	12263 => "11111111",
	12264 => "11111111",
	12265 => "11111111",
	12266 => "11111111",
	12267 => "11111111",
	12268 => "11111111",
	12269 => "11111111",
	12270 => "11111111",
	12271 => "11111111",
	12272 => "11111111",
	12273 => "11111111",
	12274 => "11111111",
	12275 => "11111111",
	12276 => "11111111",
	12277 => "11111111",
	12278 => "11111111",
	12279 => "11111111",
	12288 => "11111111",
	12289 => "11111111",
	12290 => "11111111",
	12291 => "11111111",
	12292 => "11111111",
	12293 => "11111111",
	12294 => "11111111",
	12295 => "11111111",
	12296 => "11111111",
	12297 => "11111111",
	12298 => "11111111",
	12299 => "11111111",
	12300 => "11111111",
	12301 => "11111111",
	12302 => "11111111",
	12303 => "11111111",
	12304 => "11111111",
	12305 => "11111111",
	12306 => "11111111",
	12307 => "11111111",
	12308 => "11111111",
	12309 => "11111111",
	12310 => "11111111",
	12311 => "11111111",
	12312 => "11111111",
	12313 => "11111111",
	12314 => "11111111",
	12315 => "11111111",
	12316 => "11111111",
	12317 => "11111111",
	12318 => "11111111",
	12319 => "11111111",
	12320 => "11111111",
	12321 => "11111111",
	12322 => "11111111",
	12323 => "11111111",
	12324 => "11111111",
	12325 => "11111111",
	12326 => "11111111",
	12327 => "11111111",
	12328 => "11111111",
	12329 => "11111111",
	12330 => "11111111",
	12331 => "11111111",
	12332 => "11111111",
	12333 => "11111111",
	12334 => "11111111",
	12335 => "11111111",
	12336 => "11111111",
	12337 => "11111111",
	12338 => "11111111",
	12339 => "11111111",
	12340 => "11111111",
	12341 => "11111111",
	12342 => "11111111",
	12343 => "11111111",
	12344 => "11111111",
	12345 => "11111111",
	12346 => "11111111",
	12347 => "11111111",
	12348 => "11111111",
	12349 => "11111111",
	12350 => "11111111",
	12351 => "11111111",
	12352 => "11111111",
	12353 => "11111111",
	12354 => "11111111",
	12355 => "11111111",
	12356 => "11111111",
	12357 => "11111111",
	12358 => "11111111",
	12359 => "11111111",
	12360 => "11111111",
	12361 => "11111111",
	12362 => "11111111",
	12363 => "11111111",
	12364 => "11111111",
	12365 => "11111111",
	12366 => "11111111",
	12367 => "11111111",
	12368 => "11111111",
	12369 => "11111111",
	12370 => "11111111",
	12371 => "11111111",
	12372 => "11111111",
	12373 => "11111111",
	12374 => "11111111",
	12375 => "11111111",
	12376 => "11111111",
	12377 => "11111111",
	12378 => "11111111",
	12379 => "11111111",
	12380 => "11111111",
	12381 => "11111111",
	12382 => "11111111",
	12383 => "11111111",
	12384 => "11111111",
	12385 => "11111111",
	12386 => "11111111",
	12387 => "11111111",
	12388 => "11111111",
	12389 => "11111111",
	12390 => "11111111",
	12391 => "11111111",
	12392 => "11111111",
	12393 => "11111111",
	12394 => "11111111",
	12395 => "11111111",
	12396 => "11111111",
	12397 => "11111111",
	12398 => "11111111",
	12399 => "11111111",
	12400 => "11111111",
	12401 => "11111111",
	12402 => "11111111",
	12403 => "11111111",
	12404 => "11111111",
	12405 => "11111111",
	12406 => "11111111",
	12407 => "11111111",
	12416 => "11111111",
	12417 => "11111111",
	12418 => "11111111",
	12419 => "11111111",
	12420 => "11111111",
	12421 => "11111111",
	12422 => "11111111",
	12423 => "11111111",
	12424 => "11111111",
	12425 => "11111111",
	12426 => "11111111",
	12427 => "11111111",
	12428 => "11111111",
	12429 => "11111111",
	12430 => "11111111",
	12431 => "11111111",
	12432 => "11111111",
	12433 => "11111111",
	12434 => "11111111",
	12435 => "11111111",
	12436 => "11111111",
	12437 => "11111111",
	12438 => "11111111",
	12439 => "11111111",
	12440 => "11111111",
	12441 => "11111111",
	12442 => "11111111",
	12443 => "11111111",
	12444 => "11111111",
	12445 => "11111111",
	12446 => "11111111",
	12447 => "11111111",
	12448 => "11111111",
	12449 => "11111111",
	12450 => "11111111",
	12451 => "11111111",
	12452 => "11111111",
	12453 => "11111111",
	12454 => "11111111",
	12455 => "11111111",
	12456 => "11111111",
	12457 => "11111111",
	12458 => "11111111",
	12459 => "11111111",
	12460 => "11111111",
	12461 => "11111111",
	12462 => "11111111",
	12463 => "11111111",
	12464 => "11111111",
	12465 => "11111111",
	12466 => "11111111",
	12467 => "11111111",
	12468 => "11111111",
	12469 => "11111111",
	12470 => "11111111",
	12471 => "11111111",
	12472 => "11111111",
	12473 => "11111111",
	12474 => "11111111",
	12475 => "11111111",
	12476 => "11111111",
	12477 => "11111111",
	12478 => "11111111",
	12479 => "11111111",
	12480 => "11111111",
	12481 => "11111111",
	12482 => "11111111",
	12483 => "11111111",
	12484 => "11111111",
	12485 => "11111111",
	12486 => "11111111",
	12487 => "11111111",
	12488 => "11111111",
	12489 => "11111111",
	12490 => "11111111",
	12491 => "11111111",
	12492 => "11111111",
	12493 => "11111111",
	12494 => "11111111",
	12495 => "11111111",
	12496 => "11111111",
	12497 => "11111111",
	12498 => "11111111",
	12499 => "11111111",
	12500 => "11111111",
	12501 => "11111111",
	12502 => "11111111",
	12503 => "11111111",
	12504 => "11111111",
	12505 => "11111111",
	12506 => "11111111",
	12507 => "11111111",
	12508 => "11111111",
	12509 => "11111111",
	12510 => "11111111",
	12511 => "11111111",
	12512 => "11111111",
	12513 => "11111111",
	12514 => "11111111",
	12515 => "11111111",
	12516 => "11111111",
	12517 => "11111111",
	12518 => "11111111",
	12519 => "11111111",
	12520 => "11111111",
	12521 => "11111111",
	12522 => "11111111",
	12523 => "11111111",
	12524 => "11111111",
	12525 => "11111111",
	12526 => "11111111",
	12527 => "11111111",
	12528 => "11111111",
	12529 => "11111111",
	12530 => "11111111",
	12531 => "11111111",
	12532 => "11111111",
	12533 => "11111111",
	12534 => "11111111",
	12535 => "11111111",
	12544 => "11111111",
	12545 => "11111111",
	12546 => "11111111",
	12547 => "11111111",
	12548 => "11111111",
	12549 => "11111111",
	12550 => "11111111",
	12551 => "11111111",
	12552 => "11111111",
	12553 => "11111111",
	12554 => "11111111",
	12555 => "11111111",
	12556 => "11111111",
	12557 => "11111111",
	12558 => "11111111",
	12559 => "11111111",
	12560 => "11111111",
	12561 => "11111111",
	12562 => "11111111",
	12563 => "11111111",
	12564 => "11111111",
	12565 => "11111111",
	12566 => "11111111",
	12567 => "11111111",
	12568 => "11111111",
	12569 => "11111111",
	12570 => "11111111",
	12571 => "11111111",
	12572 => "11111111",
	12573 => "11111111",
	12574 => "11111111",
	12575 => "11111111",
	12576 => "11111111",
	12577 => "11111111",
	12578 => "11111111",
	12579 => "11111111",
	12580 => "11111111",
	12581 => "11111111",
	12582 => "11111111",
	12583 => "11111111",
	12584 => "11111111",
	12585 => "11111111",
	12586 => "11111111",
	12587 => "11111111",
	12588 => "11111111",
	12589 => "11111111",
	12590 => "11111111",
	12591 => "11111111",
	12592 => "11111111",
	12593 => "11111111",
	12594 => "11111111",
	12595 => "11111111",
	12596 => "11111111",
	12597 => "11111111",
	12598 => "11111111",
	12599 => "11111111",
	12600 => "11111111",
	12601 => "11111111",
	12602 => "11111111",
	12603 => "11111111",
	12604 => "11111111",
	12605 => "11111111",
	12606 => "11111111",
	12607 => "11111111",
	12608 => "11111111",
	12609 => "11111111",
	12610 => "11111111",
	12611 => "11111111",
	12612 => "11111111",
	12613 => "11111111",
	12614 => "11111111",
	12615 => "11111111",
	12616 => "11111111",
	12617 => "11111111",
	12618 => "11111111",
	12619 => "11111111",
	12620 => "11111111",
	12621 => "11111111",
	12622 => "11111111",
	12623 => "11111111",
	12624 => "11111111",
	12625 => "11111111",
	12626 => "11111111",
	12627 => "11111111",
	12628 => "11111111",
	12629 => "11111111",
	12630 => "11111111",
	12631 => "11111111",
	12632 => "11111111",
	12633 => "11111111",
	12634 => "11111111",
	12635 => "11111111",
	12636 => "11111111",
	12637 => "11111111",
	12638 => "11111111",
	12639 => "11111111",
	12640 => "11111111",
	12641 => "11111111",
	12642 => "11111111",
	12643 => "11111111",
	12644 => "11111111",
	12645 => "11111111",
	12646 => "11111111",
	12647 => "11111111",
	12648 => "11111111",
	12649 => "11111111",
	12650 => "11111111",
	12651 => "11111111",
	12652 => "11111111",
	12653 => "11111111",
	12654 => "11111111",
	12655 => "11111111",
	12656 => "11111111",
	12657 => "11111111",
	12658 => "11111111",
	12659 => "11111111",
	12660 => "11111111",
	12661 => "11111111",
	12662 => "11111111",
	12663 => "11111111",
	12672 => "11111111",
	12673 => "11111111",
	12674 => "11111111",
	12675 => "11111111",
	12676 => "11111111",
	12677 => "11111111",
	12678 => "11111111",
	12679 => "11111111",
	12680 => "11111111",
	12681 => "11111111",
	12682 => "11111111",
	12683 => "11111111",
	12684 => "11111111",
	12685 => "11111111",
	12686 => "11111111",
	12687 => "11111111",
	12688 => "11111111",
	12689 => "11111111",
	12690 => "11111111",
	12691 => "11111111",
	12692 => "11111111",
	12693 => "11111111",
	12694 => "11111111",
	12695 => "11111111",
	12696 => "11111111",
	12697 => "11111111",
	12698 => "11111111",
	12699 => "11111111",
	12700 => "11111111",
	12701 => "11111111",
	12702 => "11111111",
	12703 => "11111111",
	12704 => "11111111",
	12705 => "11111111",
	12706 => "11111111",
	12707 => "11111111",
	12708 => "11111111",
	12709 => "11111111",
	12710 => "11111111",
	12711 => "11111111",
	12712 => "11111111",
	12713 => "11111111",
	12714 => "11111111",
	12715 => "11111111",
	12716 => "11111111",
	12717 => "11111111",
	12718 => "11111111",
	12719 => "11111111",
	12720 => "11111111",
	12721 => "11111111",
	12722 => "11111111",
	12723 => "11111111",
	12724 => "11111111",
	12725 => "11111111",
	12726 => "11111111",
	12727 => "11111111",
	12728 => "11111111",
	12729 => "11111111",
	12730 => "11111111",
	12731 => "11111111",
	12732 => "11111111",
	12733 => "11111111",
	12734 => "11111111",
	12735 => "11111111",
	12736 => "11111111",
	12737 => "11111111",
	12738 => "11111111",
	12739 => "11111111",
	12740 => "11111111",
	12741 => "11111111",
	12742 => "11111111",
	12743 => "11111111",
	12744 => "11111111",
	12745 => "11111111",
	12746 => "11111111",
	12747 => "11111111",
	12748 => "11111111",
	12749 => "11111111",
	12750 => "11111111",
	12751 => "11111111",
	12752 => "11111111",
	12753 => "11111111",
	12754 => "11111111",
	12755 => "11111111",
	12756 => "11111111",
	12757 => "11111111",
	12758 => "11111111",
	12759 => "11111111",
	12760 => "11111111",
	12761 => "11111111",
	12762 => "11111111",
	12763 => "11111111",
	12764 => "11111111",
	12765 => "11111111",
	12766 => "11111111",
	12767 => "11111111",
	12768 => "11111111",
	12769 => "11111111",
	12770 => "11111111",
	12771 => "11111111",
	12772 => "11111111",
	12773 => "11111111",
	12774 => "11111111",
	12775 => "11111111",
	12776 => "11111111",
	12777 => "11111111",
	12778 => "11111111",
	12779 => "11111111",
	12780 => "11111111",
	12781 => "11111111",
	12782 => "11111111",
	12783 => "11111111",
	12784 => "11111111",
	12785 => "11111111",
	12786 => "11111111",
	12787 => "11111111",
	12788 => "11111111",
	12789 => "11111111",
	12790 => "11111111",
	12791 => "11111111",
	12800 => "11111111",
	12801 => "11111111",
	12802 => "11111111",
	12803 => "11111111",
	12804 => "11111111",
	12805 => "11111111",
	12806 => "11111111",
	12807 => "11111111",
	12808 => "11111111",
	12809 => "11111111",
	12810 => "11111111",
	12811 => "11111111",
	12812 => "11111111",
	12813 => "11111111",
	12814 => "11111111",
	12815 => "11111111",
	12816 => "11111111",
	12817 => "11111111",
	12818 => "11111111",
	12819 => "11111111",
	12820 => "11111111",
	12821 => "11111111",
	12822 => "11111111",
	12823 => "11111111",
	12824 => "11111111",
	12825 => "11111111",
	12826 => "11111111",
	12827 => "11111111",
	12828 => "11111111",
	12829 => "11111111",
	12830 => "11111111",
	12831 => "11111111",
	12832 => "11111111",
	12833 => "11111111",
	12834 => "11111111",
	12835 => "11111111",
	12836 => "11111111",
	12837 => "11111111",
	12838 => "11111111",
	12839 => "11111111",
	12840 => "11111111",
	12841 => "11111111",
	12842 => "11111111",
	12843 => "11111111",
	12844 => "11111111",
	12845 => "11111111",
	12846 => "11111111",
	12847 => "11111111",
	12848 => "11111111",
	12849 => "11111111",
	12850 => "11111111",
	12851 => "11111111",
	12852 => "11111111",
	12853 => "11111111",
	12854 => "11111111",
	12855 => "11111111",
	12856 => "11111111",
	12857 => "11111111",
	12858 => "11111111",
	12859 => "11111111",
	12860 => "11111111",
	12861 => "11111111",
	12862 => "11111111",
	12863 => "11111111",
	12864 => "11111111",
	12865 => "11111111",
	12866 => "11111111",
	12867 => "11111111",
	12868 => "11111111",
	12869 => "11111111",
	12870 => "11111111",
	12871 => "11111111",
	12872 => "11111111",
	12873 => "11111111",
	12874 => "11111111",
	12875 => "11111111",
	12876 => "11111111",
	12877 => "11111111",
	12878 => "11111111",
	12879 => "11111111",
	12880 => "11111111",
	12881 => "11111111",
	12882 => "11111111",
	12883 => "11111111",
	12884 => "11111111",
	12885 => "11111111",
	12886 => "11111111",
	12887 => "11111111",
	12888 => "11111111",
	12889 => "11111111",
	12890 => "11111111",
	12891 => "11111111",
	12892 => "11111111",
	12893 => "11111111",
	12894 => "11111111",
	12895 => "11111111",
	12896 => "11111111",
	12897 => "11111111",
	12898 => "11111111",
	12899 => "11111111",
	12900 => "11111111",
	12901 => "11111111",
	12902 => "11111111",
	12903 => "11111111",
	12904 => "11111111",
	12905 => "11111111",
	12906 => "11111111",
	12907 => "11111111",
	12908 => "11111111",
	12909 => "11111111",
	12910 => "11111111",
	12911 => "11111111",
	12912 => "11111111",
	12913 => "11111111",
	12914 => "11111111",
	12915 => "11111111",
	12916 => "11111111",
	12917 => "11111111",
	12918 => "11111111",
	12919 => "11111111",
	12928 => "11111111",
	12929 => "11111111",
	12930 => "11111111",
	12931 => "11111111",
	12932 => "11111111",
	12933 => "11111111",
	12934 => "11111111",
	12935 => "11111111",
	12936 => "11111111",
	12937 => "11111111",
	12938 => "11111111",
	12939 => "11111111",
	12940 => "11111111",
	12941 => "11111111",
	12942 => "11111111",
	12943 => "11111111",
	12944 => "11111111",
	12945 => "11111111",
	12946 => "11111111",
	12947 => "11111111",
	12948 => "11111111",
	12949 => "11111111",
	12950 => "11111111",
	12951 => "11111111",
	12952 => "11111111",
	12953 => "11111111",
	12954 => "11111111",
	12955 => "11111111",
	12956 => "11111111",
	12957 => "11111111",
	12958 => "11111111",
	12959 => "11111111",
	12960 => "11111111",
	12961 => "11111111",
	12962 => "11111111",
	12963 => "11111111",
	12964 => "11111111",
	12965 => "11111111",
	12966 => "11111111",
	12967 => "11111111",
	12968 => "11111111",
	12969 => "11111111",
	12970 => "11111111",
	12971 => "11111111",
	12972 => "11111111",
	12973 => "11111111",
	12974 => "11111111",
	12975 => "11111111",
	12976 => "11111111",
	12977 => "11111111",
	12978 => "11111111",
	12979 => "11111111",
	12980 => "11111111",
	12981 => "11111111",
	12982 => "11111111",
	12983 => "11111111",
	12984 => "11111111",
	12985 => "11111111",
	12986 => "11111111",
	12987 => "11111111",
	12988 => "11111111",
	12989 => "11111111",
	12990 => "11111111",
	12991 => "11111111",
	12992 => "11111111",
	12993 => "11111111",
	12994 => "11111111",
	12995 => "11111111",
	12996 => "11111111",
	12997 => "11111111",
	12998 => "11111111",
	12999 => "11111111",
	13000 => "11111111",
	13001 => "11111111",
	13002 => "11111111",
	13003 => "11111111",
	13004 => "11111111",
	13005 => "11111111",
	13006 => "11111111",
	13007 => "11111111",
	13008 => "11111111",
	13009 => "11111111",
	13010 => "11111111",
	13011 => "11111111",
	13012 => "11111111",
	13013 => "11111111",
	13014 => "11111111",
	13015 => "11111111",
	13016 => "11111111",
	13017 => "11111111",
	13018 => "11111111",
	13019 => "11111111",
	13020 => "11111111",
	13021 => "11111111",
	13022 => "11111111",
	13023 => "11111111",
	13024 => "11111111",
	13025 => "11111111",
	13026 => "11111111",
	13027 => "11111111",
	13028 => "11111111",
	13029 => "11111111",
	13030 => "11111111",
	13031 => "11111111",
	13032 => "11111111",
	13033 => "11111111",
	13034 => "11111111",
	13035 => "11111111",
	13036 => "11111111",
	13037 => "11111111",
	13038 => "11111111",
	13039 => "11111111",
	13040 => "11111111",
	13041 => "11111111",
	13042 => "11111111",
	13043 => "11111111",
	13044 => "11111111",
	13045 => "11111111",
	13046 => "11111111",
	13047 => "11111111",
	13056 => "11111111",
	13057 => "11111111",
	13058 => "11111111",
	13059 => "11111111",
	13060 => "11111111",
	13061 => "11111111",
	13062 => "11111111",
	13063 => "11111111",
	13064 => "11111111",
	13065 => "11111111",
	13066 => "11111111",
	13067 => "11111111",
	13068 => "11111111",
	13069 => "11111111",
	13070 => "11111111",
	13071 => "11111111",
	13072 => "11111111",
	13073 => "11111111",
	13074 => "11111111",
	13075 => "11111111",
	13076 => "11111111",
	13077 => "11111111",
	13078 => "11111111",
	13079 => "11111111",
	13080 => "11111111",
	13081 => "11111111",
	13082 => "11111111",
	13083 => "11111111",
	13084 => "11111111",
	13085 => "11111111",
	13086 => "11111111",
	13087 => "11111111",
	13088 => "11111111",
	13089 => "11111111",
	13090 => "11111111",
	13091 => "11111111",
	13092 => "11111111",
	13093 => "11111111",
	13094 => "11111111",
	13095 => "11111111",
	13096 => "11111111",
	13097 => "11111111",
	13098 => "11111111",
	13099 => "11111111",
	13100 => "11111111",
	13101 => "11111111",
	13102 => "11111111",
	13103 => "11111111",
	13104 => "11111111",
	13105 => "11111111",
	13106 => "11111111",
	13107 => "11111111",
	13108 => "11111111",
	13109 => "11111111",
	13110 => "11111111",
	13111 => "11111111",
	13112 => "11111111",
	13113 => "11111111",
	13114 => "11111111",
	13115 => "11111111",
	13116 => "11111111",
	13117 => "11111111",
	13118 => "11111111",
	13119 => "11111111",
	13120 => "11111111",
	13121 => "11111111",
	13122 => "11111111",
	13123 => "11111111",
	13124 => "11111111",
	13125 => "11111111",
	13126 => "11111111",
	13127 => "11111111",
	13128 => "11111111",
	13129 => "11111111",
	13130 => "11111111",
	13131 => "11111111",
	13132 => "11111111",
	13133 => "11111111",
	13134 => "11111111",
	13135 => "11111111",
	13136 => "11111111",
	13137 => "11111111",
	13138 => "11111111",
	13139 => "11111111",
	13140 => "11111111",
	13141 => "11111111",
	13142 => "11111111",
	13143 => "11111111",
	13144 => "11111111",
	13145 => "11111111",
	13146 => "11111111",
	13147 => "11111111",
	13148 => "11111111",
	13149 => "11111111",
	13150 => "11111111",
	13151 => "11111111",
	13152 => "11111111",
	13153 => "11111111",
	13154 => "11111111",
	13155 => "11111111",
	13156 => "11111111",
	13157 => "11111111",
	13158 => "11111111",
	13159 => "11111111",
	13160 => "11111111",
	13161 => "11111111",
	13162 => "11111111",
	13163 => "11111111",
	13164 => "11111111",
	13165 => "11111111",
	13166 => "11111111",
	13167 => "11111111",
	13168 => "11111111",
	13169 => "11111111",
	13170 => "11111111",
	13171 => "11111111",
	13172 => "11111111",
	13173 => "11111111",
	13174 => "11111111",
	13175 => "11111111",
	13184 => "11111111",
	13185 => "11111111",
	13186 => "11111111",
	13187 => "11111111",
	13188 => "11111111",
	13189 => "11111111",
	13190 => "11111111",
	13191 => "11111111",
	13192 => "11111111",
	13193 => "11111111",
	13194 => "11111111",
	13195 => "11111111",
	13196 => "11111111",
	13197 => "11111111",
	13198 => "11111111",
	13199 => "11111111",
	13200 => "11111111",
	13201 => "11111111",
	13202 => "11111111",
	13203 => "11111111",
	13204 => "11111111",
	13205 => "11111111",
	13206 => "11111111",
	13207 => "11111111",
	13208 => "11111111",
	13209 => "11111111",
	13210 => "11111111",
	13211 => "11111111",
	13212 => "11111111",
	13213 => "11111111",
	13214 => "11111111",
	13215 => "11111111",
	13216 => "11111111",
	13217 => "11111111",
	13218 => "11111111",
	13219 => "11111111",
	13220 => "11111111",
	13221 => "11111111",
	13222 => "11111111",
	13223 => "11111111",
	13224 => "11111111",
	13225 => "11111111",
	13226 => "11111111",
	13227 => "11111111",
	13228 => "11111111",
	13229 => "11111111",
	13230 => "11111111",
	13231 => "11111111",
	13232 => "11111111",
	13233 => "11111111",
	13234 => "11111111",
	13235 => "11111111",
	13236 => "11111111",
	13237 => "11111111",
	13238 => "11111111",
	13239 => "11111111",
	13240 => "11111111",
	13241 => "11111111",
	13242 => "11111111",
	13243 => "11111111",
	13244 => "11111111",
	13245 => "11111111",
	13246 => "11111111",
	13247 => "11111111",
	13248 => "11111111",
	13249 => "11111111",
	13250 => "11111111",
	13251 => "11111111",
	13252 => "11111111",
	13253 => "11111111",
	13254 => "11111111",
	13255 => "11111111",
	13256 => "11111111",
	13257 => "11111111",
	13258 => "11111111",
	13259 => "11111111",
	13260 => "11111111",
	13261 => "11111111",
	13262 => "11111111",
	13263 => "11111111",
	13264 => "11111111",
	13265 => "11111111",
	13266 => "11111111",
	13267 => "11111111",
	13268 => "11111111",
	13269 => "11111111",
	13270 => "11111111",
	13271 => "11111111",
	13272 => "11111111",
	13273 => "11111111",
	13274 => "11111111",
	13275 => "11111111",
	13276 => "11111111",
	13277 => "11111111",
	13278 => "11111111",
	13279 => "11111111",
	13280 => "11111111",
	13281 => "11111111",
	13282 => "11111111",
	13283 => "11111111",
	13284 => "11111111",
	13285 => "11111111",
	13286 => "11111111",
	13287 => "11111111",
	13288 => "11111111",
	13289 => "11111111",
	13290 => "11111111",
	13291 => "11111111",
	13292 => "11111111",
	13293 => "11111111",
	13294 => "11111111",
	13295 => "11111111",
	13296 => "11111111",
	13297 => "11111111",
	13298 => "11111111",
	13299 => "11111111",
	13300 => "11111111",
	13301 => "11111111",
	13302 => "11111111",
	13303 => "11111111",
	13312 => "11111111",
	13313 => "11111111",
	13314 => "11111111",
	13315 => "11111111",
	13316 => "11111111",
	13317 => "11111111",
	13318 => "11111111",
	13319 => "11111111",
	13320 => "11111111",
	13321 => "11111111",
	13322 => "11111111",
	13323 => "11111111",
	13324 => "11111111",
	13325 => "11111111",
	13326 => "11111111",
	13327 => "11111111",
	13328 => "11111111",
	13329 => "11111111",
	13330 => "11111111",
	13331 => "11111111",
	13332 => "11111111",
	13333 => "11111111",
	13334 => "11111111",
	13335 => "11111111",
	13336 => "11111111",
	13337 => "11111111",
	13338 => "11111111",
	13339 => "11111111",
	13340 => "11111111",
	13341 => "11111111",
	13342 => "11111111",
	13343 => "11111111",
	13344 => "11111111",
	13345 => "11111111",
	13346 => "11111111",
	13347 => "11111111",
	13348 => "11111111",
	13349 => "11111111",
	13350 => "11111111",
	13351 => "11111111",
	13352 => "11111111",
	13353 => "11111111",
	13354 => "11111111",
	13355 => "11111111",
	13356 => "11111111",
	13357 => "11111111",
	13358 => "11111111",
	13359 => "11111111",
	13360 => "11111111",
	13361 => "11111111",
	13362 => "11111111",
	13363 => "11111111",
	13364 => "11111111",
	13365 => "11111111",
	13366 => "11111111",
	13367 => "11111111",
	13368 => "11111111",
	13369 => "11111111",
	13370 => "11111111",
	13371 => "11111111",
	13372 => "11111111",
	13373 => "11111111",
	13374 => "11111111",
	13375 => "11111111",
	13376 => "11111111",
	13377 => "11111111",
	13378 => "11111111",
	13379 => "11111111",
	13380 => "11111111",
	13381 => "11111111",
	13382 => "11111111",
	13383 => "11111111",
	13384 => "11111111",
	13385 => "11111111",
	13386 => "11111111",
	13387 => "11111111",
	13388 => "11111111",
	13389 => "11111111",
	13390 => "11111111",
	13391 => "11111111",
	13392 => "11111111",
	13393 => "11111111",
	13394 => "11111111",
	13395 => "11111111",
	13396 => "11111111",
	13397 => "11111111",
	13398 => "11111111",
	13399 => "11111111",
	13400 => "11111111",
	13401 => "11111111",
	13402 => "11111111",
	13403 => "11111111",
	13404 => "11111111",
	13405 => "11111111",
	13406 => "11111111",
	13407 => "11111111",
	13408 => "11111111",
	13409 => "11111111",
	13410 => "11111111",
	13411 => "11111111",
	13412 => "11111111",
	13413 => "11111111",
	13414 => "11111111",
	13415 => "11111111",
	13416 => "11111111",
	13417 => "11111111",
	13418 => "11111111",
	13419 => "11111111",
	13420 => "11111111",
	13421 => "11111111",
	13422 => "11111111",
	13423 => "11111111",
	13424 => "11111111",
	13425 => "11111111",
	13426 => "11111111",
	13427 => "11111111",
	13428 => "11111111",
	13429 => "11111111",
	13430 => "11111111",
	13431 => "11111111",
	13440 => "11111111",
	13441 => "11111111",
	13442 => "11111111",
	13443 => "11111111",
	13444 => "11111111",
	13445 => "11111111",
	13446 => "11111111",
	13447 => "11111111",
	13448 => "11111111",
	13449 => "11111111",
	13450 => "11111111",
	13451 => "11111111",
	13452 => "11111111",
	13453 => "11111111",
	13454 => "11111111",
	13455 => "11111111",
	13456 => "11111111",
	13457 => "11111111",
	13458 => "11111111",
	13459 => "11111111",
	13460 => "11111111",
	13461 => "11111111",
	13462 => "11111111",
	13463 => "11111111",
	13464 => "11111111",
	13465 => "11111111",
	13466 => "11111111",
	13467 => "11111111",
	13468 => "11111111",
	13469 => "11111111",
	13470 => "11111111",
	13471 => "11111111",
	13472 => "11111111",
	13473 => "11111111",
	13474 => "11111111",
	13475 => "11111111",
	13476 => "11111111",
	13477 => "11111111",
	13478 => "11111111",
	13479 => "11111111",
	13480 => "11111111",
	13481 => "11111111",
	13482 => "11111111",
	13483 => "11111111",
	13484 => "11111111",
	13485 => "11111111",
	13486 => "11111111",
	13487 => "11111111",
	13488 => "11111111",
	13489 => "11111111",
	13490 => "11111111",
	13491 => "11111111",
	13492 => "11111111",
	13493 => "11111111",
	13494 => "11111111",
	13495 => "11111111",
	13496 => "11111111",
	13497 => "11111111",
	13498 => "11111111",
	13499 => "11111111",
	13500 => "11111111",
	13501 => "11111111",
	13502 => "11111111",
	13503 => "11111111",
	13504 => "11111111",
	13505 => "11111111",
	13506 => "11111111",
	13507 => "11111111",
	13508 => "11111111",
	13509 => "11111111",
	13510 => "11111111",
	13511 => "11111111",
	13512 => "11111111",
	13513 => "11111111",
	13514 => "11111111",
	13515 => "11111111",
	13516 => "11111111",
	13517 => "11111111",
	13518 => "11111111",
	13519 => "11111111",
	13520 => "11111111",
	13521 => "11111111",
	13522 => "11111111",
	13523 => "11111111",
	13524 => "11111111",
	13525 => "11111111",
	13526 => "11111111",
	13527 => "11111111",
	13528 => "11111111",
	13529 => "11111111",
	13530 => "11111111",
	13531 => "11111111",
	13532 => "11111111",
	13533 => "11111111",
	13534 => "11111111",
	13535 => "11111111",
	13536 => "11111111",
	13537 => "11111111",
	13538 => "11111111",
	13539 => "11111111",
	13540 => "11111111",
	13541 => "11111111",
	13542 => "11111111",
	13543 => "11111111",
	13544 => "11111111",
	13545 => "11111111",
	13546 => "11111111",
	13547 => "11111111",
	13548 => "11111111",
	13549 => "11111111",
	13550 => "11111111",
	13551 => "11111111",
	13552 => "11111111",
	13553 => "11111111",
	13554 => "11111111",
	13555 => "11111111",
	13556 => "11111111",
	13557 => "11111111",
	13558 => "11111111",
	13559 => "11111111",
	13568 => "11111111",
	13569 => "11111111",
	13570 => "11111111",
	13571 => "11111111",
	13572 => "11111111",
	13573 => "11111111",
	13574 => "11111111",
	13575 => "11111111",
	13576 => "11111111",
	13577 => "11111111",
	13578 => "11111111",
	13579 => "11111111",
	13580 => "11111111",
	13581 => "11111111",
	13582 => "11111111",
	13583 => "11111111",
	13584 => "11111111",
	13585 => "11111111",
	13586 => "11111111",
	13587 => "11111111",
	13588 => "11111111",
	13589 => "11111111",
	13590 => "11111111",
	13591 => "11111111",
	13592 => "11111111",
	13593 => "11111111",
	13594 => "11111111",
	13595 => "11111111",
	13596 => "11111111",
	13597 => "11111111",
	13598 => "11111111",
	13599 => "11111111",
	13600 => "11111111",
	13601 => "11111111",
	13602 => "11111111",
	13603 => "11111111",
	13604 => "11111111",
	13605 => "11111111",
	13606 => "11111111",
	13607 => "11111111",
	13608 => "11111111",
	13609 => "11111111",
	13610 => "11111111",
	13611 => "11111111",
	13612 => "11111111",
	13613 => "11111111",
	13614 => "11111111",
	13615 => "11111111",
	13616 => "11111111",
	13617 => "11111111",
	13618 => "11111111",
	13619 => "11111111",
	13620 => "11111111",
	13621 => "11111111",
	13622 => "11111111",
	13623 => "11111111",
	13624 => "11111111",
	13625 => "11111111",
	13626 => "11111111",
	13627 => "11111111",
	13628 => "11111111",
	13629 => "11111111",
	13630 => "11111111",
	13631 => "11111111",
	13632 => "11111111",
	13633 => "11111111",
	13634 => "11111111",
	13635 => "11111111",
	13636 => "11111111",
	13637 => "11111111",
	13638 => "11111111",
	13639 => "11111111",
	13640 => "11111111",
	13641 => "11111111",
	13642 => "11111111",
	13643 => "11111111",
	13644 => "11111111",
	13645 => "11111111",
	13646 => "11111111",
	13647 => "11111111",
	13648 => "11111111",
	13649 => "11111111",
	13650 => "11111111",
	13651 => "11111111",
	13652 => "11111111",
	13653 => "11111111",
	13654 => "11111111",
	13655 => "11111111",
	13656 => "11111111",
	13657 => "11111111",
	13658 => "11111111",
	13659 => "11111111",
	13660 => "11111111",
	13661 => "11111111",
	13662 => "11111111",
	13663 => "11111111",
	13664 => "11111111",
	13665 => "11111111",
	13666 => "11111111",
	13667 => "11111111",
	13668 => "11111111",
	13669 => "11111111",
	13670 => "11111111",
	13671 => "11111111",
	13672 => "11111111",
	13673 => "11111111",
	13674 => "11111111",
	13675 => "11111111",
	13676 => "11111111",
	13677 => "11111111",
	13678 => "11111111",
	13679 => "11111111",
	13680 => "11111111",
	13681 => "11111111",
	13682 => "11111111",
	13683 => "11111111",
	13684 => "11111111",
	13685 => "11111111",
	13686 => "11111111",
	13687 => "11111111",
	13696 => "11111111",
	13697 => "11111111",
	13698 => "11111111",
	13699 => "11111111",
	13700 => "11111111",
	13701 => "11111111",
	13702 => "11111111",
	13703 => "11111111",
	13704 => "11111111",
	13705 => "11111111",
	13706 => "11111111",
	13707 => "11111111",
	13708 => "11111111",
	13709 => "11111111",
	13710 => "11111111",
	13711 => "11111111",
	13712 => "11111111",
	13713 => "11111111",
	13714 => "11111111",
	13715 => "11111111",
	13716 => "11111111",
	13717 => "11111111",
	13718 => "11111111",
	13719 => "11111111",
	13720 => "11111111",
	13721 => "11111111",
	13722 => "11111111",
	13723 => "11111111",
	13724 => "11111111",
	13725 => "11111111",
	13726 => "11111111",
	13727 => "11111111",
	13728 => "11111111",
	13729 => "11111111",
	13730 => "11111111",
	13731 => "11111111",
	13732 => "11111111",
	13733 => "11111111",
	13734 => "11111111",
	13735 => "11111111",
	13736 => "11111111",
	13737 => "11111111",
	13738 => "11111111",
	13739 => "11111111",
	13740 => "11111111",
	13741 => "11111111",
	13742 => "11111111",
	13743 => "11111111",
	13744 => "11111111",
	13745 => "11111111",
	13746 => "11111111",
	13747 => "11111111",
	13748 => "11111111",
	13749 => "11111111",
	13750 => "11111111",
	13751 => "11111111",
	13752 => "11111111",
	13753 => "11111111",
	13754 => "11111111",
	13755 => "11111111",
	13756 => "11111111",
	13757 => "11111111",
	13758 => "11111111",
	13759 => "11111111",
	13760 => "11111111",
	13761 => "11111111",
	13762 => "11111111",
	13763 => "11111111",
	13764 => "11111111",
	13765 => "11111111",
	13766 => "11111111",
	13767 => "11111111",
	13768 => "11111111",
	13769 => "11111111",
	13770 => "11111111",
	13771 => "11111111",
	13772 => "11111111",
	13773 => "11111111",
	13774 => "11111111",
	13775 => "11111111",
	13776 => "11111111",
	13777 => "11111111",
	13778 => "11111111",
	13779 => "11111111",
	13780 => "11111111",
	13781 => "11111111",
	13782 => "11111111",
	13783 => "11111111",
	13784 => "11111111",
	13785 => "11111111",
	13786 => "11111111",
	13787 => "11111111",
	13788 => "11111111",
	13789 => "11111111",
	13790 => "11111111",
	13791 => "11111111",
	13792 => "11111111",
	13793 => "11111111",
	13794 => "11111111",
	13795 => "11111111",
	13796 => "11111111",
	13797 => "11111111",
	13798 => "11111111",
	13799 => "11111111",
	13800 => "11111111",
	13801 => "11111111",
	13802 => "11111111",
	13803 => "11111111",
	13804 => "11111111",
	13805 => "11111111",
	13806 => "11111111",
	13807 => "11111111",
	13808 => "11111111",
	13809 => "11111111",
	13810 => "11111111",
	13811 => "11111111",
	13812 => "11111111",
	13813 => "11111111",
	13814 => "11111111",
	13815 => "11111111",
	13824 => "11111111",
	13825 => "11111111",
	13826 => "11111111",
	13827 => "11111111",
	13828 => "11111111",
	13829 => "11111111",
	13830 => "11111111",
	13831 => "11111111",
	13832 => "11111111",
	13833 => "11111111",
	13834 => "11111111",
	13835 => "11111111",
	13836 => "11111111",
	13837 => "11111111",
	13838 => "11111111",
	13839 => "11111111",
	13840 => "11111111",
	13841 => "11111111",
	13842 => "11111111",
	13843 => "11111111",
	13844 => "11111111",
	13845 => "11111111",
	13846 => "11111111",
	13847 => "11111111",
	13848 => "11111111",
	13849 => "11111111",
	13850 => "11111111",
	13851 => "11111111",
	13852 => "11111111",
	13853 => "11111111",
	13854 => "11111111",
	13855 => "11111111",
	13856 => "11111111",
	13857 => "11111111",
	13858 => "11111111",
	13859 => "11111111",
	13860 => "11111111",
	13861 => "11111111",
	13862 => "11111111",
	13863 => "11111111",
	13864 => "11111111",
	13865 => "11111111",
	13866 => "11111111",
	13867 => "11111111",
	13868 => "11111111",
	13869 => "11111111",
	13870 => "11111111",
	13871 => "11111111",
	13872 => "11111111",
	13873 => "11111111",
	13874 => "11111111",
	13875 => "11111111",
	13876 => "11111111",
	13877 => "11111111",
	13878 => "11111111",
	13879 => "11111111",
	13880 => "11111111",
	13881 => "11111111",
	13882 => "11111111",
	13883 => "11111111",
	13884 => "11111111",
	13885 => "11111111",
	13886 => "11111111",
	13887 => "11111111",
	13888 => "11111111",
	13889 => "11111111",
	13890 => "11111111",
	13891 => "11111111",
	13892 => "11111111",
	13893 => "11111111",
	13894 => "11111111",
	13895 => "11111111",
	13896 => "11111111",
	13897 => "11111111",
	13898 => "11111111",
	13899 => "11111111",
	13900 => "11111111",
	13901 => "11111111",
	13902 => "11111111",
	13903 => "11111111",
	13904 => "11111111",
	13905 => "11111111",
	13906 => "11111111",
	13907 => "11111111",
	13908 => "11111111",
	13909 => "11111111",
	13910 => "11111111",
	13911 => "11111111",
	13912 => "11111111",
	13913 => "11111111",
	13914 => "11111111",
	13915 => "11111111",
	13916 => "11111111",
	13917 => "11111111",
	13918 => "11111111",
	13919 => "11111111",
	13920 => "11111111",
	13921 => "11111111",
	13922 => "11111111",
	13923 => "11111111",
	13924 => "11111111",
	13925 => "11111111",
	13926 => "11111111",
	13927 => "11111111",
	13928 => "11111111",
	13929 => "11111111",
	13930 => "11111111",
	13931 => "11111111",
	13932 => "11111111",
	13933 => "11111111",
	13934 => "11111111",
	13935 => "11111111",
	13936 => "11111111",
	13937 => "11111111",
	13938 => "11111111",
	13939 => "11111111",
	13940 => "11111111",
	13941 => "11111111",
	13942 => "11111111",
	13943 => "11111111",
	13952 => "11111111",
	13953 => "11111111",
	13954 => "11111111",
	13955 => "11111111",
	13956 => "11111111",
	13957 => "11111111",
	13958 => "11111111",
	13959 => "11111111",
	13960 => "11111111",
	13961 => "11111111",
	13962 => "11111111",
	13963 => "11111111",
	13964 => "11111111",
	13965 => "11111111",
	13966 => "11111111",
	13967 => "11111111",
	13968 => "11111111",
	13969 => "11111111",
	13970 => "11111111",
	13971 => "11111111",
	13972 => "11111111",
	13973 => "11111111",
	13974 => "11111111",
	13975 => "11111111",
	13976 => "11111111",
	13977 => "11111111",
	13978 => "11111111",
	13979 => "11111111",
	13980 => "11111111",
	13981 => "11111111",
	13982 => "11111111",
	13983 => "11111111",
	13984 => "11111111",
	13985 => "11111111",
	13986 => "11111111",
	13987 => "11111111",
	13988 => "11111111",
	13989 => "11111111",
	13990 => "11111111",
	13991 => "11111111",
	13992 => "11111111",
	13993 => "11111111",
	13994 => "11111111",
	13995 => "11111111",
	13996 => "11111111",
	13997 => "11111111",
	13998 => "11111111",
	13999 => "11111111",
	14000 => "11111111",
	14001 => "11111111",
	14002 => "11111111",
	14003 => "11111111",
	14004 => "11111111",
	14005 => "11111111",
	14006 => "11111111",
	14007 => "11111111",
	14008 => "11111111",
	14009 => "11111111",
	14010 => "11111111",
	14011 => "11111111",
	14012 => "11111111",
	14013 => "11111111",
	14014 => "11111111",
	14015 => "11111111",
	14016 => "11111111",
	14017 => "11111111",
	14018 => "11111111",
	14019 => "11111111",
	14020 => "11111111",
	14021 => "11111111",
	14022 => "11111111",
	14023 => "11111111",
	14024 => "11111111",
	14025 => "11111111",
	14026 => "11111111",
	14027 => "11111111",
	14028 => "11111111",
	14029 => "11111111",
	14030 => "11111111",
	14031 => "11111111",
	14032 => "11111111",
	14033 => "11111111",
	14034 => "11111111",
	14035 => "11111111",
	14036 => "11111111",
	14037 => "11111111",
	14038 => "11111111",
	14039 => "11111111",
	14040 => "11111111",
	14041 => "11111111",
	14042 => "11111111",
	14043 => "11111111",
	14044 => "11111111",
	14045 => "11111111",
	14046 => "11111111",
	14047 => "11111111",
	14048 => "11111111",
	14049 => "11111111",
	14050 => "11111111",
	14051 => "11111111",
	14052 => "11111111",
	14053 => "11111111",
	14054 => "11111111",
	14055 => "11111111",
	14056 => "11111111",
	14057 => "11111111",
	14058 => "11111111",
	14059 => "11111111",
	14060 => "11111111",
	14061 => "11111111",
	14062 => "11111111",
	14063 => "11111111",
	14064 => "11111111",
	14065 => "11111111",
	14066 => "11111111",
	14067 => "11111111",
	14068 => "11111111",
	14069 => "11111111",
	14070 => "11111111",
	14071 => "11111111",
	14080 => "11111111",
	14081 => "11111111",
	14082 => "11111111",
	14083 => "11111111",
	14084 => "11111111",
	14085 => "11111111",
	14086 => "11111111",
	14087 => "11111111",
	14088 => "11111111",
	14089 => "11111111",
	14090 => "11111111",
	14091 => "11111111",
	14092 => "11111111",
	14093 => "11111111",
	14094 => "11111111",
	14095 => "11111111",
	14096 => "11111111",
	14097 => "11111111",
	14098 => "11111111",
	14099 => "11111111",
	14100 => "11111111",
	14101 => "11111111",
	14102 => "11111111",
	14103 => "11111111",
	14104 => "11111111",
	14105 => "11111111",
	14106 => "11111111",
	14107 => "11111111",
	14108 => "11111111",
	14109 => "11111111",
	14110 => "11111111",
	14111 => "11111111",
	14112 => "11111111",
	14113 => "11111111",
	14114 => "11111111",
	14115 => "11111111",
	14116 => "11111111",
	14117 => "11111111",
	14118 => "11111111",
	14119 => "11111111",
	14120 => "11111111",
	14121 => "11111111",
	14122 => "11111111",
	14123 => "11111111",
	14124 => "11111111",
	14125 => "11111111",
	14126 => "11111111",
	14127 => "11111111",
	14128 => "11111111",
	14129 => "11111111",
	14130 => "11111111",
	14131 => "11111111",
	14132 => "11111111",
	14133 => "11111111",
	14134 => "11111111",
	14135 => "11111111",
	14136 => "11111111",
	14137 => "11111111",
	14138 => "11111111",
	14139 => "11111111",
	14140 => "11111111",
	14141 => "11111111",
	14142 => "11111111",
	14143 => "11111111",
	14144 => "11111111",
	14145 => "11111111",
	14146 => "11111111",
	14147 => "11111111",
	14148 => "11111111",
	14149 => "11111111",
	14150 => "11111111",
	14151 => "11111111",
	14152 => "11111111",
	14153 => "11111111",
	14154 => "11111111",
	14155 => "11111111",
	14156 => "11111111",
	14157 => "11111111",
	14158 => "11111111",
	14159 => "11111111",
	14160 => "11111111",
	14161 => "11111111",
	14162 => "11111111",
	14163 => "11111111",
	14164 => "11111111",
	14165 => "11111111",
	14166 => "11111111",
	14167 => "11111111",
	14168 => "11111111",
	14169 => "11111111",
	14170 => "11111111",
	14171 => "11111111",
	14172 => "11111111",
	14173 => "11111111",
	14174 => "11111111",
	14175 => "11111111",
	14176 => "11111111",
	14177 => "11111111",
	14178 => "11111111",
	14179 => "11111111",
	14180 => "11111111",
	14181 => "11111111",
	14182 => "11111111",
	14183 => "11111111",
	14184 => "11111111",
	14185 => "11111111",
	14186 => "11111111",
	14187 => "11111111",
	14188 => "11111111",
	14189 => "11111111",
	14190 => "11111111",
	14191 => "11111111",
	14192 => "11111111",
	14193 => "11111111",
	14194 => "11111111",
	14195 => "11111111",
	14196 => "11111111",
	14197 => "11111111",
	14198 => "11111111",
	14199 => "11111111",
	14208 => "11111111",
	14209 => "11111111",
	14210 => "11111111",
	14211 => "11111111",
	14212 => "11111111",
	14213 => "11111111",
	14214 => "11111111",
	14215 => "11111111",
	14216 => "11111111",
	14217 => "11111111",
	14218 => "11111111",
	14219 => "11111111",
	14220 => "11111111",
	14221 => "11111111",
	14222 => "11111111",
	14223 => "11111111",
	14224 => "11111111",
	14225 => "11111111",
	14226 => "11111111",
	14227 => "11111111",
	14228 => "11111111",
	14229 => "11111111",
	14230 => "11111111",
	14231 => "11111111",
	14232 => "11111111",
	14233 => "11111111",
	14234 => "11111111",
	14235 => "11111111",
	14236 => "11111111",
	14237 => "11111111",
	14238 => "11111111",
	14239 => "11111111",
	14240 => "11111111",
	14241 => "11111111",
	14242 => "11111111",
	14243 => "11111111",
	14244 => "11111111",
	14245 => "11111111",
	14246 => "11111111",
	14247 => "11111111",
	14248 => "11111111",
	14249 => "11111111",
	14250 => "11111111",
	14251 => "11111111",
	14252 => "11111111",
	14253 => "11111111",
	14254 => "11111111",
	14255 => "11111111",
	14256 => "11111111",
	14257 => "11111111",
	14258 => "11111111",
	14259 => "11111111",
	14260 => "11111111",
	14261 => "11111111",
	14262 => "11111111",
	14263 => "11111111",
	14264 => "11111111",
	14265 => "11111111",
	14266 => "11111111",
	14267 => "11111111",
	14268 => "11111111",
	14269 => "11111111",
	14270 => "11111111",
	14271 => "11111111",
	14272 => "11111111",
	14273 => "11111111",
	14274 => "11111111",
	14275 => "11111111",
	14276 => "11111111",
	14277 => "11111111",
	14278 => "11111111",
	14279 => "11111111",
	14280 => "11111111",
	14281 => "11111111",
	14282 => "11111111",
	14283 => "11111111",
	14284 => "11111111",
	14285 => "11111111",
	14286 => "11111111",
	14287 => "11111111",
	14288 => "11111111",
	14289 => "11111111",
	14290 => "11111111",
	14291 => "11111111",
	14292 => "11111111",
	14293 => "11111111",
	14294 => "11111111",
	14295 => "11111111",
	14296 => "11111111",
	14297 => "11111111",
	14298 => "11111111",
	14299 => "11111111",
	14300 => "11111111",
	14301 => "11111111",
	14302 => "11111111",
	14303 => "11111111",
	14304 => "11111111",
	14305 => "11111111",
	14306 => "11111111",
	14307 => "11111111",
	14308 => "11111111",
	14309 => "11111111",
	14310 => "11111111",
	14311 => "11111111",
	14312 => "11111111",
	14313 => "11111111",
	14314 => "11111111",
	14315 => "11111111",
	14316 => "11111111",
	14317 => "11111111",
	14318 => "11111111",
	14319 => "11111111",
	14320 => "11111111",
	14321 => "11111111",
	14322 => "11111111",
	14323 => "11111111",
	14324 => "11111111",
	14325 => "11111111",
	14326 => "11111111",
	14327 => "11111111",
	14336 => "11111111",
	14337 => "11111111",
	14338 => "11111111",
	14339 => "11111111",
	14340 => "11111111",
	14341 => "11111111",
	14342 => "11111111",
	14343 => "11111111",
	14344 => "11111111",
	14345 => "11111111",
	14346 => "11111111",
	14347 => "11111111",
	14348 => "11111111",
	14349 => "11111111",
	14350 => "11111111",
	14351 => "11111111",
	14352 => "11111111",
	14353 => "11111111",
	14354 => "11111111",
	14355 => "11111111",
	14356 => "11111111",
	14357 => "11111111",
	14358 => "11111111",
	14359 => "11111111",
	14360 => "11111111",
	14361 => "11111111",
	14362 => "11111111",
	14363 => "11111111",
	14364 => "11111111",
	14365 => "11111111",
	14366 => "11111111",
	14367 => "11111111",
	14368 => "11111111",
	14369 => "11111111",
	14370 => "11111111",
	14371 => "11111111",
	14372 => "11111111",
	14373 => "11111111",
	14374 => "11111111",
	14375 => "11111111",
	14376 => "11111111",
	14377 => "11111111",
	14378 => "11111111",
	14379 => "11111111",
	14380 => "11111111",
	14381 => "11111111",
	14382 => "11111111",
	14383 => "11111111",
	14384 => "11111111",
	14385 => "11111111",
	14386 => "11111111",
	14387 => "11111111",
	14388 => "11111111",
	14389 => "11111111",
	14390 => "11111111",
	14391 => "11111111",
	14392 => "11111111",
	14393 => "11111111",
	14394 => "11111111",
	14395 => "11111111",
	14396 => "11111111",
	14397 => "11111111",
	14398 => "11111111",
	14399 => "11111111",
	14400 => "11111111",
	14401 => "11111111",
	14402 => "11111111",
	14403 => "11111111",
	14404 => "11111111",
	14405 => "11111111",
	14406 => "11111111",
	14407 => "11111111",
	14408 => "11111111",
	14409 => "11111111",
	14410 => "11111111",
	14411 => "11111111",
	14412 => "11111111",
	14413 => "11111111",
	14414 => "11111111",
	14415 => "11111111",
	14416 => "11111111",
	14417 => "11111111",
	14418 => "11111111",
	14419 => "11111111",
	14420 => "11111111",
	14421 => "11111111",
	14422 => "11111111",
	14423 => "11111111",
	14424 => "11111111",
	14425 => "11111111",
	14426 => "11111111",
	14427 => "11111111",
	14428 => "11111111",
	14429 => "11111111",
	14430 => "11111111",
	14431 => "11111111",
	14432 => "11111111",
	14433 => "11111111",
	14434 => "11111111",
	14435 => "11111111",
	14436 => "11111111",
	14437 => "11111111",
	14438 => "11111111",
	14439 => "11111111",
	14440 => "11111111",
	14441 => "11111111",
	14442 => "11111111",
	14443 => "11111111",
	14444 => "11111111",
	14445 => "11111111",
	14446 => "11111111",
	14447 => "11111111",
	14448 => "11111111",
	14449 => "11111111",
	14450 => "11111111",
	14451 => "11111111",
	14452 => "11111111",
	14453 => "11111111",
	14454 => "11111111",
	14455 => "11111111",
	14464 => "11111111",
	14465 => "11111111",
	14466 => "11111111",
	14467 => "11111111",
	14468 => "11111111",
	14469 => "11111111",
	14470 => "11111111",
	14471 => "11111111",
	14472 => "11111111",
	14473 => "11111111",
	14474 => "11111111",
	14475 => "11111111",
	14476 => "11111111",
	14477 => "11111111",
	14478 => "11111111",
	14479 => "11111111",
	14480 => "11111111",
	14481 => "11111111",
	14482 => "11111111",
	14483 => "11111111",
	14484 => "11111111",
	14485 => "11111111",
	14486 => "11111111",
	14487 => "11111111",
	14488 => "11111111",
	14489 => "11111111",
	14490 => "11111111",
	14491 => "11111111",
	14492 => "11111111",
	14493 => "11111111",
	14494 => "11111111",
	14495 => "11111111",
	14496 => "11111111",
	14497 => "11111111",
	14498 => "11111111",
	14499 => "11111111",
	14500 => "11111111",
	14501 => "11111111",
	14502 => "11111111",
	14503 => "11111111",
	14504 => "11111111",
	14505 => "11111111",
	14506 => "11111111",
	14507 => "11111111",
	14508 => "11111111",
	14509 => "11111111",
	14510 => "11111111",
	14511 => "11111111",
	14512 => "11111111",
	14513 => "11111111",
	14514 => "11111111",
	14515 => "11111111",
	14516 => "11111111",
	14517 => "11111111",
	14518 => "11111111",
	14519 => "11111111",
	14520 => "11111111",
	14521 => "11111111",
	14522 => "11111111",
	14523 => "11111111",
	14524 => "11111111",
	14525 => "11111111",
	14526 => "11111111",
	14527 => "11111111",
	14528 => "11111111",
	14529 => "11111111",
	14530 => "11111111",
	14531 => "11111111",
	14532 => "11111111",
	14533 => "11111111",
	14534 => "11111111",
	14535 => "11111111",
	14536 => "11111111",
	14537 => "11111111",
	14538 => "11111111",
	14539 => "11111111",
	14540 => "11111111",
	14541 => "11111111",
	14542 => "11111111",
	14543 => "11111111",
	14544 => "11111111",
	14545 => "11111111",
	14546 => "11111111",
	14547 => "11111111",
	14548 => "11111111",
	14549 => "11111111",
	14550 => "11111111",
	14551 => "11111111",
	14552 => "11111111",
	14553 => "11111111",
	14554 => "11111111",
	14555 => "11111111",
	14556 => "11111111",
	14557 => "11111111",
	14558 => "11111111",
	14559 => "11111111",
	14560 => "11111111",
	14561 => "11111111",
	14562 => "11111111",
	14563 => "11111111",
	14564 => "11111111",
	14565 => "11111111",
	14566 => "11111111",
	14567 => "11111111",
	14568 => "11111111",
	14569 => "11111111",
	14570 => "11111111",
	14571 => "11111111",
	14572 => "11111111",
	14573 => "11111111",
	14574 => "11111111",
	14575 => "11111111",
	14576 => "11111111",
	14577 => "11111111",
	14578 => "11111111",
	14579 => "11111111",
	14580 => "11111111",
	14581 => "11111111",
	14582 => "11111111",
	14583 => "11111111",
	14592 => "11111111",
	14593 => "11111111",
	14594 => "11111111",
	14595 => "11111111",
	14596 => "11111111",
	14597 => "11111111",
	14598 => "11111111",
	14599 => "11111111",
	14600 => "11111111",
	14601 => "11111111",
	14602 => "11111111",
	14603 => "11111111",
	14604 => "11111111",
	14605 => "11111111",
	14606 => "11111111",
	14607 => "11111111",
	14608 => "11111111",
	14609 => "11111111",
	14610 => "11111111",
	14611 => "11111111",
	14612 => "11111111",
	14613 => "11111111",
	14614 => "11111111",
	14615 => "11111111",
	14616 => "11111111",
	14617 => "11111111",
	14618 => "11111111",
	14619 => "11111111",
	14620 => "11111111",
	14621 => "11111111",
	14622 => "11111111",
	14623 => "11111111",
	14624 => "11111111",
	14625 => "11111111",
	14626 => "11111111",
	14627 => "11111111",
	14628 => "11111111",
	14629 => "11111111",
	14630 => "11111111",
	14631 => "11111111",
	14632 => "11111111",
	14633 => "11111111",
	14634 => "11111111",
	14635 => "11111111",
	14636 => "11111111",
	14637 => "11111111",
	14638 => "11111111",
	14639 => "11111111",
	14640 => "11111111",
	14641 => "11111111",
	14642 => "11111111",
	14643 => "11111111",
	14644 => "11111111",
	14645 => "11111111",
	14646 => "11111111",
	14647 => "11111111",
	14648 => "11111111",
	14649 => "11111111",
	14650 => "11111111",
	14651 => "11111111",
	14652 => "11111111",
	14653 => "11111111",
	14654 => "11111111",
	14655 => "11111111",
	14656 => "11111111",
	14657 => "11111111",
	14658 => "11111111",
	14659 => "11111111",
	14660 => "11111111",
	14661 => "11111111",
	14662 => "11111111",
	14663 => "11111111",
	14664 => "11111111",
	14665 => "11111111",
	14666 => "11111111",
	14667 => "11111111",
	14668 => "11111111",
	14669 => "11111111",
	14670 => "11111111",
	14671 => "11111111",
	14672 => "11111111",
	14673 => "11111111",
	14674 => "11111111",
	14675 => "11111111",
	14676 => "11111111",
	14677 => "11111111",
	14678 => "11111111",
	14679 => "11111111",
	14680 => "11111111",
	14681 => "11111111",
	14682 => "11111111",
	14683 => "11111111",
	14684 => "11111111",
	14685 => "11111111",
	14686 => "11111111",
	14687 => "11111111",
	14688 => "11111111",
	14689 => "11111111",
	14690 => "11111111",
	14691 => "11111111",
	14692 => "11111111",
	14693 => "11111111",
	14694 => "11111111",
	14695 => "11111111",
	14696 => "11111111",
	14697 => "11111111",
	14698 => "11111111",
	14699 => "11111111",
	14700 => "11111111",
	14701 => "11111111",
	14702 => "11111111",
	14703 => "11111111",
	14704 => "11111111",
	14705 => "11111111",
	14706 => "11111111",
	14707 => "11111111",
	14708 => "11111111",
	14709 => "11111111",
	14710 => "11111111",
	14711 => "11111111",
	14720 => "11111111",
	14721 => "11111111",
	14722 => "11111111",
	14723 => "11111111",
	14724 => "11111111",
	14725 => "11111111",
	14726 => "11111111",
	14727 => "11111111",
	14728 => "11111111",
	14729 => "11111111",
	14730 => "11111111",
	14731 => "11111111",
	14732 => "11111111",
	14733 => "11111111",
	14734 => "11111111",
	14735 => "11111111",
	14736 => "11111111",
	14737 => "11111111",
	14738 => "11111111",
	14739 => "11111111",
	14740 => "11111111",
	14741 => "11111111",
	14742 => "11111111",
	14743 => "11111111",
	14744 => "11111111",
	14745 => "11111111",
	14746 => "11111111",
	14747 => "11111111",
	14748 => "11111111",
	14749 => "11111111",
	14750 => "11111111",
	14751 => "11111111",
	14752 => "11111111",
	14753 => "11111111",
	14754 => "11111111",
	14755 => "11111111",
	14756 => "11111111",
	14757 => "11111111",
	14758 => "11111111",
	14759 => "11111111",
	14760 => "11111111",
	14761 => "11111111",
	14762 => "11111111",
	14763 => "11111111",
	14764 => "11111111",
	14765 => "11111111",
	14766 => "11111111",
	14767 => "11111111",
	14768 => "11111111",
	14769 => "11111111",
	14770 => "11111111",
	14771 => "11111111",
	14772 => "11111111",
	14773 => "11111111",
	14774 => "11111111",
	14775 => "11111111",
	14776 => "11111111",
	14777 => "11111111",
	14778 => "11111111",
	14779 => "11111111",
	14780 => "11111111",
	14781 => "11111111",
	14782 => "11111111",
	14783 => "11111111",
	14784 => "11111111",
	14785 => "11111111",
	14786 => "11111111",
	14787 => "11111111",
	14788 => "11111111",
	14789 => "11111111",
	14790 => "11111111",
	14791 => "11111111",
	14792 => "11111111",
	14793 => "11111111",
	14794 => "11111111",
	14795 => "11111111",
	14796 => "11111111",
	14797 => "11111111",
	14798 => "11111111",
	14799 => "11111111",
	14800 => "11111111",
	14801 => "11111111",
	14802 => "11111111",
	14803 => "11111111",
	14804 => "11111111",
	14805 => "11111111",
	14806 => "11111111",
	14807 => "11111111",
	14808 => "11111111",
	14809 => "11111111",
	14810 => "11111111",
	14811 => "11111111",
	14812 => "11111111",
	14813 => "11111111",
	14814 => "11111111",
	14815 => "11111111",
	14816 => "11111111",
	14817 => "11111111",
	14818 => "11111111",
	14819 => "11111111",
	14820 => "11111111",
	14821 => "11111111",
	14822 => "11111111",
	14823 => "11111111",
	14824 => "11111111",
	14825 => "11111111",
	14826 => "11111111",
	14827 => "11111111",
	14828 => "11111111",
	14829 => "11111111",
	14830 => "11111111",
	14831 => "11111111",
	14832 => "11111111",
	14833 => "11111111",
	14834 => "11111111",
	14835 => "11111111",
	14836 => "11111111",
	14837 => "11111111",
	14838 => "11111111",
	14839 => "11111111",
	14848 => "11111111",
	14849 => "11111111",
	14850 => "11111111",
	14851 => "11111111",
	14852 => "11111111",
	14853 => "11111111",
	14854 => "11111111",
	14855 => "11111111",
	14856 => "11111111",
	14857 => "11111111",
	14858 => "11111111",
	14859 => "11111111",
	14860 => "11111111",
	14861 => "11111111",
	14862 => "11111111",
	14863 => "11111111",
	14864 => "11111111",
	14865 => "11111111",
	14866 => "11111111",
	14867 => "11111111",
	14868 => "11111111",
	14869 => "11111111",
	14870 => "11111111",
	14871 => "11111111",
	14872 => "11111111",
	14873 => "11111111",
	14874 => "11111111",
	14875 => "11111111",
	14876 => "11111111",
	14877 => "11111111",
	14878 => "11111111",
	14879 => "11111111",
	14880 => "11111111",
	14881 => "11111111",
	14882 => "11111111",
	14883 => "11111111",
	14884 => "11111111",
	14885 => "11111111",
	14886 => "11111111",
	14887 => "11111111",
	14888 => "11111111",
	14889 => "11111111",
	14890 => "11111111",
	14891 => "11111111",
	14892 => "11111111",
	14893 => "11111111",
	14894 => "11111111",
	14895 => "11111111",
	14896 => "11111111",
	14897 => "11111111",
	14898 => "11111111",
	14899 => "11111111",
	14900 => "11111111",
	14901 => "11111111",
	14902 => "11111111",
	14903 => "11111111",
	14904 => "11111111",
	14905 => "11111111",
	14906 => "11111111",
	14907 => "11111111",
	14908 => "11111111",
	14909 => "11111111",
	14910 => "11111111",
	14911 => "11111111",
	14912 => "11111111",
	14913 => "11111111",
	14914 => "11111111",
	14915 => "11111111",
	14916 => "11111111",
	14917 => "11111111",
	14918 => "11111111",
	14919 => "11111111",
	14920 => "11111111",
	14921 => "11111111",
	14922 => "11111111",
	14923 => "11111111",
	14924 => "11111111",
	14925 => "11111111",
	14926 => "11111111",
	14927 => "11111111",
	14928 => "11111111",
	14929 => "11111111",
	14930 => "11111111",
	14931 => "11111111",
	14932 => "11111111",
	14933 => "11111111",
	14934 => "11111111",
	14935 => "11111111",
	14936 => "11111111",
	14937 => "11111111",
	14938 => "11111111",
	14939 => "11111111",
	14940 => "11111111",
	14941 => "11111111",
	14942 => "11111111",
	14943 => "11111111",
	14944 => "11111111",
	14945 => "11111111",
	14946 => "11111111",
	14947 => "11111111",
	14948 => "11111111",
	14949 => "11111111",
	14950 => "11111111",
	14951 => "11111111",
	14952 => "11111111",
	14953 => "11111111",
	14954 => "11111111",
	14955 => "11111111",
	14956 => "11111111",
	14957 => "11111111",
	14958 => "11111111",
	14959 => "11111111",
	14960 => "11111111",
	14961 => "11111111",
	14962 => "11111111",
	14963 => "11111111",
	14964 => "11111111",
	14965 => "11111111",
	14966 => "11111111",
	14967 => "11111111",
	14976 => "11111111",
	14977 => "11111111",
	14978 => "11111111",
	14979 => "11111111",
	14980 => "11111111",
	14981 => "11111111",
	14982 => "11111111",
	14983 => "11111111",
	14984 => "11111111",
	14985 => "11111111",
	14986 => "11111111",
	14987 => "11111111",
	14988 => "11111111",
	14989 => "11111111",
	14990 => "11111111",
	14991 => "11111111",
	14992 => "11111111",
	14993 => "11111111",
	14994 => "11111111",
	14995 => "11111111",
	14996 => "11111111",
	14997 => "11111111",
	14998 => "11111111",
	14999 => "11111111",
	15000 => "11111111",
	15001 => "11111111",
	15002 => "11111111",
	15003 => "11111111",
	15004 => "11111111",
	15005 => "11111111",
	15006 => "11111111",
	15007 => "11111111",
	15008 => "11111111",
	15009 => "11111111",
	15010 => "11111111",
	15011 => "11111111",
	15012 => "11111111",
	15013 => "11111111",
	15014 => "11111111",
	15015 => "11111111",
	15016 => "11111111",
	15017 => "11111111",
	15018 => "11111111",
	15019 => "11111111",
	15020 => "11111111",
	15021 => "11111111",
	15022 => "11111111",
	15023 => "11111111",
	15024 => "11111111",
	15025 => "11111111",
	15026 => "11111111",
	15027 => "11111111",
	15028 => "11111111",
	15029 => "11111111",
	15030 => "11111111",
	15031 => "11111111",
	15032 => "11111111",
	15033 => "11111111",
	15034 => "11111111",
	15035 => "11111111",
	15036 => "11111111",
	15037 => "11111111",
	15038 => "11111111",
	15039 => "11111111",
	15040 => "11111111",
	15041 => "11111111",
	15042 => "11111111",
	15043 => "11111111",
	15044 => "11111111",
	15045 => "11111111",
	15046 => "11111111",
	15047 => "11111111",
	15048 => "11111111",
	15049 => "11111111",
	15050 => "11111111",
	15051 => "11111111",
	15052 => "11111111",
	15053 => "11111111",
	15054 => "11111111",
	15055 => "11111111",
	15056 => "11111111",
	15057 => "11111111",
	15058 => "11111111",
	15059 => "11111111",
	15060 => "11111111",
	15061 => "11111111",
	15062 => "11111111",
	15063 => "11111111",
	15064 => "11111111",
	15065 => "11111111",
	15066 => "11111111",
	15067 => "11111111",
	15068 => "11111111",
	15069 => "11111111",
	15070 => "11111111",
	15071 => "11111111",
	15072 => "11111111",
	15073 => "11111111",
	15074 => "11111111",
	15075 => "11111111",
	15076 => "11111111",
	15077 => "11111111",
	15078 => "11111111",
	15079 => "11111111",
	15080 => "11111111",
	15081 => "11111111",
	15082 => "11111111",
	15083 => "11111111",
	15084 => "11111111",
	15085 => "11111111",
	15086 => "11111111",
	15087 => "11111111",
	15088 => "11111111",
	15089 => "11111111",
	15090 => "11111111",
	15091 => "11111111",
	15092 => "11111111",
	15093 => "11111111",
	15094 => "11111111",
	15095 => "11111111",
	15104 => "11111111",
	15105 => "11111111",
	15106 => "11111111",
	15107 => "11111111",
	15108 => "11111111",
	15109 => "11111111",
	15110 => "11111111",
	15111 => "11111111",
	15112 => "11111111",
	15113 => "11111111",
	15114 => "11111111",
	15115 => "11111111",
	15116 => "11111111",
	15117 => "11111111",
	15118 => "11111111",
	15119 => "11111111",
	15120 => "11111111",
	15121 => "11111111",
	15122 => "11111111",
	15123 => "11111111",
	15124 => "11111111",
	15125 => "11111111",
	15126 => "11111111",
	15127 => "11111111",
	15128 => "11111111",
	15129 => "11111111",
	15130 => "11111111",
	15131 => "11111111",
	15132 => "11111111",
	15133 => "11111111",
	15134 => "11111111",
	15135 => "11111111",
	15136 => "11111111",
	15137 => "11111111",
	15138 => "11111111",
	15139 => "11111111",
	15140 => "11111111",
	15141 => "11111111",
	15142 => "11111111",
	15143 => "11111111",
	15144 => "11111111",
	15145 => "11111111",
	15146 => "11111111",
	15147 => "11111111",
	15148 => "11111111",
	15149 => "11111111",
	15150 => "11111111",
	15151 => "11111111",
	15152 => "11111111",
	15153 => "11111111",
	15154 => "11111111",
	15155 => "11111111",
	15156 => "11111111",
	15157 => "11111111",
	15158 => "11111111",
	15159 => "11111111",
	15160 => "11111111",
	15161 => "11111111",
	15162 => "11111111",
	15163 => "11111111",
	15164 => "11111111",
	15165 => "11111111",
	15166 => "11111111",
	15167 => "11111111",
	15168 => "11111111",
	15169 => "11111111",
	15170 => "11111111",
	15171 => "11111111",
	15172 => "11111111",
	15173 => "11111111",
	15174 => "11111111",
	15175 => "11111111",
	15176 => "11111111",
	15177 => "11111111",
	15178 => "11111111",
	15179 => "11111111",
	15180 => "11111111",
	15181 => "11111111",
	15182 => "11111111",
	15183 => "11111111",
	15184 => "11111111",
	15185 => "11111111",
	15186 => "11111111",
	15187 => "11111111",
	15188 => "11111111",
	15189 => "11111111",
	15190 => "11111111",
	15191 => "11111111",
	15192 => "11111111",
	15193 => "11111111",
	15194 => "11111111",
	15195 => "11111111",
	15196 => "11111111",
	15197 => "11111111",
	15198 => "11111111",
	15199 => "11111111",
	15200 => "11111111",
	15201 => "11111111",
	15202 => "11111111",
	15203 => "11111111",
	15204 => "11111111",
	15205 => "11111111",
	15206 => "11111111",
	15207 => "11111111",
	15208 => "11111111",
	15209 => "11111111",
	15210 => "11111111",
	15211 => "11111111",
	15212 => "11111111",
	15213 => "11111111",
	15214 => "11111111",
	15215 => "11111111",
	15216 => "11111111",
	15217 => "11111111",
	15218 => "11111111",
	15219 => "11111111",
	15220 => "11111111",
	15221 => "11111111",
	15222 => "11111111",
	15223 => "11111111",
	15232 => "11111111",
	15233 => "11111111",
	15234 => "11111111",
	15235 => "11111111",
	15236 => "11111111",
	15237 => "11111111",
	15238 => "11111111",
	15239 => "11111111",
	15240 => "11111111",
	15241 => "11111111",
	15242 => "11111111",
	15243 => "11111111",
	15244 => "11111111",
	15245 => "11111111",
	15246 => "11111111",
	15247 => "11111111",
	15248 => "11111111",
	15249 => "11111111",
	15250 => "11111111",
	15251 => "11111111",
	15252 => "11111111",
	15253 => "11111111",
	15254 => "11111111",
	15255 => "11111111",
	15256 => "11111111",
	15257 => "11111111",
	15258 => "11111111",
	15259 => "11111111",
	15260 => "11111111",
	15261 => "11111111",
	15262 => "11111111",
	15263 => "11111111",
	15264 => "11111111",
	15265 => "11111111",
	15266 => "11111111",
	15267 => "11111111",
	15268 => "11111111",
	15269 => "11111111",
	15270 => "11111111",
	15271 => "11111111",
	15272 => "11111111",
	15273 => "11111111",
	15274 => "11111111",
	15275 => "11111111",
	15276 => "11111111",
	15277 => "11111111",
	15278 => "11111111",
	15279 => "11111111",
	15280 => "11111111",
	15281 => "11111111",
	15282 => "11111111",
	15283 => "11111111",
	15284 => "11111111",
	15285 => "11111111",
	15286 => "11111111",
	15287 => "11111111",
	15288 => "11111111",
	15289 => "11111111",
	15290 => "11111111",
	15291 => "11111111",
	15292 => "11111111",
	15293 => "11111111",
	15294 => "11111111",
	15295 => "11111111",
	15296 => "11111111",
	15297 => "11111111",
	15298 => "11111111",
	15299 => "11111111",
	15300 => "11111111",
	15301 => "11111111",
	15302 => "11111111",
	15303 => "11111111",
	15304 => "11111111",
	15305 => "11111111",
	15306 => "11111111",
	15307 => "11111111",
	15308 => "11111111",
	15309 => "11111111",
	15310 => "11111111",
	15311 => "11111111",
	15312 => "11111111",
	15313 => "11111111",
	15314 => "11111111",
	15315 => "11111111",
	15316 => "11111111",
	15317 => "11111111",
	15318 => "11111111",
	15319 => "11111111",
	15320 => "11111111",
	15321 => "11111111",
	15322 => "11111111",
	15323 => "11111111",
	15324 => "11111111",
	15325 => "11111111",
	15326 => "11111111",
	15327 => "11111111",
	15328 => "11111111",
	15329 => "11111111",
	15330 => "11111111",
	15331 => "11111111",
	15332 => "11111111",
	15333 => "11111111",
	15334 => "11111111",
	15335 => "11111111",
	15336 => "11111111",
	15337 => "11111111",
	15338 => "11111111",
	15339 => "11111111",
	15340 => "11111111",
	15341 => "11111111",
	15342 => "11111111",
	15343 => "11111111",
	15344 => "11111111",
	15345 => "11111111",
	15346 => "11111111",
	15347 => "11111111",
	15348 => "11111111",
	15349 => "11111111",
	15350 => "11111111",
	15351 => "11111111",
	15360 => "11111111",
	15361 => "11111111",
	15362 => "11111111",
	15363 => "11111111",
	15364 => "11111111",
	15365 => "11111111",
	15366 => "11111111",
	15367 => "11111111",
	15368 => "11111111",
	15369 => "11111111",
	15370 => "11111111",
	15371 => "11111111",
	15372 => "11111111",
	15373 => "11111111",
	15374 => "11111111",
	15375 => "11111111",
	15376 => "11111111",
	15377 => "11111111",
	15378 => "11111111",
	15379 => "11111111",
	15380 => "11111111",
	15381 => "11111111",
	15382 => "11111111",
	15383 => "11111111",
	15384 => "11111111",
	15385 => "11111111",
	15386 => "11111111",
	15387 => "11111111",
	15388 => "11111111",
	15389 => "11111111",
	15390 => "11111111",
	15391 => "11111111",
	15392 => "11111111",
	15393 => "11111111",
	15394 => "11111111",
	15395 => "11111111",
	15396 => "11111111",
	15397 => "11111111",
	15398 => "11111111",
	15399 => "11111111",
	15400 => "11111111",
	15401 => "11111111",
	15402 => "11111111",
	15403 => "11111111",
	15404 => "11111111",
	15405 => "11111111",
	15406 => "11111111",
	15407 => "11111111",
	15408 => "11111111",
	15409 => "11111111",
	15410 => "11111111",
	15411 => "11111111",
	15412 => "11111111",
	15413 => "11111111",
	15414 => "11111111",
	15415 => "11111111",
	15416 => "11111111",
	15417 => "11111111",
	15418 => "11111111",
	15419 => "11111111",
	15420 => "11111111",
	15421 => "11111111",
	15422 => "11111111",
	15423 => "11111111",
	15424 => "11111111",
	15425 => "11111111",
	15426 => "11111111",
	15427 => "11111111",
	15428 => "11111111",
	15429 => "11111111",
	15430 => "11111111",
	15431 => "11111111",
	15432 => "11111111",
	15433 => "11111111",
	15434 => "11111111",
	15435 => "11111111",
	15436 => "11111111",
	15437 => "11111111",
	15438 => "11111111",
	15439 => "11111111",
	15440 => "11111111",
	15441 => "11111111",
	15442 => "11111111",
	15443 => "11111111",
	15444 => "11111111",
	15445 => "11111111",
	15446 => "11111111",
	15447 => "11111111",
	15448 => "11111111",
	15449 => "11111111",
	15450 => "11111111",
	15451 => "11111111",
	15452 => "11111111",
	15453 => "11111111",
	15454 => "11111111",
	15455 => "11111111",
	15456 => "11111111",
	15457 => "11111111",
	15458 => "11111111",
	15459 => "11111111",
	15460 => "11111111",
	15461 => "11111111",
	15462 => "11111111",
	15463 => "11111111",
	15464 => "11111111",
	15465 => "11111111",
	15466 => "11111111",
	15467 => "11111111",
	15468 => "11111111",
	15469 => "11111111",
	15470 => "11111111",
	15471 => "11111111",
	15472 => "11111111",
	15473 => "11111111",
	15474 => "11111111",
	15475 => "11111111",
	15476 => "11111111",
	15477 => "11111111",
	15478 => "11111111",
	15479 => "11111111",

	others => (others => '0')
);

begin
	
	-- process ROM
	process (CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (EN = '1') then
				DATA <= ROM(conv_integer(ADDR));
			end if;
		end if;
	end process;
	
end Behavioral;

