----------------------------------------------------------------------------------
-- Company: Ensimag 
-- Engineer: S. Viardot
-- 
-- Create Date:    14:13:14 11/24/2008 
-- Design Name: 
-- Module Name:    ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: Memoire Video
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM is
    Port ( AD : in  STD_LOGIC_VECTOR (12 downto 0);
           D : out  STD_LOGIC_VECTOR (15 downto 0);
           CLK : in STD_LOGIC
			  );
end ROM;

architecture Behavioral of ROM is
 constant low_address: natural := 0;
 constant high_address: natural := 8192;  
 subtype octet is std_logic_vector( 15 downto 0 );
 type zone_memoire is
         array (natural range low_address to high_address) of octet;
 signal m: zone_memoire;
begin
m(0)<=x"0000";
m(1)<=x"0000";
m(2)<=x"0000";
m(3)<=x"0000";
m(4)<=x"0000";
m(5)<=x"0000";
m(6)<=x"0080";
m(7)<=x"0000";
m(8)<=x"0000";
m(9)<=x"0000";
m(10)<=x"0000";
m(11)<=x"0000";
m(12)<=x"1000";
m(32)<=x"0000";
m(33)<=x"0000";
m(34)<=x"0000";
m(35)<=x"0000";
m(36)<=x"0000";
m(37)<=x"0000";
m(38)<=x"0100";
m(39)<=x"0000";
m(40)<=x"0000";
m(41)<=x"0000";
m(42)<=x"0000";
m(43)<=x"0000";
m(44)<=x"0000";
m(64)<=x"0000";
m(65)<=x"0000";
m(66)<=x"0000";
m(67)<=x"0000";
m(68)<=x"0000";
m(69)<=x"0000";
m(70)<=x"00e8";
m(71)<=x"0000";
m(72)<=x"0000";
m(73)<=x"0000";
m(74)<=x"0000";
m(75)<=x"0000";
m(76)<=x"0000";
m(96)<=x"0000";
m(97)<=x"0000";
m(98)<=x"0000";
m(99)<=x"0000";
m(100)<=x"0000";
m(101)<=x"0000";
m(102)<=x"0006";
m(103)<=x"0000";
m(104)<=x"0000";
m(105)<=x"0000";
m(106)<=x"0000";
m(107)<=x"0000";
m(108)<=x"0000";
m(128)<=x"0000";
m(129)<=x"0000";
m(130)<=x"0000";
m(131)<=x"0000";
m(132)<=x"0000";
m(133)<=x"0000";
m(134)<=x"0046";
m(135)<=x"0000";
m(136)<=x"0000";
m(137)<=x"0000";
m(138)<=x"0000";
m(139)<=x"0000";
m(140)<=x"0000";
m(160)<=x"0000";
m(161)<=x"0000";
m(162)<=x"0000";
m(163)<=x"0000";
m(164)<=x"0000";
m(165)<=x"0000";
m(166)<=x"9412";
m(167)<=x"2000";
m(168)<=x"0000";
m(169)<=x"0000";
m(170)<=x"0000";
m(171)<=x"0000";
m(172)<=x"0000";
m(192)<=x"0000";
m(193)<=x"0000";
m(194)<=x"0000";
m(195)<=x"0000";
m(196)<=x"0000";
m(197)<=x"000c";
m(198)<=x"2266";
m(199)<=x"2000";
m(200)<=x"0000";
m(201)<=x"0000";
m(202)<=x"0000";
m(203)<=x"0000";
m(204)<=x"0000";
m(224)<=x"0000";
m(225)<=x"0000";
m(226)<=x"0000";
m(227)<=x"0000";
m(228)<=x"0000";
m(229)<=x"0000";
m(230)<=x"0c18";
m(231)<=x"0000";
m(232)<=x"0000";
m(233)<=x"0000";
m(234)<=x"0000";
m(235)<=x"0000";
m(236)<=x"0000";
m(256)<=x"0000";
m(257)<=x"0000";
m(258)<=x"0000";
m(259)<=x"0000";
m(260)<=x"0000";
m(261)<=x"0002";
m(262)<=x"8c36";
m(263)<=x"2000";
m(264)<=x"0000";
m(265)<=x"0000";
m(266)<=x"0000";
m(267)<=x"0000";
m(268)<=x"0000";
m(288)<=x"0000";
m(289)<=x"0000";
m(290)<=x"0000";
m(291)<=x"0000";
m(292)<=x"0000";
m(293)<=x"0059";
m(294)<=x"610d";
m(295)<=x"d900";
m(296)<=x"0000";
m(297)<=x"0000";
m(298)<=x"0000";
m(299)<=x"0000";
m(300)<=x"0000";
m(320)<=x"0000";
m(321)<=x"0000";
m(322)<=x"0000";
m(323)<=x"0000";
m(324)<=x"0000";
m(325)<=x"0801";
m(326)<=x"4019";
m(327)<=x"e500";
m(328)<=x"0000";
m(329)<=x"0000";
m(330)<=x"0000";
m(331)<=x"0000";
m(332)<=x"0000";
m(352)<=x"0000";
m(353)<=x"0000";
m(354)<=x"0000";
m(355)<=x"0000";
m(356)<=x"0000";
m(357)<=x"1102";
m(358)<=x"08da";
m(359)<=x"a910";
m(360)<=x"0000";
m(361)<=x"0000";
m(362)<=x"0000";
m(363)<=x"0000";
m(364)<=x"0000";
m(384)<=x"0000";
m(385)<=x"0000";
m(386)<=x"0000";
m(387)<=x"0000";
m(388)<=x"0000";
m(389)<=x"0822";
m(390)<=x"29bd";
m(391)<=x"e788";
m(392)<=x"0000";
m(393)<=x"0000";
m(394)<=x"0000";
m(395)<=x"0000";
m(396)<=x"0000";
m(416)<=x"0000";
m(417)<=x"0000";
m(418)<=x"0000";
m(419)<=x"0000";
m(420)<=x"0160";
m(421)<=x"8301";
m(422)<=x"197b";
m(423)<=x"7e90";
m(424)<=x"0000";
m(425)<=x"0000";
m(426)<=x"0000";
m(427)<=x"0000";
m(428)<=x"0000";
m(448)<=x"0000";
m(449)<=x"0000";
m(450)<=x"0000";
m(451)<=x"0000";
m(452)<=x"0798";
m(453)<=x"0126";
m(454)<=x"a8ff";
m(455)<=x"ba00";
m(456)<=x"0000";
m(457)<=x"0000";
m(458)<=x"0000";
m(459)<=x"0000";
m(460)<=x"0000";
m(480)<=x"0000";
m(481)<=x"0000";
m(482)<=x"0000";
m(483)<=x"0000";
m(484)<=x"29f9";
m(485)<=x"48e3";
m(486)<=x"35f9";
m(487)<=x"ff70";
m(488)<=x"0000";
m(489)<=x"0000";
m(490)<=x"0000";
m(491)<=x"0000";
m(492)<=x"0000";
m(512)<=x"0000";
m(513)<=x"0000";
m(514)<=x"0000";
m(515)<=x"0000";
m(516)<=x"8dbf";
m(517)<=x"b5e6";
m(518)<=x"effe";
m(519)<=x"7fd0";
m(520)<=x"0000";
m(521)<=x"0000";
m(522)<=x"0000";
m(523)<=x"0000";
m(524)<=x"0000";
m(544)<=x"0000";
m(545)<=x"0000";
m(546)<=x"0000";
m(547)<=x"0001";
m(548)<=x"47f7";
m(549)<=x"db7f";
m(550)<=x"b7fd";
m(551)<=x"ffa4";
m(552)<=x"0000";
m(553)<=x"0000";
m(554)<=x"0000";
m(555)<=x"0000";
m(556)<=x"0000";
m(576)<=x"0000";
m(577)<=x"0000";
m(578)<=x"0000";
m(579)<=x"0008";
m(580)<=x"3dff";
m(581)<=x"ddfe";
m(582)<=x"77ff";
m(583)<=x"7fc6";
m(584)<=x"0000";
m(585)<=x"0000";
m(586)<=x"0000";
m(587)<=x"0000";
m(588)<=x"0000";
m(608)<=x"0000";
m(609)<=x"0000";
m(610)<=x"0000";
m(611)<=x"0002";
m(612)<=x"b77e";
m(613)<=x"fbff";
m(614)<=x"ffff";
m(615)<=x"ffb2";
m(616)<=x"0000";
m(617)<=x"0000";
m(618)<=x"0000";
m(619)<=x"0000";
m(620)<=x"0000";
m(640)<=x"0000";
m(641)<=x"0000";
m(642)<=x"0000";
m(643)<=x"0037";
m(644)<=x"ffff";
m(645)<=x"bfff";
m(646)<=x"ffff";
m(647)<=x"fff8";
m(648)<=x"000a";
m(649)<=x"3800";
m(650)<=x"0000";
m(651)<=x"0000";
m(652)<=x"0000";
m(672)<=x"0000";
m(673)<=x"0000";
m(674)<=x"0000";
m(675)<=x"006e";
m(676)<=x"ded7";
m(677)<=x"f7ff";
m(678)<=x"ffff";
m(679)<=x"ffa6";
m(680)<=x"8115";
m(681)<=x"4200";
m(682)<=x"0000";
m(683)<=x"0000";
m(684)<=x"0000";
m(704)<=x"0000";
m(705)<=x"0000";
m(706)<=x"0000";
m(707)<=x"046d";
m(708)<=x"ffbd";
m(709)<=x"efff";
m(710)<=x"ffff";
m(711)<=x"ff7c";
m(712)<=x"1120";
m(713)<=x"0000";
m(714)<=x"0000";
m(715)<=x"0000";
m(716)<=x"0000";
m(736)<=x"0000";
m(737)<=x"0000";
m(738)<=x"0000";
m(739)<=x"03b7";
m(740)<=x"b5ef";
m(741)<=x"f3ff";
m(742)<=x"ffff";
m(743)<=x"ffe1";
m(744)<=x"0704";
m(745)<=x"0000";
m(746)<=x"0000";
m(747)<=x"0000";
m(748)<=x"0000";
m(768)<=x"0000";
m(769)<=x"0000";
m(770)<=x"0000";
m(771)<=x"0bf5";
m(772)<=x"feef";
m(773)<=x"bfff";
m(774)<=x"ffff";
m(775)<=x"ff91";
m(776)<=x"bb20";
m(777)<=x"0000";
m(778)<=x"0000";
m(779)<=x"0000";
m(780)<=x"0000";
m(800)<=x"0000";
m(801)<=x"0000";
m(802)<=x"0000";
m(803)<=x"225f";
m(804)<=x"f7ff";
m(805)<=x"ffff";
m(806)<=x"ffff";
m(807)<=x"ffed";
m(808)<=x"fbd8";
m(809)<=x"1100";
m(810)<=x"0000";
m(811)<=x"0000";
m(812)<=x"0000";
m(832)<=x"0000";
m(833)<=x"0000";
m(834)<=x"0000";
m(835)<=x"0ebb";
m(836)<=x"efbf";
m(837)<=x"ffff";
m(838)<=x"ffff";
m(839)<=x"fffb";
m(840)<=x"fea6";
m(841)<=x"067a";
m(842)<=x"0000";
m(843)<=x"0000";
m(844)<=x"0000";
m(864)<=x"0000";
m(865)<=x"0000";
m(866)<=x"0000";
m(867)<=x"124f";
m(868)<=x"ffff";
m(869)<=x"ffff";
m(870)<=x"ffff";
m(871)<=x"fff5";
m(872)<=x"ffc8";
m(873)<=x"6e47";
m(874)<=x"0000";
m(875)<=x"0000";
m(876)<=x"0000";
m(896)<=x"0000";
m(897)<=x"0000";
m(898)<=x"0000";
m(899)<=x"0a7f";
m(900)<=x"deff";
m(901)<=x"ffff";
m(902)<=x"ffff";
m(903)<=x"ffff";
m(904)<=x"ffb5";
m(905)<=x"d340";
m(906)<=x"6000";
m(907)<=x"0000";
m(908)<=x"0000";
m(928)<=x"0000";
m(929)<=x"0000";
m(930)<=x"0000";
m(931)<=x"0065";
m(932)<=x"ffdf";
m(933)<=x"ffff";
m(934)<=x"ffff";
m(935)<=x"ffff";
m(936)<=x"ffff";
m(937)<=x"fe98";
m(938)<=x"0000";
m(939)<=x"0000";
m(940)<=x"0000";
m(960)<=x"0000";
m(961)<=x"0000";
m(962)<=x"0000";
m(963)<=x"196f";
m(964)<=x"fbff";
m(965)<=x"ffff";
m(966)<=x"ffff";
m(967)<=x"ffff";
m(968)<=x"ffff";
m(969)<=x"e8eb";
m(970)<=x"4000";
m(971)<=x"0000";
m(972)<=x"0000";
m(992)<=x"0000";
m(993)<=x"0000";
m(994)<=x"0000";
m(995)<=x"407d";
m(996)<=x"7fff";
m(997)<=x"ffff";
m(998)<=x"ffff";
m(999)<=x"ffff";
m(1000)<=x"fffa";
m(1001)<=x"e409";
m(1002)<=x"9000";
m(1003)<=x"0000";
m(1004)<=x"0000";
m(1024)<=x"0000";
m(1025)<=x"0000";
m(1026)<=x"0000";
m(1027)<=x"01bf";
m(1028)<=x"ffff";
m(1029)<=x"ffff";
m(1030)<=x"ffff";
m(1031)<=x"ffff";
m(1032)<=x"ffff";
m(1033)<=x"ff00";
m(1034)<=x"0200";
m(1035)<=x"0000";
m(1036)<=x"0000";
m(1056)<=x"0000";
m(1057)<=x"0000";
m(1058)<=x"0000";
m(1059)<=x"01fb";
m(1060)<=x"bfff";
m(1061)<=x"ffff";
m(1062)<=x"ffff";
m(1063)<=x"ffff";
m(1064)<=x"ffff";
m(1065)<=x"ffa2";
m(1066)<=x"0000";
m(1067)<=x"0000";
m(1068)<=x"0000";
m(1088)<=x"0000";
m(1089)<=x"0000";
m(1090)<=x"0000";
m(1091)<=x"0bef";
m(1092)<=x"bfff";
m(1093)<=x"ffff";
m(1094)<=x"ffff";
m(1095)<=x"ffff";
m(1096)<=x"ffff";
m(1097)<=x"ffe0";
m(1098)<=x"0000";
m(1099)<=x"0000";
m(1100)<=x"0000";
m(1120)<=x"0000";
m(1121)<=x"0000";
m(1122)<=x"0000";
m(1123)<=x"3fbc";
m(1124)<=x"dfff";
m(1125)<=x"ffff";
m(1126)<=x"ffff";
m(1127)<=x"ffff";
m(1128)<=x"ffff";
m(1129)<=x"fff0";
m(1130)<=x"0000";
m(1131)<=x"0000";
m(1132)<=x"0000";
m(1152)<=x"0000";
m(1153)<=x"0000";
m(1154)<=x"0000";
m(1155)<=x"5edb";
m(1156)<=x"ffff";
m(1157)<=x"ffff";
m(1158)<=x"ffff";
m(1159)<=x"ffff";
m(1160)<=x"ffff";
m(1161)<=x"fff0";
m(1162)<=x"0100";
m(1163)<=x"0000";
m(1164)<=x"0000";
m(1184)<=x"0000";
m(1185)<=x"0000";
m(1186)<=x"0000";
m(1187)<=x"27bf";
m(1188)<=x"afff";
m(1189)<=x"ffff";
m(1190)<=x"ffff";
m(1191)<=x"ffff";
m(1192)<=x"ffff";
m(1193)<=x"fffe";
m(1194)<=x"0000";
m(1195)<=x"0000";
m(1196)<=x"0000";
m(1216)<=x"0000";
m(1217)<=x"0000";
m(1218)<=x"0000";
m(1219)<=x"dd7f";
m(1220)<=x"ffff";
m(1221)<=x"ffff";
m(1222)<=x"ffff";
m(1223)<=x"ffff";
m(1224)<=x"ffff";
m(1225)<=x"fffe";
m(1226)<=x"8000";
m(1227)<=x"0000";
m(1228)<=x"0000";
m(1248)<=x"0000";
m(1249)<=x"0000";
m(1250)<=x"0010";
m(1251)<=x"4fd6";
m(1252)<=x"dfff";
m(1253)<=x"ffff";
m(1254)<=x"ffff";
m(1255)<=x"ffff";
m(1256)<=x"ffff";
m(1257)<=x"ffff";
m(1258)<=x"2a40";
m(1259)<=x"0000";
m(1260)<=x"0000";
m(1280)<=x"0000";
m(1281)<=x"0000";
m(1282)<=x"0001";
m(1283)<=x"7fdb";
m(1284)<=x"f7ff";
m(1285)<=x"ffff";
m(1286)<=x"ffff";
m(1287)<=x"ffff";
m(1288)<=x"ffff";
m(1289)<=x"ffff";
m(1290)<=x"bd20";
m(1291)<=x"0000";
m(1292)<=x"0000";
m(1312)<=x"0000";
m(1313)<=x"0000";
m(1314)<=x"000e";
m(1315)<=x"fe7f";
m(1316)<=x"ffff";
m(1317)<=x"ffff";
m(1318)<=x"ffff";
m(1319)<=x"ffff";
m(1320)<=x"ffff";
m(1321)<=x"ffff";
m(1322)<=x"f604";
m(1323)<=x"0000";
m(1324)<=x"0000";
m(1344)<=x"0000";
m(1345)<=x"0000";
m(1346)<=x"001f";
m(1347)<=x"f5dd";
m(1348)<=x"dfff";
m(1349)<=x"ffff";
m(1350)<=x"ffff";
m(1351)<=x"ffff";
m(1352)<=x"ffff";
m(1353)<=x"ffff";
m(1354)<=x"ff90";
m(1355)<=x"0000";
m(1356)<=x"0000";
m(1376)<=x"0000";
m(1377)<=x"0000";
m(1378)<=x"003d";
m(1379)<=x"ff7f";
m(1380)<=x"fdff";
m(1381)<=x"ffff";
m(1382)<=x"ffff";
m(1383)<=x"ffff";
m(1384)<=x"ffff";
m(1385)<=x"ffff";
m(1386)<=x"ff88";
m(1387)<=x"0000";
m(1388)<=x"0000";
m(1408)<=x"0000";
m(1409)<=x"0000";
m(1410)<=x"03f6";
m(1411)<=x"e6ef";
m(1412)<=x"fdff";
m(1413)<=x"ffff";
m(1414)<=x"ffff";
m(1415)<=x"ffff";
m(1416)<=x"ffff";
m(1417)<=x"ffff";
m(1418)<=x"fee4";
m(1419)<=x"0000";
m(1420)<=x"0000";
m(1440)<=x"0000";
m(1441)<=x"0000";
m(1442)<=x"0fdf";
m(1443)<=x"9db9";
m(1444)<=x"77ff";
m(1445)<=x"ffdd";
m(1446)<=x"ffef";
m(1447)<=x"ffff";
m(1448)<=x"ffff";
m(1449)<=x"ffff";
m(1450)<=x"f9e2";
m(1451)<=x"0000";
m(1452)<=x"0000";
m(1472)<=x"0000";
m(1473)<=x"0000";
m(1474)<=x"0b7f";
m(1475)<=x"fbfe";
m(1476)<=x"edff";
m(1477)<=x"ffff";
m(1478)<=x"fffe";
m(1479)<=x"ffff";
m(1480)<=x"ffff";
m(1481)<=x"ffff";
m(1482)<=x"ff18";
m(1483)<=x"0000";
m(1484)<=x"0000";
m(1504)<=x"0000";
m(1505)<=x"0000";
m(1506)<=x"06de";
m(1507)<=x"6edf";
m(1508)<=x"feff";
m(1509)<=x"fffd";
m(1510)<=x"ffff";
m(1511)<=x"ffff";
m(1512)<=x"ffff";
m(1513)<=x"ffff";
m(1514)<=x"fe58";
m(1515)<=x"0000";
m(1516)<=x"0000";
m(1536)<=x"0000";
m(1537)<=x"0000";
m(1538)<=x"1ffb";
m(1539)<=x"5bef";
m(1540)<=x"feff";
m(1541)<=x"fffb";
m(1542)<=x"feff";
m(1543)<=x"ffff";
m(1544)<=x"ffff";
m(1545)<=x"ffff";
m(1546)<=x"fa14";
m(1547)<=x"0000";
m(1548)<=x"0000";
m(1568)<=x"0000";
m(1569)<=x"0000";
m(1570)<=x"ffdd";
m(1571)<=x"bff7";
m(1572)<=x"97ff";
m(1573)<=x"f9bf";
m(1574)<=x"ff3b";
m(1575)<=x"ffff";
m(1576)<=x"ffff";
m(1577)<=x"ffff";
m(1578)<=x"ff68";
m(1579)<=x"0000";
m(1580)<=x"0000";
m(1600)<=x"0000";
m(1601)<=x"0001";
m(1602)<=x"ffa3";
m(1603)<=x"fdaf";
m(1604)<=x"ffff";
m(1605)<=x"ffff";
m(1606)<=x"e9ef";
m(1607)<=x"ffff";
m(1608)<=x"ffff";
m(1609)<=x"ffff";
m(1610)<=x"fff8";
m(1611)<=x"0000";
m(1612)<=x"0000";
m(1632)<=x"0000";
m(1633)<=x"0007";
m(1634)<=x"febe";
m(1635)<=x"a7fd";
m(1636)<=x"bfff";
m(1637)<=x"7edd";
m(1638)<=x"bf77";
m(1639)<=x"ffff";
m(1640)<=x"ffff";
m(1641)<=x"ffff";
m(1642)<=x"ff85";
m(1643)<=x"0000";
m(1644)<=x"0000";
m(1664)<=x"0000";
m(1665)<=x"000f";
m(1666)<=x"7e5e";
m(1667)<=x"9bff";
m(1668)<=x"6fff";
m(1669)<=x"dfde";
m(1670)<=x"3cdd";
m(1671)<=x"ffff";
m(1672)<=x"ffff";
m(1673)<=x"ffff";
m(1674)<=x"ff80";
m(1675)<=x"0000";
m(1676)<=x"0000";
m(1696)<=x"0000";
m(1697)<=x"0035";
m(1698)<=x"d7e3";
m(1699)<=x"ffd4";
m(1700)<=x"7dff";
m(1701)<=x"ff7e";
m(1702)<=x"e7bb";
m(1703)<=x"ffff";
m(1704)<=x"ffff";
m(1705)<=x"ffff";
m(1706)<=x"ffe0";
m(1707)<=x"0000";
m(1708)<=x"0000";
m(1728)<=x"0000";
m(1729)<=x"0038";
m(1730)<=x"59a9";
m(1731)<=x"9dff";
m(1732)<=x"bfff";
m(1733)<=x"fff5";
m(1734)<=x"6db5";
m(1735)<=x"ffff";
m(1736)<=x"ffff";
m(1737)<=x"ffff";
m(1738)<=x"ffe6";
m(1739)<=x"0000";
m(1740)<=x"0000";
m(1760)<=x"0000";
m(1761)<=x"0009";
m(1762)<=x"3556";
m(1763)<=x"737b";
m(1764)<=x"ebff";
m(1765)<=x"ffee";
m(1766)<=x"d72f";
m(1767)<=x"fdff";
m(1768)<=x"ffff";
m(1769)<=x"ffff";
m(1770)<=x"fff0";
m(1771)<=x"0000";
m(1772)<=x"0000";
m(1792)<=x"0000";
m(1793)<=x"0018";
m(1794)<=x"355d";
m(1795)<=x"a6dc";
m(1796)<=x"fef7";
m(1797)<=x"fb77";
m(1798)<=x"6d5b";
m(1799)<=x"bfdf";
m(1800)<=x"efff";
m(1801)<=x"ffff";
m(1802)<=x"ff98";
m(1803)<=x"0000";
m(1804)<=x"0000";
m(1824)<=x"0000";
m(1825)<=x"0009";
m(1826)<=x"8ba6";
m(1827)<=x"59ab";
m(1828)<=x"cfed";
m(1829)<=x"ffec";
m(1830)<=x"66be";
m(1831)<=x"fbff";
m(1832)<=x"ffff";
m(1833)<=x"ffff";
m(1834)<=x"fff8";
m(1835)<=x"0000";
m(1836)<=x"0000";
m(1856)<=x"0000";
m(1857)<=x"0010";
m(1858)<=x"6f91";
m(1859)<=x"b656";
m(1860)<=x"76ff";
m(1861)<=x"fdff";
m(1862)<=x"f5db";
m(1863)<=x"d7bf";
m(1864)<=x"ffff";
m(1865)<=x"ffff";
m(1866)<=x"fffe";
m(1867)<=x"0000";
m(1868)<=x"0000";
m(1888)<=x"0000";
m(1889)<=x"0002";
m(1890)<=x"bc6d";
m(1891)<=x"eda9";
m(1892)<=x"5fd6";
m(1893)<=x"dff6";
m(1894)<=x"9d7f";
m(1895)<=x"bffd";
m(1896)<=x"ffff";
m(1897)<=x"ffff";
m(1898)<=x"fff9";
m(1899)<=x"0000";
m(1900)<=x"0000";
m(1920)<=x"0000";
m(1921)<=x"0001";
m(1922)<=x"afd6";
m(1923)<=x"6d49";
m(1924)<=x"effe";
m(1925)<=x"7fe7";
m(1926)<=x"9e67";
m(1927)<=x"ff5b";
m(1928)<=x"f7ff";
m(1929)<=x"ffff";
m(1930)<=x"fffc";
m(1931)<=x"0000";
m(1932)<=x"0000";
m(1952)<=x"0000";
m(1953)<=x"001f";
m(1954)<=x"fda9";
m(1955)<=x"1225";
m(1956)<=x"162b";
m(1957)<=x"efbd";
m(1958)<=x"ebff";
m(1959)<=x"b7ff";
m(1960)<=x"bfff";
m(1961)<=x"ffff";
m(1962)<=x"ffff";
m(1963)<=x"0000";
m(1964)<=x"0000";
m(1984)<=x"0000";
m(1985)<=x"001f";
m(1986)<=x"f552";
m(1987)<=x"bbc5";
m(1988)<=x"aabe";
m(1989)<=x"b7fe";
m(1990)<=x"bedf";
m(1991)<=x"5ebe";
m(1992)<=x"fdff";
m(1993)<=x"ffff";
m(1994)<=x"ffff";
m(1995)<=x"8000";
m(1996)<=x"0000";
m(2016)<=x"0000";
m(2017)<=x"003f";
m(2018)<=x"fea9";
m(2019)<=x"441a";
m(2020)<=x"5551";
m(2021)<=x"bfe7";
m(2022)<=x"f7ff";
m(2023)<=x"ffdb";
m(2024)<=x"db7f";
m(2025)<=x"ffff";
m(2026)<=x"fffb";
m(2027)<=x"8000";
m(2028)<=x"0000";
m(2048)<=x"0000";
m(2049)<=x"00ff";
m(2050)<=x"f67a";
m(2051)<=x"e596";
m(2052)<=x"9aad";
m(2053)<=x"dbff";
m(2054)<=x"dfff";
m(2055)<=x"ffff";
m(2056)<=x"ffff";
m(2057)<=x"ffff";
m(2058)<=x"fffb";
m(2059)<=x"4000";
m(2060)<=x"0000";
m(2080)<=x"0000";
m(2081)<=x"00ff";
m(2082)<=x"fdc5";
m(2083)<=x"1400";
m(2084)<=x"6596";
m(2085)<=x"7f9e";
m(2086)<=x"7fff";
m(2087)<=x"ffff";
m(2088)<=x"ffff";
m(2089)<=x"ffff";
m(2090)<=x"ffff";
m(2091)<=x"4000";
m(2092)<=x"0000";
m(2112)<=x"0000";
m(2113)<=x"01ff";
m(2114)<=x"8562";
m(2115)<=x"0029";
m(2116)<=x"812a";
m(2117)<=x"b6ff";
m(2118)<=x"feff";
m(2119)<=x"ffff";
m(2120)<=x"ffff";
m(2121)<=x"ffff";
m(2122)<=x"fffe";
m(2123)<=x"2000";
m(2124)<=x"0000";
m(2144)<=x"0000";
m(2145)<=x"03ff";
m(2146)<=x"ffa4";
m(2147)<=x"1606";
m(2148)<=x"5a5d";
m(2149)<=x"af7b";
m(2150)<=x"ffff";
m(2151)<=x"ffff";
m(2152)<=x"ffff";
m(2153)<=x"ffff";
m(2154)<=x"fffa";
m(2155)<=x"5000";
m(2156)<=x"0000";
m(2176)<=x"0000";
m(2177)<=x"07fe";
m(2178)<=x"ffa0";
m(2179)<=x"a4a4";
m(2180)<=x"8a43";
m(2181)<=x"ddff";
m(2182)<=x"ffff";
m(2183)<=x"ffff";
m(2184)<=x"ffff";
m(2185)<=x"ffff";
m(2186)<=x"fffc";
m(2187)<=x"0800";
m(2188)<=x"0000";
m(2208)<=x"0000";
m(2209)<=x"03ff";
m(2210)<=x"ba5a";
m(2211)<=x"0809";
m(2212)<=x"e4be";
m(2213)<=x"bfff";
m(2214)<=x"ffff";
m(2215)<=x"ffff";
m(2216)<=x"ffff";
m(2217)<=x"ffff";
m(2218)<=x"fff9";
m(2219)<=x"0000";
m(2220)<=x"0000";
m(2240)<=x"0000";
m(2241)<=x"07ff";
m(2242)<=x"dde6";
m(2243)<=x"2022";
m(2244)<=x"1d1f";
m(2245)<=x"f7f7";
m(2246)<=x"fdff";
m(2247)<=x"ffff";
m(2248)<=x"ffff";
m(2249)<=x"ffff";
m(2250)<=x"fffe";
m(2251)<=x"4200";
m(2252)<=x"0000";
m(2272)<=x"0000";
m(2273)<=x"07f7";
m(2274)<=x"5724";
m(2275)<=x"e427";
m(2276)<=x"e262";
m(2277)<=x"bfff";
m(2278)<=x"ffff";
m(2279)<=x"ffff";
m(2280)<=x"ffff";
m(2281)<=x"ffff";
m(2282)<=x"fffc";
m(2283)<=x"0800";
m(2284)<=x"0000";
m(2304)<=x"0000";
m(2305)<=x"01de";
m(2306)<=x"edd6";
m(2307)<=x"080d";
m(2308)<=x"696e";
m(2309)<=x"bfff";
m(2310)<=x"ffff";
m(2311)<=x"ffff";
m(2312)<=x"ffff";
m(2313)<=x"ffff";
m(2314)<=x"ffff";
m(2315)<=x"0000";
m(2316)<=x"0000";
m(2336)<=x"0000";
m(2337)<=x"01aa";
m(2338)<=x"996a";
m(2339)<=x"4126";
m(2340)<=x"829b";
m(2341)<=x"b7ff";
m(2342)<=x"ffff";
m(2343)<=x"ffff";
m(2344)<=x"ffff";
m(2345)<=x"ffff";
m(2346)<=x"ffff";
m(2347)<=x"0000";
m(2348)<=x"0000";
m(2368)<=x"0000";
m(2369)<=x"01e7";
m(2370)<=x"de94";
m(2371)<=x"3051";
m(2372)<=x"154e";
m(2373)<=x"ffff";
m(2374)<=x"ffff";
m(2375)<=x"ffff";
m(2376)<=x"ffff";
m(2377)<=x"ffff";
m(2378)<=x"ffff";
m(2379)<=x"0800";
m(2380)<=x"0000";
m(2400)<=x"0000";
m(2401)<=x"01c9";
m(2402)<=x"6229";
m(2403)<=x"8424";
m(2404)<=x"5ab3";
m(2405)<=x"efff";
m(2406)<=x"ffff";
m(2407)<=x"ffff";
m(2408)<=x"ffff";
m(2409)<=x"ffff";
m(2410)<=x"ffff";
m(2411)<=x"e000";
m(2412)<=x"0000";
m(2432)<=x"0000";
m(2433)<=x"01d5";
m(2434)<=x"5999";
m(2435)<=x"2c40";
m(2436)<=x"abdf";
m(2437)<=x"dfff";
m(2438)<=x"ffff";
m(2439)<=x"ffff";
m(2440)<=x"ffff";
m(2441)<=x"ffdf";
m(2442)<=x"ffff";
m(2443)<=x"f000";
m(2444)<=x"0000";
m(2464)<=x"0000";
m(2465)<=x"03f2";
m(2466)<=x"a562";
m(2467)<=x"4003";
m(2468)<=x"143b";
m(2469)<=x"ffff";
m(2470)<=x"ffff";
m(2471)<=x"ffff";
m(2472)<=x"ffff";
m(2473)<=x"ffff";
m(2474)<=x"ffff";
m(2475)<=x"f000";
m(2476)<=x"0000";
m(2496)<=x"0000";
m(2497)<=x"03f9";
m(2498)<=x"52a4";
m(2499)<=x"d808";
m(2500)<=x"32a8";
m(2501)<=x"57ff";
m(2502)<=x"ffff";
m(2503)<=x"ffff";
m(2504)<=x"ffff";
m(2505)<=x"ffff";
m(2506)<=x"ffff";
m(2507)<=x"fc00";
m(2508)<=x"0000";
m(2528)<=x"0000";
m(2529)<=x"01fe";
m(2530)<=x"9d87";
m(2531)<=x"2209";
m(2532)<=x"c895";
m(2533)<=x"ffff";
m(2534)<=x"ffff";
m(2535)<=x"ffff";
m(2536)<=x"ffff";
m(2537)<=x"ffff";
m(2538)<=x"ffff";
m(2539)<=x"fc00";
m(2540)<=x"0000";
m(2560)<=x"0000";
m(2561)<=x"03f5";
m(2562)<=x"5a64";
m(2563)<=x"2818";
m(2564)<=x"5136";
m(2565)<=x"ffff";
m(2566)<=x"ffff";
m(2567)<=x"ffff";
m(2568)<=x"ffff";
m(2569)<=x"ffef";
m(2570)<=x"ffff";
m(2571)<=x"ff00";
m(2572)<=x"0000";
m(2592)<=x"0000";
m(2593)<=x"03fe";
m(2594)<=x"8169";
m(2595)<=x"9002";
m(2596)<=x"01e7";
m(2597)<=x"ffff";
m(2598)<=x"7fff";
m(2599)<=x"ffff";
m(2600)<=x"ffff";
m(2601)<=x"ffff";
m(2602)<=x"ffff";
m(2603)<=x"fe00";
m(2604)<=x"0000";
m(2624)<=x"0000";
m(2625)<=x"07f6";
m(2626)<=x"a5d4";
m(2627)<=x"6008";
m(2628)<=x"063d";
m(2629)<=x"ffbc";
m(2630)<=x"ffbf";
m(2631)<=x"ffff";
m(2632)<=x"ffff";
m(2633)<=x"ffff";
m(2634)<=x"ffff";
m(2635)<=x"ff00";
m(2636)<=x"0000";
m(2656)<=x"0000";
m(2657)<=x"0fff";
m(2658)<=x"5b00";
m(2659)<=x"4090";
m(2660)<=x"2486";
m(2661)<=x"42d7";
m(2662)<=x"2a7d";
m(2663)<=x"ffff";
m(2664)<=x"ffff";
m(2665)<=x"ffff";
m(2666)<=x"ffff";
m(2667)<=x"fe00";
m(2668)<=x"0000";
m(2688)<=x"0000";
m(2689)<=x"1fff";
m(2690)<=x"e401";
m(2691)<=x"8000";
m(2692)<=x"6140";
m(2693)<=x"ffff";
m(2694)<=x"ff89";
m(2695)<=x"d7ff";
m(2696)<=x"ffff";
m(2697)<=x"ffff";
m(2698)<=x"ffff";
m(2699)<=x"ff00";
m(2700)<=x"0000";
m(2720)<=x"0000";
m(2721)<=x"0fef";
m(2722)<=x"62a4";
m(2723)<=x"4101";
m(2724)<=x"841f";
m(2725)<=x"ffff";
m(2726)<=x"ffff";
m(2727)<=x"ffff";
m(2728)<=x"ffff";
m(2729)<=x"fff7";
m(2730)<=x"ffff";
m(2731)<=x"ff00";
m(2732)<=x"0000";
m(2752)<=x"0000";
m(2753)<=x"1fd2";
m(2754)<=x"ba16";
m(2755)<=x"2003";
m(2756)<=x"0147";
m(2757)<=x"ffff";
m(2758)<=x"ffff";
m(2759)<=x"ffff";
m(2760)<=x"ffff";
m(2761)<=x"ffff";
m(2762)<=x"ffff";
m(2763)<=x"fe00";
m(2764)<=x"0000";
m(2784)<=x"0000";
m(2785)<=x"1f7f";
m(2786)<=x"e951";
m(2787)<=x"4418";
m(2788)<=x"6ab7";
m(2789)<=x"ffff";
m(2790)<=x"ffff";
m(2791)<=x"ffff";
m(2792)<=x"ffff";
m(2793)<=x"ff77";
m(2794)<=x"ffff";
m(2795)<=x"ff00";
m(2796)<=x"0000";
m(2816)<=x"0000";
m(2817)<=x"0fab";
m(2818)<=x"9cac";
m(2819)<=x"8018";
m(2820)<=x"22b7";
m(2821)<=x"eddf";
m(2822)<=x"ffff";
m(2823)<=x"ffff";
m(2824)<=x"ffff";
m(2825)<=x"ffff";
m(2826)<=x"ffff";
m(2827)<=x"fc00";
m(2828)<=x"0000";
m(2848)<=x"0000";
m(2849)<=x"2f7e";
m(2850)<=x"e392";
m(2851)<=x"1823";
m(2852)<=x"4808";
m(2853)<=x"5afd";
m(2854)<=x"ffff";
m(2855)<=x"ffff";
m(2856)<=x"ffff";
m(2857)<=x"ffef";
m(2858)<=x"ffff";
m(2859)<=x"f800";
m(2860)<=x"0000";
m(2880)<=x"0000";
m(2881)<=x"1ef7";
m(2882)<=x"7a41";
m(2883)<=x"a000";
m(2884)<=x"0000";
m(2885)<=x"ffe6";
m(2886)<=x"d7ff";
m(2887)<=x"ffff";
m(2888)<=x"ffff";
m(2889)<=x"fea7";
m(2890)<=x"ffff";
m(2891)<=x"f800";
m(2892)<=x"0000";
m(2912)<=x"0000";
m(2913)<=x"7fd9";
m(2914)<=x"9584";
m(2915)<=x"00a4";
m(2916)<=x"15bf";
m(2917)<=x"ffff";
m(2918)<=x"a4bb";
m(2919)<=x"ffff";
m(2920)<=x"ffff";
m(2921)<=x"ffff";
m(2922)<=x"ffff";
m(2923)<=x"f800";
m(2924)<=x"0000";
m(2944)<=x"0000";
m(2945)<=x"dfeb";
m(2946)<=x"e481";
m(2947)<=x"0018";
m(2948)<=x"b26b";
m(2949)<=x"bfff";
m(2950)<=x"ffab";
m(2951)<=x"1dff";
m(2952)<=x"ffff";
m(2953)<=x"ffff";
m(2954)<=x"ffff";
m(2955)<=x"fe00";
m(2956)<=x"0000";
m(2976)<=x"0000";
m(2977)<=x"2f7a";
m(2978)<=x"9928";
m(2979)<=x"2801";
m(2980)<=x"e809";
m(2981)<=x"ffff";
m(2982)<=x"ffff";
m(2983)<=x"deff";
m(2984)<=x"ffff";
m(2985)<=x"f9f7";
m(2986)<=x"ffff";
m(2987)<=x"f800";
m(2988)<=x"0000";
m(3008)<=x"0000";
m(3009)<=x"3bd6";
m(3010)<=x"a580";
m(3011)<=x"a003";
m(3012)<=x"41db";
m(3013)<=x"2fdb";
m(3014)<=x"ffff";
m(3015)<=x"ffff";
m(3016)<=x"ffff";
m(3017)<=x"efff";
m(3018)<=x"ffff";
m(3019)<=x"f800";
m(3020)<=x"0000";
m(3040)<=x"0000";
m(3041)<=x"3eef";
m(3042)<=x"5ab2";
m(3043)<=x"0214";
m(3044)<=x"1626";
m(3045)<=x"f56e";
m(3046)<=x"9dff";
m(3047)<=x"ffff";
m(3048)<=x"ffff";
m(3049)<=x"ff7f";
m(3050)<=x"ffff";
m(3051)<=x"ff00";
m(3052)<=x"0000";
m(3072)<=x"0000";
m(3073)<=x"2f75";
m(3074)<=x"3625";
m(3075)<=x"1024";
m(3076)<=x"051b";
m(3077)<=x"fffe";
m(3078)<=x"ae7f";
m(3079)<=x"7fff";
m(3080)<=x"ffff";
m(3081)<=x"ffff";
m(3082)<=x"ffff";
m(3083)<=x"ff80";
m(3084)<=x"0000";
m(3104)<=x"0000";
m(3105)<=x"39aa";
m(3106)<=x"81a0";
m(3107)<=x"0211";
m(3108)<=x"3855";
m(3109)<=x"bffb";
m(3110)<=x"5bdf";
m(3111)<=x"fbff";
m(3112)<=x"ffff";
m(3113)<=x"ff6f";
m(3114)<=x"ffff";
m(3115)<=x"ff80";
m(3116)<=x"0000";
m(3136)<=x"0000";
m(3137)<=x"29df";
m(3138)<=x"e244";
m(3139)<=x"8000";
m(3140)<=x"8086";
m(3141)<=x"7ffe";
m(3142)<=x"dbff";
m(3143)<=x"ffff";
m(3144)<=x"ffff";
m(3145)<=x"ff7d";
m(3146)<=x"ffff";
m(3147)<=x"ffc0";
m(3148)<=x"0000";
m(3168)<=x"0000";
m(3169)<=x"1efe";
m(3170)<=x"4924";
m(3171)<=x"103a";
m(3172)<=x"a180";
m(3173)<=x"0def";
m(3174)<=x"ae7d";
m(3175)<=x"dffb";
m(3176)<=x"ffff";
m(3177)<=x"ffaf";
m(3178)<=x"ffff";
m(3179)<=x"ffc0";
m(3180)<=x"0000";
m(3200)<=x"0000";
m(3201)<=x"0356";
m(3202)<=x"b291";
m(3203)<=x"0408";
m(3204)<=x"043a";
m(3205)<=x"ef6e";
m(3206)<=x"a2ff";
m(3207)<=x"affa";
m(3208)<=x"ffff";
m(3209)<=x"ffbf";
m(3210)<=x"ffff";
m(3211)<=x"fff0";
m(3212)<=x"0000";
m(3232)<=x"0000";
m(3233)<=x"007f";
m(3234)<=x"4d90";
m(3235)<=x"4053";
m(3236)<=x"17df";
m(3237)<=x"ffff";
m(3238)<=x"5553";
m(3239)<=x"f7ff";
m(3240)<=x"ffff";
m(3241)<=x"fdbf";
m(3242)<=x"ffff";
m(3243)<=x"fff0";
m(3244)<=x"0000";
m(3264)<=x"0000";
m(3265)<=x"0057";
m(3266)<=x"e040";
m(3267)<=x"0020";
m(3268)<=x"bf79";
m(3269)<=x"ffff";
m(3270)<=x"c6ad";
m(3271)<=x"ffff";
m(3272)<=x"ffff";
m(3273)<=x"ffff";
m(3274)<=x"ffff";
m(3275)<=x"fff0";
m(3276)<=x"0000";
m(3296)<=x"0000";
m(3297)<=x"0224";
m(3298)<=x"5588";
m(3299)<=x"6004";
m(3300)<=x"14df";
m(3301)<=x"ffff";
m(3302)<=x"fb5b";
m(3303)<=x"efff";
m(3304)<=x"ffff";
m(3305)<=x"fb7f";
m(3306)<=x"ffff";
m(3307)<=x"fff0";
m(3308)<=x"0000";
m(3328)<=x"0000";
m(3329)<=x"0021";
m(3330)<=x"2801";
m(3331)<=x"0019";
m(3332)<=x"b5d7";
m(3333)<=x"03ff";
m(3334)<=x"ffd4";
m(3335)<=x"f7ff";
m(3336)<=x"ffff";
m(3337)<=x"e7bf";
m(3338)<=x"ffff";
m(3339)<=x"fffc";
m(3340)<=x"0000";
m(3360)<=x"0000";
m(3361)<=x"0046";
m(3362)<=x"2644";
m(3363)<=x"0102";
m(3364)<=x"6011";
m(3365)<=x"7eff";
m(3366)<=x"ff9f";
m(3367)<=x"4fff";
m(3368)<=x"ffff";
m(3369)<=x"fdff";
m(3370)<=x"ffff";
m(3371)<=x"fffc";
m(3372)<=x"0000";
m(3392)<=x"0000";
m(3393)<=x"004a";
m(3394)<=x"6498";
m(3395)<=x"0009";
m(3396)<=x"b000";
m(3397)<=x"2aff";
m(3398)<=x"fffb";
m(3399)<=x"ffff";
m(3400)<=x"ffff";
m(3401)<=x"ff7f";
m(3402)<=x"ffff";
m(3403)<=x"ffbe";
m(3404)<=x"0000";
m(3424)<=x"0000";
m(3425)<=x"0015";
m(3426)<=x"db90";
m(3427)<=x"8012";
m(3428)<=x"4804";
m(3429)<=x"5fff";
m(3430)<=x"ffff";
m(3431)<=x"bfff";
m(3432)<=x"ffff";
m(3433)<=x"fdff";
m(3434)<=x"ffff";
m(3435)<=x"ff1e";
m(3436)<=x"0000";
m(3456)<=x"0000";
m(3457)<=x"0062";
m(3458)<=x"7711";
m(3459)<=x"0015";
m(3460)<=x"4000";
m(3461)<=x"13ff";
m(3462)<=x"ffff";
m(3463)<=x"e7ff";
m(3464)<=x"ffff";
m(3465)<=x"faff";
m(3466)<=x"ffff";
m(3467)<=x"ff0c";
m(3468)<=x"0000";
m(3488)<=x"0000";
m(3489)<=x"0002";
m(3490)<=x"dc48";
m(3491)<=x"064b";
m(3492)<=x"8000";
m(3493)<=x"00df";
m(3494)<=x"ffff";
m(3495)<=x"ffcf";
m(3496)<=x"ffff";
m(3497)<=x"ffff";
m(3498)<=x"ffff";
m(3499)<=x"ffbc";
m(3500)<=x"0000";
m(3520)<=x"0000";
m(3521)<=x"0048";
m(3522)<=x"3d10";
m(3523)<=x"022f";
m(3524)<=x"0000";
m(3525)<=x"02ff";
m(3526)<=x"ff7f";
m(3527)<=x"ffdf";
m(3528)<=x"ffff";
m(3529)<=x"f7ff";
m(3530)<=x"ffff";
m(3531)<=x"ffae";
m(3532)<=x"0000";
m(3552)<=x"0000";
m(3553)<=x"0220";
m(3554)<=x"0ac8";
m(3555)<=x"0018";
m(3556)<=x"0000";
m(3557)<=x"041f";
m(3558)<=x"ffff";
m(3559)<=x"6bb3";
m(3560)<=x"ffff";
m(3561)<=x"da5f";
m(3562)<=x"ffff";
m(3563)<=x"fff8";
m(3564)<=x"0000";
m(3584)<=x"0000";
m(3585)<=x"0462";
m(3586)<=x"0f00";
m(3587)<=x"0496";
m(3588)<=x"0000";
m(3589)<=x"001d";
m(3590)<=x"ffbf";
m(3591)<=x"ed06";
m(3592)<=x"ffff";
m(3593)<=x"f6ff";
m(3594)<=x"ffff";
m(3595)<=x"ffdc";
m(3596)<=x"0000";
m(3616)<=x"0000";
m(3617)<=x"0008";
m(3618)<=x"1020";
m(3619)<=x"210d";
m(3620)<=x"8800";
m(3621)<=x"0046";
m(3622)<=x"fffd";
m(3623)<=x"a600";
m(3624)<=x"097f";
m(3625)<=x"ff5f";
m(3626)<=x"ffff";
m(3627)<=x"7fdc";
m(3628)<=x"0000";
m(3648)<=x"0000";
m(3649)<=x"001a";
m(3650)<=x"0380";
m(3651)<=x"2010";
m(3652)<=x"8000";
m(3653)<=x"0095";
m(3654)<=x"7ffb";
m(3655)<=x"4000";
m(3656)<=x"017f";
m(3657)<=x"fdef";
m(3658)<=x"ffff";
m(3659)<=x"fffc";
m(3660)<=x"0000";
m(3680)<=x"0000";
m(3681)<=x"00e4";
m(3682)<=x"0000";
m(3683)<=x"0565";
m(3684)<=x"1000";
m(3685)<=x"0004";
m(3686)<=x"69dd";
m(3687)<=x"a000";
m(3688)<=x"029f";
m(3689)<=x"ffbf";
m(3690)<=x"ffff";
m(3691)<=x"fffc";
m(3692)<=x"0000";
m(3712)<=x"0000";
m(3713)<=x"0092";
m(3714)<=x"0000";
m(3715)<=x"4208";
m(3716)<=x"0000";
m(3717)<=x"0001";
m(3718)<=x"37ed";
m(3719)<=x"0800";
m(3720)<=x"001f";
m(3721)<=x"ffdf";
m(3722)<=x"ffff";
m(3723)<=x"ebfe";
m(3724)<=x"0000";
m(3744)<=x"0000";
m(3745)<=x"00e8";
m(3746)<=x"0020";
m(3747)<=x"1450";
m(3748)<=x"6000";
m(3749)<=x"0000";
m(3750)<=x"4d76";
m(3751)<=x"8000";
m(3752)<=x"0057";
m(3753)<=x"fe9f";
m(3754)<=x"fdff";
m(3755)<=x"fffc";
m(3756)<=x"0000";
m(3776)<=x"0000";
m(3777)<=x"00c6";
m(3778)<=x"0080";
m(3779)<=x"8288";
m(3780)<=x"4000";
m(3781)<=x"0001";
m(3782)<=x"2969";
m(3783)<=x"0000";
m(3784)<=x"000f";
m(3785)<=x"ffdf";
m(3786)<=x"ffff";
m(3787)<=x"fffc";
m(3788)<=x"0000";
m(3808)<=x"0000";
m(3809)<=x"01a9";
m(3810)<=x"0000";
m(3811)<=x"1820";
m(3812)<=x"0010";
m(3813)<=x"0000";
m(3814)<=x"26da";
m(3815)<=x"0000";
m(3816)<=x"0011";
m(3817)<=x"ffbf";
m(3818)<=x"ffff";
m(3819)<=x"b9fc";
m(3820)<=x"0000";
m(3840)<=x"0000";
m(3841)<=x"03e4";
m(3842)<=x"0020";
m(3843)<=x"0490";
m(3844)<=x"0000";
m(3845)<=x"0000";
m(3846)<=x"4a68";
m(3847)<=x"0000";
m(3848)<=x"0001";
m(3849)<=x"ff7f";
m(3850)<=x"ffff";
m(3851)<=x"edfe";
m(3852)<=x"0000";
m(3872)<=x"0000";
m(3873)<=x"0399";
m(3874)<=x"4000";
m(3875)<=x"aa00";
m(3876)<=x"0000";
m(3877)<=x"0000";
m(3878)<=x"1596";
m(3879)<=x"0000";
m(3880)<=x"0000";
m(3881)<=x"ffdf";
m(3882)<=x"e3fa";
m(3883)<=x"ba5c";
m(3884)<=x"0000";
m(3904)<=x"0000";
m(3905)<=x"0245";
m(3906)<=x"8001";
m(3907)<=x"2483";
m(3908)<=x"8000";
m(3909)<=x"0000";
m(3910)<=x"07dc";
m(3911)<=x"0000";
m(3912)<=x"0001";
m(3913)<=x"ffbf";
m(3914)<=x"f7ff";
m(3915)<=x"e5f8";
m(3916)<=x"0000";
m(3936)<=x"0000";
m(3937)<=x"03aa";
m(3938)<=x"0020";
m(3939)<=x"1220";
m(3940)<=x"8000";
m(3941)<=x"0000";
m(3942)<=x"2260";
m(3943)<=x"0000";
m(3944)<=x"0000";
m(3945)<=x"ffff";
m(3946)<=x"fa6f";
m(3947)<=x"fbfc";
m(3948)<=x"0000";
m(3968)<=x"0000";
m(3969)<=x"04d3";
m(3970)<=x"0000";
m(3971)<=x"1848";
m(3972)<=x"0000";
m(3973)<=x"0000";
m(3974)<=x"0bf0";
m(3975)<=x"0000";
m(3976)<=x"0700";
m(3977)<=x"5fef";
m(3978)<=x"f7ad";
m(3979)<=x"ad7a";
m(3980)<=x"0000";
m(4000)<=x"0000";
m(4001)<=x"054a";
m(4002)<=x"e008";
m(4003)<=x"4512";
m(4004)<=x"0000";
m(4005)<=x"0000";
m(4006)<=x"55e0";
m(4007)<=x"0000";
m(4008)<=x"0006";
m(4009)<=x"bdff";
m(4010)<=x"fff7";
m(4011)<=x"d3fd";
m(4012)<=x"0000";
m(4032)<=x"0000";
m(4033)<=x"05bd";
m(4034)<=x"8000";
m(4035)<=x"a944";
m(4036)<=x"0000";
m(4037)<=x"1001";
m(4038)<=x"4bf0";
m(4039)<=x"0000";
m(4040)<=x"0006";
m(4041)<=x"7bff";
m(4042)<=x"ffff";
m(4043)<=x"9dd8";
m(4044)<=x"0000";
m(4064)<=x"0000";
m(4065)<=x"024b";
m(4066)<=x"c000";
m(4067)<=x"8250";
m(4068)<=x"0000";
m(4069)<=x"0000";
m(4070)<=x"17f8";
m(4071)<=x"0000";
m(4072)<=x"0002";
m(4073)<=x"7fff";
m(4074)<=x"fffd";
m(4075)<=x"aafe";
m(4076)<=x"0000";
m(4096)<=x"0000";
m(4097)<=x"013b";
m(4098)<=x"a008";
m(4099)<=x"2508";
m(4100)<=x"0940";
m(4101)<=x"2188";
m(4102)<=x"9ffc";
m(4103)<=x"00c0";
m(4104)<=x"0002";
m(4105)<=x"3fff";
m(4106)<=x"ffff";
m(4107)<=x"2d7c";
m(4108)<=x"8000";
m(4128)<=x"0000";
m(4129)<=x"08ee";
m(4130)<=x"601a";
m(4131)<=x"a660";
m(4132)<=x"0190";
m(4133)<=x"0859";
m(4134)<=x"4ffe";
m(4135)<=x"0040";
m(4136)<=x"0803";
m(4137)<=x"9fff";
m(4138)<=x"ffbb";
m(4139)<=x"e7fa";
m(4140)<=x"0000";
m(4160)<=x"0000";
m(4161)<=x"01ee";
m(4162)<=x"e510";
m(4163)<=x"09c6";
m(4164)<=x"1166";
m(4165)<=x"19a4";
m(4166)<=x"affe";
m(4167)<=x"8080";
m(4168)<=x"1901";
m(4169)<=x"3fef";
m(4170)<=x"fefa";
m(4171)<=x"adfd";
m(4172)<=x"0000";
m(4192)<=x"0000";
m(4193)<=x"0335";
m(4194)<=x"603e";
m(4195)<=x"5220";
m(4196)<=x"483f";
m(4197)<=x"e401";
m(4198)<=x"5fff";
m(4199)<=x"3c60";
m(4200)<=x"1f09";
m(4201)<=x"bfff";
m(4202)<=x"dfef";
m(4203)<=x"d75e";
m(4204)<=x"2000";
m(4224)<=x"0000";
m(4225)<=x"0a58";
m(4226)<=x"7236";
m(4227)<=x"a800";
m(4228)<=x"900d";
m(4229)<=x"8045";
m(4230)<=x"5fff";
m(4231)<=x"39f1";
m(4232)<=x"ff8d";
m(4233)<=x"ffef";
m(4234)<=x"ffff";
m(4235)<=x"6dfc";
m(4236)<=x"0000";
m(4256)<=x"0000";
m(4257)<=x"017a";
m(4258)<=x"e0bd";
m(4259)<=x"93ba";
m(4260)<=x"2c00";
m(4261)<=x"021a";
m(4262)<=x"2fff";
m(4263)<=x"ec3f";
m(4264)<=x"fd87";
m(4265)<=x"fffc";
m(4266)<=x"bfff";
m(4267)<=x"d75f";
m(4268)<=x"8000";
m(4288)<=x"0000";
m(4289)<=x"01bb";
m(4290)<=x"7916";
m(4291)<=x"4a20";
m(4292)<=x"9400";
m(4293)<=x"0016";
m(4294)<=x"bfff";
m(4295)<=x"f205";
m(4296)<=x"7441";
m(4297)<=x"ffc5";
m(4298)<=x"7fff";
m(4299)<=x"cdfe";
m(4300)<=x"a000";
m(4320)<=x"0000";
m(4321)<=x"0962";
m(4322)<=x"d876";
m(4323)<=x"984b";
m(4324)<=x"2a40";
m(4325)<=x"082a";
m(4326)<=x"5fff";
m(4327)<=x"e400";
m(4328)<=x"02f2";
m(4329)<=x"fff0";
m(4330)<=x"bfff";
m(4331)<=x"bf9d";
m(4332)<=x"4000";
m(4352)<=x"0000";
m(4353)<=x"0129";
m(4354)<=x"5876";
m(4355)<=x"4e8b";
m(4356)<=x"aa02";
m(4357)<=x"40db";
m(4358)<=x"afff";
m(4359)<=x"fd80";
m(4360)<=x"27f7";
m(4361)<=x"fff0";
m(4362)<=x"7fdf";
m(4363)<=x"df5e";
m(4364)<=x"8000";
m(4384)<=x"0000";
m(4385)<=x"01b5";
m(4386)<=x"c8f7";
m(4387)<=x"3166";
m(4388)<=x"59ec";
m(4389)<=x"02a8";
m(4390)<=x"5fff";
m(4391)<=x"f828";
m(4392)<=x"8bff";
m(4393)<=x"ffe1";
m(4394)<=x"9fff";
m(4395)<=x"ff9e";
m(4396)<=x"4000";
m(4416)<=x"0000";
m(4417)<=x"0229";
m(4418)<=x"b567";
m(4419)<=x"94f6";
m(4420)<=x"745a";
m(4421)<=x"8866";
m(4422)<=x"7fff";
m(4423)<=x"f165";
m(4424)<=x"17ff";
m(4425)<=x"fff5";
m(4426)<=x"bfff";
m(4427)<=x"f6b7";
m(4428)<=x"2000";
m(4448)<=x"0000";
m(4449)<=x"0099";
m(4450)<=x"dc7d";
m(4451)<=x"6a0d";
m(4452)<=x"4b70";
m(4453)<=x"13bd";
m(4454)<=x"7fff";
m(4455)<=x"fe09";
m(4456)<=x"dfef";
m(4457)<=x"fff3";
m(4458)<=x"dfff";
m(4459)<=x"ff9e";
m(4460)<=x"8000";
m(4480)<=x"0000";
m(4481)<=x"0025";
m(4482)<=x"b4da";
m(4483)<=x"aba2";
m(4484)<=x"4624";
m(4485)<=x"2998";
m(4486)<=x"5fff";
m(4487)<=x"fd8f";
m(4488)<=x"ffff";
m(4489)<=x"fffa";
m(4490)<=x"7fff";
m(4491)<=x"ff92";
m(4492)<=x"0000";
m(4512)<=x"0000";
m(4513)<=x"021a";
m(4514)<=x"da7f";
m(4515)<=x"544f";
m(4516)<=x"bda1";
m(4517)<=x"476e";
m(4518)<=x"9fff";
m(4519)<=x"ff55";
m(4520)<=x"ffff";
m(4521)<=x"fff1";
m(4522)<=x"67ff";
m(4523)<=x"fffd";
m(4524)<=x"c000";
m(4544)<=x"0000";
m(4545)<=x"2296";
m(4546)<=x"b446";
m(4547)<=x"6a55";
m(4548)<=x"7655";
m(4549)<=x"deb5";
m(4550)<=x"9fff";
m(4551)<=x"ffc1";
m(4552)<=x"ffff";
m(4553)<=x"fff7";
m(4554)<=x"ffff";
m(4555)<=x"f7e6";
m(4556)<=x"8000";
m(4576)<=x"0000";
m(4577)<=x"0009";
m(4578)<=x"a3a7";
m(4579)<=x"94ad";
m(4580)<=x"c94a";
m(4581)<=x"295a";
m(4582)<=x"6fff";
m(4583)<=x"ff54";
m(4584)<=x"3fff";
m(4585)<=x"fff4";
m(4586)<=x"bfff";
m(4587)<=x"ffeb";
m(4588)<=x"0000";
m(4608)<=x"0000";
m(4609)<=x"00b1";
m(4610)<=x"f257";
m(4611)<=x"9957";
m(4612)<=x"cac2";
m(4613)<=x"5d5a";
m(4614)<=x"9fff";
m(4615)<=x"fff1";
m(4616)<=x"9dff";
m(4617)<=x"fffe";
m(4618)<=x"7fff";
m(4619)<=x"fff6";
m(4620)<=x"0000";
m(4640)<=x"0000";
m(4641)<=x"0109";
m(4642)<=x"2c21";
m(4643)<=x"a6aa";
m(4644)<=x"6819";
m(4645)<=x"b225";
m(4646)<=x"afff";
m(4647)<=x"fffd";
m(4648)<=x"ff7f";
m(4649)<=x"fff7";
m(4650)<=x"bfff";
m(4651)<=x"fffa";
m(4652)<=x"6000";
m(4672)<=x"0000";
m(4673)<=x"0015";
m(4674)<=x"e56b";
m(4675)<=x"d619";
m(4676)<=x"a299";
m(4677)<=x"a998";
m(4678)<=x"dfff";
m(4679)<=x"fffd";
m(4680)<=x"efff";
m(4681)<=x"fff2";
m(4682)<=x"bfff";
m(4683)<=x"ffba";
m(4684)<=x"0000";
m(4704)<=x"0000";
m(4705)<=x"0022";
m(4706)<=x"7207";
m(4707)<=x"4a64";
m(4708)<=x"5927";
m(4709)<=x"566a";
m(4710)<=x"2fff";
m(4711)<=x"fff6";
m(4712)<=x"5fff";
m(4713)<=x"ffff";
m(4714)<=x"ffff";
m(4715)<=x"fdfe";
m(4716)<=x"5000";
m(4736)<=x"0000";
m(4737)<=x"0021";
m(4738)<=x"b80b";
m(4739)<=x"958a";
m(4740)<=x"4696";
m(4741)<=x"dbd3";
m(4742)<=x"2fff";
m(4743)<=x"ffff";
m(4744)<=x"97ff";
m(4745)<=x"fffb";
m(4746)<=x"afff";
m(4747)<=x"fffc";
m(4748)<=x"8000";
m(4768)<=x"0000";
m(4769)<=x"0085";
m(4770)<=x"6197";
m(4771)<=x"e635";
m(4772)<=x"99aa";
m(4773)<=x"a6a8";
m(4774)<=x"bfff";
m(4775)<=x"ffff";
m(4776)<=x"eeff";
m(4777)<=x"fff3";
m(4778)<=x"ffff";
m(4779)<=x"fffe";
m(4780)<=x"0200";
m(4800)<=x"0000";
m(4801)<=x"008a";
m(4802)<=x"663b";
m(4803)<=x"cb66";
m(4804)<=x"6415";
m(4805)<=x"aee5";
m(4806)<=x"bfff";
m(4807)<=x"ffff";
m(4808)<=x"fa7f";
m(4809)<=x"ffff";
m(4810)<=x"ffff";
m(4811)<=x"ffea";
m(4812)<=x"0000";
m(4832)<=x"0000";
m(4833)<=x"0918";
m(4834)<=x"d907";
m(4835)<=x"b412";
m(4836)<=x"526a";
m(4837)<=x"5734";
m(4838)<=x"7fff";
m(4839)<=x"ffff";
m(4840)<=x"ffaf";
m(4841)<=x"ffff";
m(4842)<=x"efff";
m(4843)<=x"ffff";
m(4844)<=x"4000";
m(4864)<=x"0000";
m(4865)<=x"0299";
m(4866)<=x"ea0b";
m(4867)<=x"d6a4";
m(4868)<=x"b195";
m(4869)<=x"ed95";
m(4870)<=x"bfff";
m(4871)<=x"ffff";
m(4872)<=x"fcdf";
m(4873)<=x"fff7";
m(4874)<=x"efff";
m(4875)<=x"fff6";
m(4876)<=x"0000";
m(4896)<=x"0000";
m(4897)<=x"06e2";
m(4898)<=x"6111";
m(4899)<=x"ed89";
m(4900)<=x"052a";
m(4901)<=x"7ec2";
m(4902)<=x"5fff";
m(4903)<=x"ffff";
m(4904)<=x"a965";
m(4905)<=x"fff7";
m(4906)<=x"ffff";
m(4907)<=x"fffb";
m(4908)<=x"1000";
m(4928)<=x"0000";
m(4929)<=x"07ee";
m(4930)<=x"7111";
m(4931)<=x"f831";
m(4932)<=x"6c95";
m(4933)<=x"ea02";
m(4934)<=x"7fff";
m(4935)<=x"ffff";
m(4936)<=x"f6af";
m(4937)<=x"fff7";
m(4938)<=x"ffff";
m(4939)<=x"fff9";
m(4940)<=x"9000";
m(4960)<=x"0000";
m(4961)<=x"03c2";
m(4962)<=x"6201";
m(4963)<=x"ae8c";
m(4964)<=x"416b";
m(4965)<=x"be05";
m(4966)<=x"bfff";
m(4967)<=x"efff";
m(4968)<=x"fd37";
m(4969)<=x"ffff";
m(4970)<=x"ffff";
m(4971)<=x"ffd6";
m(4972)<=x"0000";
m(4992)<=x"0000";
m(4993)<=x"0306";
m(4994)<=x"6201";
m(4995)<=x"eb85";
m(4996)<=x"59aa";
m(4997)<=x"ac36";
m(4998)<=x"7fff";
m(4999)<=x"fbff";
m(5000)<=x"ffd7";
m(5001)<=x"ffff";
m(5002)<=x"ffff";
m(5003)<=x"ffdb";
m(5004)<=x"0000";
m(5024)<=x"0000";
m(5025)<=x"0604";
m(5026)<=x"c11c";
m(5027)<=x"f938";
m(5028)<=x"aa7b";
m(5029)<=x"f081";
m(5030)<=x"7fff";
m(5031)<=x"f7ff";
m(5032)<=x"fffe";
m(5033)<=x"fdff";
m(5034)<=x"ffff";
m(5035)<=x"fff9";
m(5036)<=x"0000";
m(5056)<=x"0000";
m(5057)<=x"000c";
m(5058)<=x"1099";
m(5059)<=x"dea7";
m(5060)<=x"5156";
m(5061)<=x"90a6";
m(5062)<=x"ffff";
m(5063)<=x"fbff";
m(5064)<=x"ff47";
m(5065)<=x"fbff";
m(5066)<=x"ffff";
m(5067)<=x"ffda";
m(5068)<=x"8000";
m(5088)<=x"0000";
m(5089)<=x"0411";
m(5090)<=x"9004";
m(5091)<=x"7b92";
m(5092)<=x"aedf";
m(5093)<=x"f431";
m(5094)<=x"7fff";
m(5095)<=x"f1ff";
m(5096)<=x"fffb";
m(5097)<=x"f5ff";
m(5098)<=x"ffff";
m(5099)<=x"fffd";
m(5100)<=x"0000";
m(5120)<=x"0000";
m(5121)<=x"0048";
m(5122)<=x"210c";
m(5123)<=x"fc95";
m(5124)<=x"adff";
m(5125)<=x"4052";
m(5126)<=x"7fff";
m(5127)<=x"fdff";
m(5128)<=x"ffef";
m(5129)<=x"f7ef";
m(5130)<=x"ffff";
m(5131)<=x"fff9";
m(5132)<=x"8000";
m(5152)<=x"0000";
m(5153)<=x"0004";
m(5154)<=x"56a8";
m(5155)<=x"77aa";
m(5156)<=x"9769";
m(5157)<=x"a4e1";
m(5158)<=x"bfff";
m(5159)<=x"f8ff";
m(5160)<=x"ffff";
m(5161)<=x"fcef";
m(5162)<=x"ffff";
m(5163)<=x"ffe1";
m(5164)<=x"8000";
m(5184)<=x"0000";
m(5185)<=x"0010";
m(5186)<=x"4591";
m(5187)<=x"6e95";
m(5188)<=x"5c7f";
m(5189)<=x"06a2";
m(5190)<=x"7fff";
m(5191)<=x"fa7f";
m(5192)<=x"ffff";
m(5193)<=x"e7ff";
m(5194)<=x"ffff";
m(5195)<=x"fff5";
m(5196)<=x"0000";
m(5216)<=x"0000";
m(5217)<=x"0008";
m(5218)<=x"1058";
m(5219)<=x"7b69";
m(5220)<=x"b7ec";
m(5221)<=x"0359";
m(5222)<=x"7fff";
m(5223)<=x"fc3f";
m(5224)<=x"ffff";
m(5225)<=x"e5ef";
m(5226)<=x"fdff";
m(5227)<=x"f7f0";
m(5228)<=x"8000";
m(5248)<=x"0000";
m(5249)<=x"0000";
m(5250)<=x"4000";
m(5251)<=x"6da5";
m(5252)<=x"aeda";
m(5253)<=x"0eca";
m(5254)<=x"57ff";
m(5255)<=x"fe3f";
m(5256)<=x"ffff";
m(5257)<=x"fcff";
m(5258)<=x"fddf";
m(5259)<=x"fff4";
m(5260)<=x"0000";
m(5280)<=x"0000";
m(5281)<=x"0020";
m(5282)<=x"1804";
m(5283)<=x"3a5a";
m(5284)<=x"537e";
m(5285)<=x"3a20";
m(5286)<=x"afff";
m(5287)<=x"ff8f";
m(5288)<=x"ffff";
m(5289)<=x"e3ff";
m(5290)<=x"ffff";
m(5291)<=x"ffc9";
m(5292)<=x"0000";
m(5312)<=x"0000";
m(5313)<=x"0000";
m(5314)<=x"0008";
m(5315)<=x"3b88";
m(5316)<=x"afb0";
m(5317)<=x"5620";
m(5318)<=x"55ff";
m(5319)<=x"ff97";
m(5320)<=x"ffff";
m(5321)<=x"c57f";
m(5322)<=x"fdff";
m(5323)<=x"fff9";
m(5324)<=x"8000";
m(5344)<=x"0000";
m(5345)<=x"0000";
m(5346)<=x"0000";
m(5347)<=x"1d6d";
m(5348)<=x"55e8";
m(5349)<=x"7d00";
m(5350)<=x"0bff";
m(5351)<=x"ffcb";
m(5352)<=x"ffff";
m(5353)<=x"cbff";
m(5354)<=x"ffff";
m(5355)<=x"ffd0";
m(5356)<=x"0000";
m(5376)<=x"0000";
m(5377)<=x"0000";
m(5378)<=x"0004";
m(5379)<=x"1eaa";
m(5380)<=x"ade8";
m(5381)<=x"7700";
m(5382)<=x"4bbf";
m(5383)<=x"ffe7";
m(5384)<=x"ffff";
m(5385)<=x"dbff";
m(5386)<=x"ffff";
m(5387)<=x"ffe9";
m(5388)<=x"0000";
m(5408)<=x"0000";
m(5409)<=x"0000";
m(5410)<=x"0000";
m(5411)<=x"1b95";
m(5412)<=x"7b51";
m(5413)<=x"ad80";
m(5414)<=x"00a6";
m(5415)<=x"7fe6";
m(5416)<=x"ffff";
m(5417)<=x"cfff";
m(5418)<=x"ffff";
m(5419)<=x"fff0";
m(5420)<=x"0000";
m(5440)<=x"0000";
m(5441)<=x"0000";
m(5442)<=x"0000";
m(5443)<=x"064a";
m(5444)<=x"9d81";
m(5445)<=x"9780";
m(5446)<=x"0064";
m(5447)<=x"fff5";
m(5448)<=x"ffff";
m(5449)<=x"bfff";
m(5450)<=x"ffff";
m(5451)<=x"dff0";
m(5452)<=x"0000";
m(5472)<=x"0000";
m(5473)<=x"0000";
m(5474)<=x"0000";
m(5475)<=x"0ea3";
m(5476)<=x"7a67";
m(5477)<=x"dc40";
m(5478)<=x"000b";
m(5479)<=x"fff3";
m(5480)<=x"ffff";
m(5481)<=x"ffff";
m(5482)<=x"ffff";
m(5483)<=x"fff0";
m(5484)<=x"0000";
m(5504)<=x"0000";
m(5505)<=x"0000";
m(5506)<=x"0000";
m(5507)<=x"0d4d";
m(5508)<=x"b5c6";
m(5509)<=x"57d0";
m(5510)<=x"000f";
m(5511)<=x"fff9";
m(5512)<=x"ffff";
m(5513)<=x"ffff";
m(5514)<=x"ffff";
m(5515)<=x"ffe0";
m(5516)<=x"0000";
m(5536)<=x"0000";
m(5537)<=x"0000";
m(5538)<=x"0000";
m(5539)<=x"06b0";
m(5540)<=x"ea1f";
m(5541)<=x"b666";
m(5542)<=x"001f";
m(5543)<=x"ffff";
m(5544)<=x"7fff";
m(5545)<=x"ffff";
m(5546)<=x"ffff";
m(5547)<=x"fff8";
m(5548)<=x"0000";
m(5568)<=x"0000";
m(5569)<=x"0000";
m(5570)<=x"0000";
m(5571)<=x"2223";
m(5572)<=x"95bb";
m(5573)<=x"21c8";
m(5574)<=x"007f";
m(5575)<=x"ffff";
m(5576)<=x"7fff";
m(5577)<=x"ffff";
m(5578)<=x"ffff";
m(5579)<=x"fff8";
m(5580)<=x"0000";
m(5600)<=x"0000";
m(5601)<=x"0000";
m(5602)<=x"0000";
m(5603)<=x"a58c";
m(5604)<=x"6a24";
m(5605)<=x"de16";
m(5606)<=x"007f";
m(5607)<=x"ffff";
m(5608)<=x"bfff";
m(5609)<=x"ffff";
m(5610)<=x"ffff";
m(5611)<=x"fffd";
m(5612)<=x"0000";
m(5632)<=x"0000";
m(5633)<=x"0000";
m(5634)<=x"0001";
m(5635)<=x"410d";
m(5636)<=x"caab";
m(5637)<=x"bce5";
m(5638)<=x"037f";
m(5639)<=x"ffff";
m(5640)<=x"bfff";
m(5641)<=x"ffff";
m(5642)<=x"ffdf";
m(5643)<=x"fefa";
m(5644)<=x"a000";
m(5664)<=x"0000";
m(5665)<=x"0000";
m(5666)<=x"0004";
m(5667)<=x"0252";
m(5668)<=x"59fd";
m(5669)<=x"d310";
m(5670)<=x"ba97";
m(5671)<=x"ffff";
m(5672)<=x"efff";
m(5673)<=x"ffff";
m(5674)<=x"fffd";
m(5675)<=x"ff7a";
m(5676)<=x"5000";
m(5696)<=x"0000";
m(5697)<=x"0000";
m(5698)<=x"0002";
m(5699)<=x"0220";
m(5700)<=x"807a";
m(5701)<=x"4529";
m(5702)<=x"58db";
m(5703)<=x"ffff";
m(5704)<=x"dfff";
m(5705)<=x"ffff";
m(5706)<=x"f7f7";
m(5707)<=x"fdf4";
m(5708)<=x"1c00";
m(5728)<=x"0000";
m(5729)<=x"0000";
m(5730)<=x"0004";
m(5731)<=x"0189";
m(5732)<=x"5740";
m(5733)<=x"92c5";
m(5734)<=x"bb3f";
m(5735)<=x"ffff";
m(5736)<=x"cfff";
m(5737)<=x"ffff";
m(5738)<=x"ffb6";
m(5739)<=x"ff91";
m(5740)<=x"81d4";
m(5760)<=x"0000";
m(5761)<=x"0000";
m(5762)<=x"0001";
m(5763)<=x"02a2";
m(5764)<=x"8691";
m(5765)<=x"1b1d";
m(5766)<=x"757d";
m(5767)<=x"ffff";
m(5768)<=x"dfff";
m(5769)<=x"ffff";
m(5770)<=x"fbfc";
m(5771)<=x"ff7c";
m(5772)<=x"8015";
m(5792)<=x"0000";
m(5793)<=x"0000";
m(5794)<=x"0008";
m(5795)<=x"0200";
m(5796)<=x"1299";
m(5797)<=x"8065";
m(5798)<=x"7b2f";
m(5799)<=x"ffff";
m(5800)<=x"e7ff";
m(5801)<=x"ffff";
m(5802)<=x"f7df";
m(5803)<=x"7ed8";
m(5804)<=x"2a67";
m(5824)<=x"0000";
m(5825)<=x"0000";
m(5826)<=x"0000";
m(5827)<=x"0302";
m(5828)<=x"6602";
m(5829)<=x"812a";
m(5830)<=x"73f7";
m(5831)<=x"ffff";
m(5832)<=x"ffff";
m(5833)<=x"ffff";
m(5834)<=x"f9ff";
m(5835)<=x"a71a";
m(5836)<=x"0152";
m(5856)<=x"0000";
m(5857)<=x"0000";
m(5858)<=x"0020";
m(5859)<=x"0310";
m(5860)<=x"0091";
m(5861)<=x"1043";
m(5862)<=x"dbb6";
m(5863)<=x"ffff";
m(5864)<=x"e7ff";
m(5865)<=x"ffff";
m(5866)<=x"fafe";
m(5867)<=x"ff4a";
m(5868)<=x"4809";
m(5888)<=x"0000";
m(5889)<=x"0000";
m(5890)<=x"0004";
m(5891)<=x"0708";
m(5892)<=x"1180";
m(5893)<=x"0046";
m(5894)<=x"e567";
m(5895)<=x"dfff";
m(5896)<=x"efff";
m(5897)<=x"ffff";
m(5898)<=x"0e7b";
m(5899)<=x"fe08";
m(5900)<=x"0220";
m(5920)<=x"0000";
m(5921)<=x"0000";
m(5922)<=x"0000";
m(5923)<=x"0780";
m(5924)<=x"0100";
m(5925)<=x"2029";
m(5926)<=x"bba8";
m(5927)<=x"bdff";
m(5928)<=x"ffff";
m(5929)<=x"ffff";
m(5930)<=x"88be";
m(5931)<=x"3f82";
m(5932)<=x"100b";
m(5952)<=x"0000";
m(5953)<=x"0000";
m(5954)<=x"0040";
m(5955)<=x"0780";
m(5956)<=x"0400";
m(5957)<=x"0050";
m(5958)<=x"81b1";
m(5959)<=x"5dff";
m(5960)<=x"ffff";
m(5961)<=x"ffff";
m(5962)<=x"82ef";
m(5963)<=x"1700";
m(5964)<=x"1002";
m(5984)<=x"0000";
m(5985)<=x"0000";
m(5986)<=x"0008";
m(5987)<=x"0788";
m(5988)<=x"0000";
m(5989)<=x"0045";
m(5990)<=x"e191";
m(5991)<=x"fbff";
m(5992)<=x"c7ff";
m(5993)<=x"ffff";
m(5994)<=x"8a58";
m(5995)<=x"5f90";
m(5996)<=x"0850";
m(6016)<=x"0000";
m(6017)<=x"0000";
m(6018)<=x"0050";
m(6019)<=x"07c0";
m(6020)<=x"0000";
m(6021)<=x"0000";
m(6022)<=x"c051";
m(6023)<=x"6afe";
m(6024)<=x"0fff";
m(6025)<=x"ffff";
m(6026)<=x"01f6";
m(6027)<=x"3f88";
m(6028)<=x"0004";
m(6048)<=x"0000";
m(6049)<=x"0000";
m(6050)<=x"0001";
m(6051)<=x"07e0";
m(6052)<=x"0000";
m(6053)<=x"0005";
m(6054)<=x"0010";
m(6055)<=x"11f8";
m(6056)<=x"0677";
m(6057)<=x"ffff";
m(6058)<=x"806d";
m(6059)<=x"87a0";
m(6060)<=x"0021";
m(6080)<=x"0000";
m(6081)<=x"0000";
m(6082)<=x"0000";
m(6083)<=x"07f0";
m(6084)<=x"0000";
m(6085)<=x"0000";
m(6086)<=x"0000";
m(6087)<=x"9950";
m(6088)<=x"2dff";
m(6089)<=x"ffff";
m(6090)<=x"0012";
m(6091)<=x"055a";
m(6092)<=x"0000";
m(6112)<=x"0000";
m(6113)<=x"0000";
m(6114)<=x"0048";
m(6115)<=x"07f8";
m(6116)<=x"0000";
m(6117)<=x"0000";
m(6118)<=x"0000";
m(6119)<=x"0530";
m(6120)<=x"1d77";
m(6121)<=x"ffff";
m(6122)<=x"0000";
m(6123)<=x"0002";
m(6124)<=x"2448";
m(6144)<=x"0000";
m(6145)<=x"0000";
m(6146)<=x"0000";
m(6147)<=x"03fc";
m(6148)<=x"0001";
m(6149)<=x"4000";
m(6150)<=x"0000";
m(6151)<=x"0270";
m(6152)<=x"1be7";
m(6153)<=x"ffff";
m(6154)<=x"0000";
m(6155)<=x"0000";
m(6156)<=x"0002";
m(6176)<=x"0000";
m(6177)<=x"0000";
m(6178)<=x"0002";
m(6179)<=x"3ffe";
m(6180)<=x"0010";
m(6181)<=x"0000";
m(6182)<=x"0000";
m(6183)<=x"99f0";
m(6184)<=x"10f7";
m(6185)<=x"ffff";
m(6186)<=x"0000";
m(6187)<=x"0000";
m(6188)<=x"0000";
m(6208)<=x"0000";
m(6209)<=x"0000";
m(6210)<=x"0040";
m(6211)<=x"1fff";
m(6212)<=x"0000";
m(6213)<=x"8000";
m(6214)<=x"0000";
m(6215)<=x"23f0";
m(6216)<=x"439f";
m(6217)<=x"ffff";
m(6218)<=x"0000";
m(6219)<=x"1000";
m(6220)<=x"0000";
m(6240)<=x"0000";
m(6241)<=x"0000";
m(6242)<=x"0004";
m(6243)<=x"1fff";
m(6244)<=x"0089";
m(6245)<=x"1000";
m(6246)<=x"0000";
m(6247)<=x"1df8";
m(6248)<=x"09bf";
m(6249)<=x"ffff";
m(6250)<=x"0594";
m(6251)<=x"0000";
m(6252)<=x"0000";
m(6272)<=x"0000";
m(6273)<=x"0000";
m(6274)<=x"0010";
m(6275)<=x"1fff";
m(6276)<=x"8090";
m(6277)<=x"0800";
m(6278)<=x"0000";
m(6279)<=x"57f8";
m(6280)<=x"835f";
m(6281)<=x"ffff";
m(6282)<=x"1b00";
m(6283)<=x"1000";
m(6284)<=x"0000";
m(6304)<=x"0000";
m(6305)<=x"0000";
m(6306)<=x"0000";
m(6307)<=x"1fff";
m(6308)<=x"c005";
m(6309)<=x"a220";
m(6310)<=x"0000";
m(6311)<=x"2a94";
m(6312)<=x"0e3f";
m(6313)<=x"ffff";
m(6314)<=x"6c58";
m(6315)<=x"0000";
m(6316)<=x"0000";
m(6336)<=x"0000";
m(6337)<=x"0000";
m(6338)<=x"0010";
m(6339)<=x"1fff";
m(6340)<=x"c008";
m(6341)<=x"0840";
m(6342)<=x"0000";
m(6343)<=x"66f8";
m(6344)<=x"0e7f";
m(6345)<=x"fffc";
m(6346)<=x"1ba0";
m(6347)<=x"8000";
m(6348)<=x"0000";
m(6368)<=x"0000";
m(6369)<=x"0000";
m(6370)<=x"0080";
m(6371)<=x"1fff";
m(6372)<=x"c009";
m(6373)<=x"a690";
m(6374)<=x"0002";
m(6375)<=x"1bfc";
m(6376)<=x"3e1f";
m(6377)<=x"fffc";
m(6378)<=x"2d02";
m(6379)<=x"0000";
m(6380)<=x"0000";
m(6400)<=x"0000";
m(6401)<=x"0000";
m(6402)<=x"0000";
m(6403)<=x"07ff";
m(6404)<=x"f008";
m(6405)<=x"856d";
m(6406)<=x"5fff";
m(6407)<=x"fbfc";
m(6408)<=x"3e97";
m(6409)<=x"fff9";
m(6410)<=x"5658";
m(6411)<=x"0000";
m(6412)<=x"0000";
m(6432)<=x"0000";
m(6433)<=x"0000";
m(6434)<=x"0000";
m(6435)<=x"07ff";
m(6436)<=x"f002";
m(6437)<=x"326f";
m(6438)<=x"f9ff";
m(6439)<=x"fff0";
m(6440)<=x"3c0f";
m(6441)<=x"fff8";
m(6442)<=x"6882";
m(6443)<=x"4000";
m(6444)<=x"0000";
m(6464)<=x"0000";
m(6465)<=x"0000";
m(6466)<=x"0000";
m(6467)<=x"03ff";
m(6468)<=x"f800";
m(6469)<=x"2bfb";
m(6470)<=x"fbff";
m(6471)<=x"ffe0";
m(6472)<=x"9c1f";
m(6473)<=x"fff0";
m(6474)<=x"1322";
m(6475)<=x"4000";
m(6476)<=x"0000";
m(6496)<=x"0000";
m(6497)<=x"0000";
m(6498)<=x"0000";
m(6499)<=x"00ff";
m(6500)<=x"f800";
m(6501)<=x"459f";
m(6502)<=x"ffff";
m(6503)<=x"ffc0";
m(6504)<=x"780f";
m(6505)<=x"fff1";
m(6506)<=x"8888";
m(6507)<=x"0000";
m(6508)<=x"0000";
m(6528)<=x"0000";
m(6529)<=x"0000";
m(6530)<=x"0000";
m(6531)<=x"00f8";
m(6532)<=x"fc00";
m(6533)<=x"0a5f";
m(6534)<=x"d6ff";
m(6535)<=x"ffc0";
m(6536)<=x"3c0f";
m(6537)<=x"fff0";
m(6538)<=x"3005";
m(6539)<=x"0000";
m(6540)<=x"0000";
m(6560)<=x"0000";
m(6561)<=x"0000";
m(6562)<=x"0000";
m(6563)<=x"00e0";
m(6564)<=x"fe00";
m(6565)<=x"51d6";
m(6566)<=x"ffff";
m(6567)<=x"ff80";
m(6568)<=x"7803";
m(6569)<=x"ffc5";
m(6570)<=x"8d50";
m(6571)<=x"8000";
m(6572)<=x"0000";
m(6592)<=x"0000";
m(6593)<=x"0000";
m(6594)<=x"0000";
m(6595)<=x"0001";
m(6596)<=x"fc00";
m(6597)<=x"0465";
m(6598)<=x"ebff";
m(6599)<=x"ff00";
m(6600)<=x"f803";
m(6601)<=x"7fc4";
m(6602)<=x"5005";
m(6603)<=x"0000";
m(6604)<=x"0000";
m(6624)<=x"0000";
m(6625)<=x"0000";
m(6626)<=x"0000";
m(6627)<=x"0001";
m(6628)<=x"fe00";
m(6629)<=x"1314";
m(6630)<=x"393f";
m(6631)<=x"ff00";
m(6632)<=x"f881";
m(6633)<=x"bfc1";
m(6634)<=x"4494";
m(6635)<=x"0000";
m(6636)<=x"0000";
m(6656)<=x"0000";
m(6657)<=x"0000";
m(6658)<=x"0000";
m(6659)<=x"0003";
m(6660)<=x"fe00";
m(6661)<=x"0049";
m(6662)<=x"002f";
m(6663)<=x"fc00";
m(6664)<=x"f000";
m(6665)<=x"8fc9";
m(6666)<=x"3012";
m(6667)<=x"0000";
m(6668)<=x"0000";
m(6688)<=x"0000";
m(6689)<=x"0000";
m(6690)<=x"0000";
m(6691)<=x"0002";
m(6692)<=x"fe00";
m(6693)<=x"0020";
m(6694)<=x"00a5";
m(6695)<=x"b041";
m(6696)<=x"f000";
m(6697)<=x"cf84";
m(6698)<=x"0848";
m(6699)<=x"0000";
m(6700)<=x"0000";
m(6720)<=x"0000";
m(6721)<=x"0000";
m(6722)<=x"0000";
m(6723)<=x"0000";
m(6724)<=x"fe00";
m(6725)<=x"0040";
m(6726)<=x"0009";
m(6727)<=x"63c1";
m(6728)<=x"f000";
m(6729)<=x"efb6";
m(6730)<=x"4104";
m(6731)<=x"0000";
m(6732)<=x"0000";
m(6752)<=x"0000";
m(6753)<=x"0000";
m(6754)<=x"0000";
m(6755)<=x"0000";
m(6756)<=x"3f00";
m(6757)<=x"0000";
m(6758)<=x"0000";
m(6759)<=x"8783";
m(6760)<=x"e000";
m(6761)<=x"3f0a";
m(6762)<=x"2014";
m(6763)<=x"0000";
m(6764)<=x"0000";
m(6784)<=x"0000";
m(6785)<=x"0000";
m(6786)<=x"0000";
m(6787)<=x"0000";
m(6788)<=x"0700";
m(6789)<=x"0000";
m(6790)<=x"0000";
m(6791)<=x"0383";
m(6792)<=x"f000";
m(6793)<=x"3742";
m(6794)<=x"0008";
m(6795)<=x"0000";
m(6796)<=x"0000";
m(6816)<=x"0000";
m(6817)<=x"0000";
m(6818)<=x"0000";
m(6819)<=x"0000";
m(6820)<=x"03c0";
m(6821)<=x"0000";
m(6822)<=x"0000";
m(6823)<=x"0183";
m(6824)<=x"f000";
m(6825)<=x"18b6";
m(6826)<=x"6464";
m(6827)<=x"0000";
m(6828)<=x"0000";
m(6848)<=x"0000";
m(6849)<=x"0000";
m(6850)<=x"0000";
m(6851)<=x"0000";
m(6852)<=x"00e0";
m(6853)<=x"0000";
m(6854)<=x"0003";
m(6855)<=x"4407";
m(6856)<=x"f000";
m(6857)<=x"0ca0";
m(6858)<=x"2028";
m(6859)<=x"0000";
m(6860)<=x"0000";
m(6880)<=x"0000";
m(6881)<=x"0000";
m(6882)<=x"0000";
m(6883)<=x"0000";
m(6884)<=x"0020";
m(6885)<=x"0000";
m(6886)<=x"000f";
m(6887)<=x"860f";
m(6888)<=x"f000";
m(6889)<=x"0ddc";
m(6890)<=x"0010";
m(6891)<=x"0000";
m(6892)<=x"0000";
m(6912)<=x"0000";
m(6913)<=x"0000";
m(6914)<=x"0000";
m(6915)<=x"0000";
m(6916)<=x"0000";
m(6917)<=x"0000";
m(6918)<=x"0003";
m(6919)<=x"dc07";
m(6920)<=x"fc00";
m(6921)<=x"0ce0";
m(6922)<=x"0090";
m(6923)<=x"0000";
m(6924)<=x"0000";
m(6944)<=x"0000";
m(6945)<=x"0000";
m(6946)<=x"0000";
m(6947)<=x"0000";
m(6948)<=x"0000";
m(6949)<=x"0000";
m(6950)<=x"0000";
m(6951)<=x"e40f";
m(6952)<=x"fe00";
m(6953)<=x"0826";
m(6954)<=x"0020";
m(6955)<=x"0000";
m(6956)<=x"0000";
m(6976)<=x"0000";
m(6977)<=x"0000";
m(6978)<=x"0000";
m(6979)<=x"0000";
m(6980)<=x"0000";
m(6981)<=x"0000";
m(6982)<=x"0000";
m(6983)<=x"701f";
m(6984)<=x"fe00";
m(6985)<=x"00b0";
m(6986)<=x"0000";
m(6987)<=x"0000";
m(6988)<=x"0000";
m(7008)<=x"0000";
m(7009)<=x"0000";
m(7010)<=x"0000";
m(7011)<=x"0000";
m(7012)<=x"0000";
m(7013)<=x"0000";
m(7014)<=x"0000";
m(7015)<=x"381f";
m(7016)<=x"ff00";
m(7017)<=x"000c";
m(7018)<=x"0000";
m(7019)<=x"0000";
m(7020)<=x"0000";
m(7040)<=x"0000";
m(7041)<=x"0000";
m(7042)<=x"0000";
m(7043)<=x"0000";
m(7044)<=x"0000";
m(7045)<=x"0000";
m(7046)<=x"0000";
m(7047)<=x"001f";
m(7048)<=x"fe00";
m(7049)<=x"0010";
m(7050)<=x"0000";
m(7051)<=x"0000";
m(7052)<=x"0000";
m(7072)<=x"0000";
m(7073)<=x"0000";
m(7074)<=x"0000";
m(7075)<=x"0000";
m(7076)<=x"0000";
m(7077)<=x"0000";
m(7078)<=x"0000";
m(7079)<=x"001a";
m(7080)<=x"0808";
m(7081)<=x"0084";
m(7082)<=x"0040";
m(7083)<=x"0000";
m(7084)<=x"0000";
m(7104)<=x"0000";
m(7105)<=x"0000";
m(7106)<=x"0000";
m(7107)<=x"0000";
m(7108)<=x"0000";
m(7109)<=x"0000";
m(7110)<=x"0000";
m(7111)<=x"0000";
m(7112)<=x"0004";
m(7113)<=x"c102";
m(7114)<=x"0000";
m(7115)<=x"0000";
m(7116)<=x"0000";
m(7136)<=x"0000";
m(7137)<=x"0000";
m(7138)<=x"0000";
m(7139)<=x"0000";
m(7140)<=x"0000";
m(7141)<=x"0000";
m(7142)<=x"0000";
m(7143)<=x"0000";
m(7144)<=x"0007";
m(7145)<=x"e010";
m(7146)<=x"0000";
m(7147)<=x"0000";
m(7148)<=x"0000";
m(7168)<=x"0000";
m(7169)<=x"0000";
m(7170)<=x"0000";
m(7171)<=x"0000";
m(7172)<=x"0000";
m(7173)<=x"0000";
m(7174)<=x"0000";
m(7175)<=x"0000";
m(7176)<=x"0001";
m(7177)<=x"f000";
m(7178)<=x"0000";
m(7179)<=x"0000";
m(7180)<=x"0000";
m(7200)<=x"0000";
m(7201)<=x"0000";
m(7202)<=x"0000";
m(7203)<=x"0000";
m(7204)<=x"0000";
m(7205)<=x"0000";
m(7206)<=x"0000";
m(7207)<=x"0000";
m(7208)<=x"0001";
m(7209)<=x"7000";
m(7210)<=x"0000";
m(7211)<=x"0000";
m(7212)<=x"0000";
m(7232)<=x"0000";
m(7233)<=x"0000";
m(7234)<=x"0000";
m(7235)<=x"0000";
m(7236)<=x"0000";
m(7237)<=x"0000";
m(7238)<=x"0000";
m(7239)<=x"0000";
m(7240)<=x"0000";
m(7241)<=x"f810";
m(7242)<=x"0000";
m(7243)<=x"0000";
m(7244)<=x"0000";
m(7264)<=x"0000";
m(7265)<=x"0000";
m(7266)<=x"0000";
m(7267)<=x"0000";
m(7268)<=x"0000";
m(7269)<=x"0000";
m(7270)<=x"0000";
m(7271)<=x"0000";
m(7272)<=x"0000";
m(7273)<=x"7802";
m(7274)<=x"0000";
m(7275)<=x"0000";
m(7276)<=x"0000";
m(7296)<=x"0000";
m(7297)<=x"0000";
m(7298)<=x"0000";
m(7299)<=x"0000";
m(7300)<=x"0000";
m(7301)<=x"0000";
m(7302)<=x"0000";
m(7303)<=x"0000";
m(7304)<=x"0000";
m(7305)<=x"3840";
m(7306)<=x"0000";
m(7307)<=x"0000";
m(7308)<=x"0000";
m(7328)<=x"0000";
m(7329)<=x"0000";
m(7330)<=x"0000";
m(7331)<=x"0000";
m(7332)<=x"0000";
m(7333)<=x"0000";
m(7334)<=x"0000";
m(7335)<=x"0000";
m(7336)<=x"0000";
m(7337)<=x"1e80";
m(7338)<=x"0000";
m(7339)<=x"0000";
m(7340)<=x"0000";
m(7360)<=x"0000";
m(7361)<=x"0000";
m(7362)<=x"0000";
m(7363)<=x"0000";
m(7364)<=x"0000";
m(7365)<=x"0000";
m(7366)<=x"0000";
m(7367)<=x"0000";
m(7368)<=x"0000";
m(7369)<=x"1f48";
m(7370)<=x"0000";
m(7371)<=x"0000";
m(7372)<=x"0000";
m(7392)<=x"0000";
m(7393)<=x"0000";
m(7394)<=x"0000";
m(7395)<=x"0000";
m(7396)<=x"0000";
m(7397)<=x"0000";
m(7398)<=x"0000";
m(7399)<=x"0000";
m(7400)<=x"0000";
m(7401)<=x"1c80";
m(7402)<=x"0000";
m(7403)<=x"0000";
m(7404)<=x"0000";
m(7424)<=x"0000";
m(7425)<=x"0000";
m(7426)<=x"0000";
m(7427)<=x"0000";
m(7428)<=x"0000";
m(7429)<=x"0000";
m(7430)<=x"0000";
m(7431)<=x"0000";
m(7432)<=x"0000";
m(7433)<=x"0f80";
m(7434)<=x"0000";
m(7435)<=x"0000";
m(7436)<=x"0000";
m(7456)<=x"0000";
m(7457)<=x"0000";
m(7458)<=x"0000";
m(7459)<=x"0000";
m(7460)<=x"0000";
m(7461)<=x"0000";
m(7462)<=x"0000";
m(7463)<=x"0000";
m(7464)<=x"0026";
m(7465)<=x"be30";
m(7466)<=x"0000";
m(7467)<=x"0000";
m(7468)<=x"0000";
m(7488)<=x"0000";
m(7489)<=x"0000";
m(7490)<=x"0000";
m(7491)<=x"0000";
m(7492)<=x"0000";
m(7493)<=x"0000";
m(7494)<=x"0000";
m(7495)<=x"0000";
m(7496)<=x"0025";
m(7497)<=x"7f80";
m(7498)<=x"0000";
m(7499)<=x"0000";
m(7500)<=x"0000";
m(7520)<=x"0000";
m(7521)<=x"0000";
m(7522)<=x"0000";
m(7523)<=x"0000";
m(7524)<=x"0000";
m(7525)<=x"0000";
m(7526)<=x"0000";
m(7527)<=x"0000";
m(7528)<=x"0000";
m(7529)<=x"4be0";
m(7530)<=x"0000";
m(7531)<=x"0000";
m(7532)<=x"0000";
m(7552)<=x"0000";
m(7553)<=x"0000";
m(7554)<=x"0000";
m(7555)<=x"0000";
m(7556)<=x"0000";
m(7557)<=x"0000";
m(7558)<=x"0000";
m(7559)<=x"0000";
m(7560)<=x"0001";
m(7561)<=x"7700";
m(7562)<=x"0000";
m(7563)<=x"0000";
m(7564)<=x"0000";
m(7584)<=x"0000";
m(7585)<=x"0000";
m(7586)<=x"0000";
m(7587)<=x"0000";
m(7588)<=x"0000";
m(7589)<=x"0000";
m(7590)<=x"0000";
m(7591)<=x"0000";
m(7592)<=x"0000";
m(7593)<=x"4180";
m(7594)<=x"0000";
m(7595)<=x"0000";
m(7596)<=x"0000";
m(7616)<=x"0000";
m(7617)<=x"0000";
m(7618)<=x"0000";
m(7619)<=x"0000";
m(7620)<=x"0000";
m(7621)<=x"0000";
m(7622)<=x"0000";
m(7623)<=x"0000";
m(7624)<=x"0006";
m(7625)<=x"0180";
m(7626)<=x"0000";
m(7627)<=x"0000";
m(7628)<=x"0000";
m(7648)<=x"0000";
m(7649)<=x"0000";
m(7650)<=x"0000";
m(7651)<=x"0000";
m(7652)<=x"0000";
m(7653)<=x"0000";
m(7654)<=x"0000";
m(7655)<=x"0000";
m(7656)<=x"0000";
m(7657)<=x"01c0";
m(7658)<=x"0000";
m(7659)<=x"0000";
m(7660)<=x"0000";
m(7680)<=x"0000";
m(7681)<=x"0000";
m(7682)<=x"0000";
m(7683)<=x"0000";
m(7684)<=x"0000";
m(7685)<=x"0000";
m(7686)<=x"0000";
m(7687)<=x"0000";
m(7688)<=x"0000";
m(7689)<=x"00e0";
m(7690)<=x"0000";
m(7691)<=x"0000";
m(7692)<=x"0000";
m(7712)<=x"0000";
m(7713)<=x"0000";
m(7714)<=x"0000";
m(7715)<=x"0000";
m(7716)<=x"0000";
m(7717)<=x"0000";
m(7718)<=x"0000";
m(7719)<=x"0000";
m(7720)<=x"0000";
m(7721)<=x"0060";
m(7722)<=x"0000";
m(7723)<=x"0000";
m(7724)<=x"0000";
m(7744)<=x"0000";
m(7745)<=x"0000";
m(7746)<=x"0000";
m(7747)<=x"0000";
m(7748)<=x"0000";
m(7749)<=x"0000";
m(7750)<=x"0000";
m(7751)<=x"0000";
m(7752)<=x"0000";
m(7753)<=x"0000";
m(7754)<=x"0000";
m(7755)<=x"0000";
m(7756)<=x"0000";
m(7776)<=x"0000";
m(7777)<=x"0000";
m(7778)<=x"0000";
m(7779)<=x"0000";
m(7780)<=x"0000";
m(7781)<=x"0000";
m(7782)<=x"0000";
m(7783)<=x"0000";
m(7784)<=x"0000";
m(7785)<=x"0000";
m(7786)<=x"0000";
m(7787)<=x"0000";
m(7788)<=x"0000";
m(7808)<=x"0000";
m(7809)<=x"0000";
m(7810)<=x"0000";
m(7811)<=x"0000";
m(7812)<=x"0000";
m(7813)<=x"0000";
m(7814)<=x"0000";
m(7815)<=x"0000";
m(7816)<=x"0000";
m(7817)<=x"0200";
m(7818)<=x"0000";
m(7819)<=x"0000";
m(7820)<=x"0000";
m(7840)<=x"0000";
m(7841)<=x"0000";
m(7842)<=x"0000";
m(7843)<=x"0000";
m(7844)<=x"0000";
m(7845)<=x"0000";
m(7846)<=x"0000";
m(7847)<=x"0000";
m(7848)<=x"0000";
m(7849)<=x"0000";
m(7850)<=x"0000";
m(7851)<=x"0000";
m(7852)<=x"0000";
m(7872)<=x"0000";
m(7873)<=x"0000";
m(7874)<=x"0000";
m(7875)<=x"0000";
m(7876)<=x"0000";
m(7877)<=x"0000";
m(7878)<=x"0000";
m(7879)<=x"0000";
m(7880)<=x"0000";
m(7881)<=x"0000";
m(7882)<=x"0000";
m(7883)<=x"0000";
m(7884)<=x"0000";
m(7904)<=x"0000";
m(7905)<=x"0000";
m(7906)<=x"0000";
m(7907)<=x"0000";
m(7908)<=x"0000";
m(7909)<=x"0000";
m(7910)<=x"0000";
m(7911)<=x"0000";
m(7912)<=x"0000";
m(7913)<=x"0000";
m(7914)<=x"0000";
m(7915)<=x"0000";
m(7916)<=x"0000";
m(7936)<=x"0000";
m(7937)<=x"0000";
m(7938)<=x"0000";
m(7939)<=x"0000";
m(7940)<=x"0000";
m(7941)<=x"0000";
m(7942)<=x"0000";
m(7943)<=x"0000";
m(7944)<=x"0000";
m(7945)<=x"0000";
m(7946)<=x"0000";
m(7947)<=x"0000";
m(7948)<=x"0000";
m(7968)<=x"0000";
m(7969)<=x"0000";
m(7970)<=x"0000";
m(7971)<=x"0000";
m(7972)<=x"0000";
m(7973)<=x"0000";
m(7974)<=x"0000";
m(7975)<=x"0000";
m(7976)<=x"0000";
m(7977)<=x"0000";
m(7978)<=x"0000";
m(7979)<=x"0000";
m(7980)<=x"0000";
m(8000)<=x"0000";
m(8001)<=x"0000";
m(8002)<=x"0000";
m(8003)<=x"0000";
m(8004)<=x"0000";
m(8005)<=x"0000";
m(8006)<=x"0000";
m(8007)<=x"0000";
m(8008)<=x"0000";
m(8009)<=x"0000";
m(8010)<=x"0000";
m(8011)<=x"0000";
m(8012)<=x"0000";

   process(CLK)
	 begin 
		if (CLK'event AND CLK='1') then
			D <= m(conv_integer(AD));
		end if;
	end process;
end Behavioral;

