----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:16:29 04/19/2013 
-- Design Name: 
-- Module Name:    VRAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity VRAM is
	port (Clk		: in 	std_logic;
			CE			: in 	std_logic;
			Enable_w	: in 	std_logic;
			Addr_w	: in 	std_logic_vector	(18 downto 0);
			Addr_r	: in 	std_logic_vector	(18 downto 0);
			Data_in	: in 	std_logic_vector	(7 downto 0);
			Data_out	: out std_logic_vector	(7 downto 0));
end VRAM;

architecture Behavioral of VRAM is
	type ram_type is array ((2**19)-1 downto 0) of std_logic_vector (7 downto 0);
	signal VRAM: ram_type := (
		19555 => x"FF",
		20579 => x"FF",
		21603 => x"FF",
		22627 => x"FF",
		23651 => x"FF",
		24675 => x"FF",
		25699 => x"FF",
		26723 => x"FF",
		27747 => x"FF",
		28771 => x"FF",
		29795 => x"FF",
		30819 => x"FF",
		31843 => x"FF",
		32867 => x"FF",
		33891 => x"FF",
		34915 => x"FF",
		35939 => x"FF",
		36963 => x"FF",
		37987 => x"FF",
		39011 => x"FF",
		40035 => x"FF",
		41059 => x"FF",
		42083 => x"FF",
		43107 => x"FF",
		44131 => x"FF",
		45155 => x"FF",
		46179 => x"FF",
		47203 => x"FF",
		48227 => x"FF",
		49251 => x"FF",
		50275 => x"FF",
		51299 => x"FF",
		52323 => x"FF",
		53347 => x"FF",
		54371 => x"FF",
		55395 => x"FF",
		56419 => x"FF",
		57443 => x"FF",
		58467 => x"FF",
		59491 => x"FF",
		60515 => x"FF",
		61539 => x"FF",
		62563 => x"FF",
		63587 => x"FF",
		64611 => x"FF",
		65635 => x"FF",
		66659 => x"FF",
		67683 => x"FF",
		68707 => x"FF",
		69731 => x"FF",
		70755 => x"FF",
		71779 => x"FF",
		72803 => x"FF",
		73827 => x"FF",
		74851 => x"FF",
		75875 => x"FF",
		76899 => x"FF",
		77923 => x"FF",
		78947 => x"FF",
		79971 => x"FF",
		80995 => x"FF",
		82019 => x"FF",
		83043 => x"FF",
		84067 => x"FF",
		85091 => x"FF",
		86115 => x"FF",
		87139 => x"FF",
		88163 => x"FF",
		89187 => x"FF",
		90211 => x"FF",
		91235 => x"FF",
		92259 => x"FF",
		93283 => x"FF",
		94307 => x"FF",
		95331 => x"FF",
		96355 => x"FF",
		97379 => x"FF",
		98403 => x"FF",
		99427 => x"FF",
		100451 => x"FF",
		101475 => x"FF",
		102499 => x"FF",
		103523 => x"FF",
		104547 => x"FF",
		105571 => x"FF",
		106595 => x"FF",
		107619 => x"FF",
		108643 => x"FF",
		109667 => x"FF",
		110691 => x"FF",
		111715 => x"FF",
		112739 => x"FF",
		113763 => x"FF",
		114787 => x"FF",
		115811 => x"FF",
		116835 => x"FF",
		117859 => x"FF",
		118883 => x"FF",
		119907 => x"FF",
		120931 => x"FF",
		121955 => x"FF",
		122979 => x"FF",
		124003 => x"FF",
		125027 => x"FF",
		126051 => x"FF",
		127075 => x"FF",
		128099 => x"FF",
		129123 => x"FF",
		130147 => x"FF",
		131171 => x"FF",
		132195 => x"FF",
		133219 => x"FF",
		134243 => x"FF",
		135267 => x"FF",
		136291 => x"FF",
		137315 => x"FF",
		138339 => x"FF",
		139363 => x"FF",
		140387 => x"FF",
		141411 => x"FF",
		142435 => x"FF",
		143459 => x"FF",
		144483 => x"FF",
		145507 => x"FF",
		146531 => x"FF",
		147555 => x"FF",
		148579 => x"FF",
		149603 => x"FF",
		150627 => x"FF",
		151651 => x"FF",
		152675 => x"FF",
		153699 => x"FF",
		154723 => x"FF",
		155747 => x"FF",
		156771 => x"FF",
		157795 => x"FF",
		158819 => x"FF",
		159843 => x"FF",
		160867 => x"FF",
		161891 => x"FF",
		162915 => x"FF",
		163939 => x"FF",
		164963 => x"FF",
		165987 => x"FF",
		167011 => x"FF",
		168035 => x"FF",
		169059 => x"FF",
		170083 => x"FF",
		171107 => x"FF",
		172131 => x"FF",
		173155 => x"FF",
		174179 => x"FF",
		175203 => x"FF",
		176227 => x"FF",
		177251 => x"FF",
		178275 => x"FF",
		179299 => x"FF",
		180323 => x"FF",
		181347 => x"FF",
		182371 => x"FF",
		183395 => x"FF",
		184419 => x"FF",
		185443 => x"FF",
		186467 => x"FF",
		187491 => x"FF",
		188515 => x"FF",
		189539 => x"FF",
		190563 => x"FF",
		191587 => x"FF",
		192611 => x"FF",
		193635 => x"FF",
		194659 => x"FF",
		195683 => x"FF",
		196707 => x"FF",
		197731 => x"FF",
		198755 => x"FF",
		199779 => x"FF",
		200803 => x"FF",
		201827 => x"FF",
		202851 => x"FF",
		203875 => x"FF",
		204899 => x"FF",
		205923 => x"FF",
		206947 => x"FF",
		207971 => x"FF",
		208995 => x"FF",
		210019 => x"FF",
		211043 => x"FF",
		212067 => x"FF",
		213091 => x"FF",
		214115 => x"FF",
		215139 => x"FF",
		216163 => x"FF",
		217187 => x"FF",
		218211 => x"FF",
		219235 => x"FF",
		220259 => x"FF",
		221283 => x"FF",
		222307 => x"FF",
		223331 => x"FF",
		224355 => x"FF",
		225379 => x"FF",
		226403 => x"FF",
		227427 => x"FF",
		228451 => x"FF",
		229475 => x"FF",
		230499 => x"FF",
		231523 => x"FF",
		232547 => x"FF",
		233571 => x"FF",
		234595 => x"FF",
		235619 => x"FF",
		236643 => x"FF",
		237667 => x"FF",
		238691 => x"FF",
		239715 => x"FF",
		240739 => x"FF",
		241763 => x"FF",
		242787 => x"FF",
		243811 => x"FF",
		244835 => x"FF",
		245859 => x"FF",
		246883 => x"FF",
		247907 => x"FF",
		248931 => x"FF",
		249955 => x"FF",
		250979 => x"FF",
		252003 => x"FF",
		253027 => x"FF",
		254051 => x"FF",
		255075 => x"FF",
		256099 => x"FF",
		257123 => x"FF",
		258147 => x"FF",
		259171 => x"FF",
		260195 => x"FF",
		261219 => x"FF",
		262243 => x"FF",
		263267 => x"FF",
		264291 => x"FF",
		265315 => x"FF",
		266339 => x"FF",
		267363 => x"FF",
		268387 => x"FF",
		269411 => x"FF",
		270435 => x"FF",
		271459 => x"FF",
		272483 => x"FF",
		273507 => x"FF",
		274531 => x"FF",
		275555 => x"FF",
		276579 => x"FF",
		277603 => x"FF",
		278627 => x"FF",
		279651 => x"FF",
		280675 => x"FF",
		281699 => x"FF",
		282723 => x"FF",
		283747 => x"FF",
		284771 => x"FF",
		285795 => x"FF",
		286819 => x"FF",
		287843 => x"FF",
		288867 => x"FF",
		289891 => x"FF",
		290915 => x"FF",
		291939 => x"FF",
		292963 => x"FF",
		293987 => x"FF",
		295011 => x"FF",
		296035 => x"FF",
		297059 => x"FF",
		298083 => x"FF",
		299107 => x"FF",
		300131 => x"FF",
		301155 => x"FF",
		302179 => x"FF",
		303203 => x"FF",
		304227 => x"FF",
		305251 => x"FF",
		306275 => x"FF",
		307299 => x"FF",
		308323 => x"FF",
		309347 => x"FF",
		310371 => x"FF",
		311395 => x"FF",
		312419 => x"FF",
		313443 => x"FF",
		314467 => x"FF",
		315491 => x"FF",
		316515 => x"FF",
		317539 => x"FF",
		318563 => x"FF",
		319587 => x"FF",
		320611 => x"FF",
		321635 => x"FF",
		322659 => x"FF",
		323683 => x"FF",
		324707 => x"FF",
		325731 => x"FF",
		326755 => x"FF",
		327779 => x"FF",
		328803 => x"FF",
		329827 => x"FF",
		330851 => x"FF",
		331875 => x"FF",
		332899 => x"FF",
		333923 => x"FF",
		334947 => x"FF",
		335971 => x"FF",
		336995 => x"FF",
		338019 => x"FF",
		339043 => x"FF",
		340067 => x"FF",
		341091 => x"FF",
		342115 => x"FF",
		343139 => x"FF",
		344163 => x"FF",
		345187 => x"FF",
		346211 => x"FF",
		347235 => x"FF",
		348259 => x"FF",
		349283 => x"FF",
		350307 => x"FF",
		351331 => x"FF",
		352355 => x"FF",
		353379 => x"FF",
		354403 => x"FF",
		355427 => x"FF",
		356451 => x"FF",
		357475 => x"FF",
		358499 => x"FF",
		359523 => x"FF",
		360547 => x"FF",
		361571 => x"FF",
		362595 => x"FF",
		363619 => x"FF",
		364643 => x"FF",
		365667 => x"FF",
		366691 => x"FF",
		367715 => x"FF",
		368739 => x"FF",
		369763 => x"FF",
		370787 => x"FF",
		371811 => x"FF",
		372835 => x"FF",
		373859 => x"FF",
		374883 => x"FF",
		375907 => x"FF",
		376931 => x"FF",
		377955 => x"FF",
		378979 => x"FF",
		380003 => x"FF",
		381027 => x"FF",
		382051 => x"FF",
		383075 => x"FF",
		384099 => x"FF",
		385123 => x"FF",
		386147 => x"FF",
		387171 => x"FF",
		388195 => x"FF",
		389219 => x"FF",
		390243 => x"FF",
		391267 => x"FF",
		392291 => x"FF",
		393315 => x"FF",
		394339 => x"FF",
		395363 => x"FF",
		396387 => x"FF",
		397411 => x"FF",
		398435 => x"FF",
		399459 => x"FF",
		400483 => x"FF",
		401507 => x"FF",
		402531 => x"FF",
		403555 => x"FF",
		404579 => x"FF",
		405603 => x"FF",
		406627 => x"FF",
		407651 => x"FF",
		408675 => x"FF",
		409699 => x"FF",
		410723 => x"FF",
		411747 => x"FF",
		412771 => x"FF",
		413795 => x"FF",
		414819 => x"FF",
		415843 => x"FF",
		416867 => x"FF",
		417891 => x"FF",
		418915 => x"FF",
		419939 => x"FF",
		420963 => x"FF",
		421987 => x"FF",
		423011 => x"FF",
		424035 => x"FF",
		425059 => x"FF",
		426083 => x"FF",
		427107 => x"FF",
		428131 => x"FF",
		429155 => x"FF",
		430179 => x"FF",
		431203 => x"FF",
		432227 => x"FF",
		433251 => x"FF",
		434275 => x"FF",
		435299 => x"FF",
		436323 => x"FF",
		437347 => x"FF",
		438371 => x"FF",
		439395 => x"FF",
		440419 => x"FF",
		441443 => x"FF",
		442467 => x"FF",
		443491 => x"FF",
		444515 => x"FF",
		445539 => x"FF",
		446563 => x"FF",
		447587 => x"FF",
		448611 => x"FF",
		449635 => x"FF",
		450659 => x"FF",
		451683 => x"FF",
		452707 => x"FF",
		453731 => x"FF",
		454755 => x"FF",
		455779 => x"FF",
		456803 => x"FF",
		457827 => x"FF",
		458851 => x"FF",
		459875 => x"FF",
		460899 => x"FF",
		461923 => x"FF",
		462947 => x"FF",
		463971 => x"FF",
		464995 => x"FF",
		466019 => x"FF",
		467043 => x"FF",
		468067 => x"FF",
		469091 => x"FF",
		19556 => x"FF",
		20580 => x"FF",
		21604 => x"FF",
		22628 => x"FF",
		23652 => x"FF",
		24676 => x"FF",
		25700 => x"FF",
		26724 => x"FF",
		27748 => x"FF",
		28772 => x"FF",
		29796 => x"FF",
		30820 => x"FF",
		31844 => x"FF",
		32868 => x"FF",
		33892 => x"FF",
		34916 => x"FF",
		35940 => x"FF",
		36964 => x"FF",
		37988 => x"FF",
		39012 => x"FF",
		40036 => x"FF",
		41060 => x"FF",
		42084 => x"FF",
		43108 => x"FF",
		44132 => x"FF",
		45156 => x"FF",
		46180 => x"FF",
		47204 => x"FF",
		48228 => x"FF",
		49252 => x"FF",
		50276 => x"FF",
		51300 => x"FF",
		52324 => x"FF",
		53348 => x"FF",
		54372 => x"FF",
		55396 => x"FF",
		56420 => x"FF",
		57444 => x"FF",
		58468 => x"FF",
		59492 => x"FF",
		60516 => x"FF",
		61540 => x"FF",
		62564 => x"FF",
		63588 => x"FF",
		64612 => x"FF",
		65636 => x"FF",
		66660 => x"FF",
		67684 => x"FF",
		68708 => x"FF",
		69732 => x"FF",
		70756 => x"FF",
		71780 => x"FF",
		72804 => x"FF",
		73828 => x"FF",
		74852 => x"FF",
		75876 => x"FF",
		76900 => x"FF",
		77924 => x"FF",
		78948 => x"FF",
		79972 => x"FF",
		80996 => x"FF",
		82020 => x"FF",
		83044 => x"FF",
		84068 => x"FF",
		85092 => x"FF",
		86116 => x"FF",
		87140 => x"FF",
		88164 => x"FF",
		89188 => x"FF",
		90212 => x"FF",
		91236 => x"FF",
		92260 => x"FF",
		93284 => x"FF",
		94308 => x"FF",
		95332 => x"FF",
		96356 => x"FF",
		97380 => x"FF",
		98404 => x"FF",
		99428 => x"FF",
		100452 => x"FF",
		101476 => x"FF",
		102500 => x"FF",
		103524 => x"FF",
		104548 => x"FF",
		105572 => x"FF",
		106596 => x"FF",
		107620 => x"FF",
		108644 => x"FF",
		109668 => x"FF",
		110692 => x"FF",
		111716 => x"FF",
		112740 => x"FF",
		113764 => x"FF",
		114788 => x"FF",
		115812 => x"FF",
		116836 => x"FF",
		117860 => x"FF",
		118884 => x"FF",
		119908 => x"FF",
		120932 => x"FF",
		121956 => x"FF",
		122980 => x"FF",
		124004 => x"FF",
		125028 => x"FF",
		126052 => x"FF",
		127076 => x"FF",
		128100 => x"FF",
		129124 => x"FF",
		130148 => x"FF",
		131172 => x"FF",
		132196 => x"FF",
		133220 => x"FF",
		134244 => x"FF",
		135268 => x"FF",
		136292 => x"FF",
		137316 => x"FF",
		138340 => x"FF",
		139364 => x"FF",
		140388 => x"FF",
		141412 => x"FF",
		142436 => x"FF",
		143460 => x"FF",
		144484 => x"FF",
		145508 => x"FF",
		146532 => x"FF",
		147556 => x"FF",
		148580 => x"FF",
		149604 => x"FF",
		150628 => x"FF",
		151652 => x"FF",
		152676 => x"FF",
		153700 => x"FF",
		154724 => x"FF",
		155748 => x"FF",
		156772 => x"FF",
		157796 => x"FF",
		158820 => x"FF",
		159844 => x"FF",
		160868 => x"FF",
		161892 => x"FF",
		162916 => x"FF",
		163940 => x"FF",
		164964 => x"FF",
		165988 => x"FF",
		167012 => x"FF",
		168036 => x"FF",
		169060 => x"FF",
		170084 => x"FF",
		171108 => x"FF",
		172132 => x"FF",
		173156 => x"FF",
		174180 => x"FF",
		175204 => x"FF",
		176228 => x"FF",
		177252 => x"FF",
		178276 => x"FF",
		179300 => x"FF",
		180324 => x"FF",
		181348 => x"FF",
		182372 => x"FF",
		183396 => x"FF",
		184420 => x"FF",
		185444 => x"FF",
		186468 => x"FF",
		187492 => x"FF",
		188516 => x"FF",
		189540 => x"FF",
		190564 => x"FF",
		191588 => x"FF",
		192612 => x"FF",
		193636 => x"FF",
		194660 => x"FF",
		195684 => x"FF",
		196708 => x"FF",
		197732 => x"FF",
		198756 => x"FF",
		199780 => x"FF",
		200804 => x"FF",
		201828 => x"FF",
		202852 => x"FF",
		203876 => x"FF",
		204900 => x"FF",
		205924 => x"FF",
		206948 => x"FF",
		207972 => x"FF",
		208996 => x"FF",
		210020 => x"FF",
		211044 => x"FF",
		212068 => x"FF",
		213092 => x"FF",
		214116 => x"FF",
		215140 => x"FF",
		216164 => x"FF",
		217188 => x"FF",
		218212 => x"FF",
		219236 => x"FF",
		220260 => x"FF",
		221284 => x"FF",
		222308 => x"FF",
		223332 => x"FF",
		224356 => x"FF",
		225380 => x"FF",
		226404 => x"FF",
		227428 => x"FF",
		228452 => x"FF",
		229476 => x"FF",
		230500 => x"FF",
		231524 => x"FF",
		232548 => x"FF",
		233572 => x"FF",
		234596 => x"FF",
		235620 => x"FF",
		236644 => x"FF",
		237668 => x"FF",
		238692 => x"FF",
		239716 => x"FF",
		240740 => x"FF",
		241764 => x"FF",
		242788 => x"FF",
		243812 => x"FF",
		244836 => x"FF",
		245860 => x"FF",
		246884 => x"FF",
		247908 => x"FF",
		248932 => x"FF",
		249956 => x"FF",
		250980 => x"FF",
		252004 => x"FF",
		253028 => x"FF",
		254052 => x"FF",
		255076 => x"FF",
		256100 => x"FF",
		257124 => x"FF",
		258148 => x"FF",
		259172 => x"FF",
		260196 => x"FF",
		261220 => x"FF",
		262244 => x"FF",
		263268 => x"FF",
		264292 => x"FF",
		265316 => x"FF",
		266340 => x"FF",
		267364 => x"FF",
		268388 => x"FF",
		269412 => x"FF",
		270436 => x"FF",
		271460 => x"FF",
		272484 => x"FF",
		273508 => x"FF",
		274532 => x"FF",
		275556 => x"FF",
		276580 => x"FF",
		277604 => x"FF",
		278628 => x"FF",
		279652 => x"FF",
		280676 => x"FF",
		281700 => x"FF",
		282724 => x"FF",
		283748 => x"FF",
		284772 => x"FF",
		285796 => x"FF",
		286820 => x"FF",
		287844 => x"FF",
		288868 => x"FF",
		289892 => x"FF",
		290916 => x"FF",
		291940 => x"FF",
		292964 => x"FF",
		293988 => x"FF",
		295012 => x"FF",
		296036 => x"FF",
		297060 => x"FF",
		298084 => x"FF",
		299108 => x"FF",
		300132 => x"FF",
		301156 => x"FF",
		302180 => x"FF",
		303204 => x"FF",
		304228 => x"FF",
		305252 => x"FF",
		306276 => x"FF",
		307300 => x"FF",
		308324 => x"FF",
		309348 => x"FF",
		310372 => x"FF",
		311396 => x"FF",
		312420 => x"FF",
		313444 => x"FF",
		314468 => x"FF",
		315492 => x"FF",
		316516 => x"FF",
		317540 => x"FF",
		318564 => x"FF",
		319588 => x"FF",
		320612 => x"FF",
		321636 => x"FF",
		322660 => x"FF",
		323684 => x"FF",
		324708 => x"FF",
		325732 => x"FF",
		326756 => x"FF",
		327780 => x"FF",
		328804 => x"FF",
		329828 => x"FF",
		330852 => x"FF",
		331876 => x"FF",
		332900 => x"FF",
		333924 => x"FF",
		334948 => x"FF",
		335972 => x"FF",
		336996 => x"FF",
		338020 => x"FF",
		339044 => x"FF",
		340068 => x"FF",
		341092 => x"FF",
		342116 => x"FF",
		343140 => x"FF",
		344164 => x"FF",
		345188 => x"FF",
		346212 => x"FF",
		347236 => x"FF",
		348260 => x"FF",
		349284 => x"FF",
		350308 => x"FF",
		351332 => x"FF",
		352356 => x"FF",
		353380 => x"FF",
		354404 => x"FF",
		355428 => x"FF",
		356452 => x"FF",
		357476 => x"FF",
		358500 => x"FF",
		359524 => x"FF",
		360548 => x"FF",
		361572 => x"FF",
		362596 => x"FF",
		363620 => x"FF",
		364644 => x"FF",
		365668 => x"FF",
		366692 => x"FF",
		367716 => x"FF",
		368740 => x"FF",
		369764 => x"FF",
		370788 => x"FF",
		371812 => x"FF",
		372836 => x"FF",
		373860 => x"FF",
		374884 => x"FF",
		375908 => x"FF",
		376932 => x"FF",
		377956 => x"FF",
		378980 => x"FF",
		380004 => x"FF",
		381028 => x"FF",
		382052 => x"FF",
		383076 => x"FF",
		384100 => x"FF",
		385124 => x"FF",
		386148 => x"FF",
		387172 => x"FF",
		388196 => x"FF",
		389220 => x"FF",
		390244 => x"FF",
		391268 => x"FF",
		392292 => x"FF",
		393316 => x"FF",
		394340 => x"FF",
		395364 => x"FF",
		396388 => x"FF",
		397412 => x"FF",
		398436 => x"FF",
		399460 => x"FF",
		400484 => x"FF",
		401508 => x"FF",
		402532 => x"FF",
		403556 => x"FF",
		404580 => x"FF",
		405604 => x"FF",
		406628 => x"FF",
		407652 => x"FF",
		408676 => x"FF",
		409700 => x"FF",
		410724 => x"FF",
		411748 => x"FF",
		412772 => x"FF",
		413796 => x"FF",
		414820 => x"FF",
		415844 => x"FF",
		416868 => x"FF",
		417892 => x"FF",
		418916 => x"FF",
		419940 => x"FF",
		420964 => x"FF",
		421988 => x"FF",
		423012 => x"FF",
		424036 => x"FF",
		425060 => x"FF",
		426084 => x"FF",
		427108 => x"FF",
		428132 => x"FF",
		429156 => x"FF",
		430180 => x"FF",
		431204 => x"FF",
		432228 => x"FF",
		433252 => x"FF",
		434276 => x"FF",
		435300 => x"FF",
		436324 => x"FF",
		437348 => x"FF",
		438372 => x"FF",
		439396 => x"FF",
		440420 => x"FF",
		441444 => x"FF",
		442468 => x"FF",
		443492 => x"FF",
		444516 => x"FF",
		445540 => x"FF",
		446564 => x"FF",
		447588 => x"FF",
		448612 => x"FF",
		449636 => x"FF",
		450660 => x"FF",
		451684 => x"FF",
		452708 => x"FF",
		453732 => x"FF",
		454756 => x"FF",
		455780 => x"FF",
		456804 => x"FF",
		457828 => x"FF",
		458852 => x"FF",
		459876 => x"FF",
		460900 => x"FF",
		461924 => x"FF",
		462948 => x"FF",
		463972 => x"FF",
		464996 => x"FF",
		466020 => x"FF",
		467044 => x"FF",
		468068 => x"FF",
		469092 => x"FF",
		19557 => x"FF",
		20581 => x"FF",
		21605 => x"FF",
		22629 => x"FF",
		23653 => x"FF",
		24677 => x"FF",
		25701 => x"FF",
		26725 => x"FF",
		27749 => x"FF",
		28773 => x"FF",
		29797 => x"FF",
		30821 => x"FF",
		31845 => x"FF",
		32869 => x"FF",
		33893 => x"FF",
		34917 => x"FF",
		35941 => x"FF",
		36965 => x"FF",
		37989 => x"FF",
		39013 => x"FF",
		40037 => x"FF",
		41061 => x"FF",
		42085 => x"FF",
		43109 => x"FF",
		44133 => x"FF",
		45157 => x"FF",
		46181 => x"FF",
		47205 => x"FF",
		48229 => x"FF",
		49253 => x"FF",
		50277 => x"FF",
		51301 => x"FF",
		52325 => x"FF",
		53349 => x"FF",
		54373 => x"FF",
		55397 => x"FF",
		56421 => x"FF",
		57445 => x"FF",
		58469 => x"FF",
		59493 => x"FF",
		60517 => x"FF",
		61541 => x"FF",
		62565 => x"FF",
		63589 => x"FF",
		64613 => x"FF",
		65637 => x"FF",
		66661 => x"FF",
		67685 => x"FF",
		68709 => x"FF",
		69733 => x"FF",
		70757 => x"FF",
		71781 => x"FF",
		72805 => x"FF",
		73829 => x"FF",
		74853 => x"FF",
		75877 => x"FF",
		76901 => x"FF",
		77925 => x"FF",
		78949 => x"FF",
		79973 => x"FF",
		80997 => x"FF",
		82021 => x"FF",
		83045 => x"FF",
		84069 => x"FF",
		85093 => x"FF",
		86117 => x"FF",
		87141 => x"FF",
		88165 => x"FF",
		89189 => x"FF",
		90213 => x"FF",
		91237 => x"FF",
		92261 => x"FF",
		93285 => x"FF",
		94309 => x"FF",
		95333 => x"FF",
		96357 => x"FF",
		97381 => x"FF",
		98405 => x"FF",
		99429 => x"FF",
		100453 => x"FF",
		101477 => x"FF",
		102501 => x"FF",
		103525 => x"FF",
		104549 => x"FF",
		105573 => x"FF",
		106597 => x"FF",
		107621 => x"FF",
		108645 => x"FF",
		109669 => x"FF",
		110693 => x"FF",
		111717 => x"FF",
		112741 => x"FF",
		113765 => x"FF",
		114789 => x"FF",
		115813 => x"FF",
		116837 => x"FF",
		117861 => x"FF",
		118885 => x"FF",
		119909 => x"FF",
		120933 => x"FF",
		121957 => x"FF",
		122981 => x"FF",
		124005 => x"FF",
		125029 => x"FF",
		126053 => x"FF",
		127077 => x"FF",
		128101 => x"FF",
		129125 => x"FF",
		130149 => x"FF",
		131173 => x"FF",
		132197 => x"FF",
		133221 => x"FF",
		134245 => x"FF",
		135269 => x"FF",
		136293 => x"FF",
		137317 => x"FF",
		138341 => x"FF",
		139365 => x"FF",
		140389 => x"FF",
		141413 => x"FF",
		142437 => x"FF",
		143461 => x"FF",
		144485 => x"FF",
		145509 => x"FF",
		146533 => x"FF",
		147557 => x"FF",
		148581 => x"FF",
		149605 => x"FF",
		150629 => x"FF",
		151653 => x"FF",
		152677 => x"FF",
		153701 => x"FF",
		154725 => x"FF",
		155749 => x"FF",
		156773 => x"FF",
		157797 => x"FF",
		158821 => x"FF",
		159845 => x"FF",
		160869 => x"FF",
		161893 => x"FF",
		162917 => x"FF",
		163941 => x"FF",
		164965 => x"FF",
		165989 => x"FF",
		167013 => x"FF",
		168037 => x"FF",
		169061 => x"FF",
		170085 => x"FF",
		171109 => x"FF",
		172133 => x"FF",
		173157 => x"FF",
		174181 => x"FF",
		175205 => x"FF",
		176229 => x"FF",
		177253 => x"FF",
		178277 => x"FF",
		179301 => x"FF",
		180325 => x"FF",
		181349 => x"FF",
		182373 => x"FF",
		183397 => x"FF",
		184421 => x"FF",
		185445 => x"FF",
		186469 => x"FF",
		187493 => x"FF",
		188517 => x"FF",
		189541 => x"FF",
		190565 => x"FF",
		191589 => x"FF",
		192613 => x"FF",
		193637 => x"FF",
		194661 => x"FF",
		195685 => x"FF",
		196709 => x"FF",
		197733 => x"FF",
		198757 => x"FF",
		199781 => x"FF",
		200805 => x"FF",
		201829 => x"FF",
		202853 => x"FF",
		203877 => x"FF",
		204901 => x"FF",
		205925 => x"FF",
		206949 => x"FF",
		207973 => x"FF",
		208997 => x"FF",
		210021 => x"FF",
		211045 => x"FF",
		212069 => x"FF",
		213093 => x"FF",
		214117 => x"FF",
		215141 => x"FF",
		216165 => x"FF",
		217189 => x"FF",
		218213 => x"FF",
		219237 => x"FF",
		220261 => x"FF",
		221285 => x"FF",
		222309 => x"FF",
		223333 => x"FF",
		224357 => x"FF",
		225381 => x"FF",
		226405 => x"FF",
		227429 => x"FF",
		228453 => x"FF",
		229477 => x"FF",
		230501 => x"FF",
		231525 => x"FF",
		232549 => x"FF",
		233573 => x"FF",
		234597 => x"FF",
		235621 => x"FF",
		236645 => x"FF",
		237669 => x"FF",
		238693 => x"FF",
		239717 => x"FF",
		240741 => x"FF",
		241765 => x"FF",
		242789 => x"FF",
		243813 => x"FF",
		244837 => x"FF",
		245861 => x"FF",
		246885 => x"FF",
		247909 => x"FF",
		248933 => x"FF",
		249957 => x"FF",
		250981 => x"FF",
		252005 => x"FF",
		253029 => x"FF",
		254053 => x"FF",
		255077 => x"FF",
		256101 => x"FF",
		257125 => x"FF",
		258149 => x"FF",
		259173 => x"FF",
		260197 => x"FF",
		261221 => x"FF",
		262245 => x"FF",
		263269 => x"FF",
		264293 => x"FF",
		265317 => x"FF",
		266341 => x"FF",
		267365 => x"FF",
		268389 => x"FF",
		269413 => x"FF",
		270437 => x"FF",
		271461 => x"FF",
		272485 => x"FF",
		273509 => x"FF",
		274533 => x"FF",
		275557 => x"FF",
		276581 => x"FF",
		277605 => x"FF",
		278629 => x"FF",
		279653 => x"FF",
		280677 => x"FF",
		281701 => x"FF",
		282725 => x"FF",
		283749 => x"FF",
		284773 => x"FF",
		285797 => x"FF",
		286821 => x"FF",
		287845 => x"FF",
		288869 => x"FF",
		289893 => x"FF",
		290917 => x"FF",
		291941 => x"FF",
		292965 => x"FF",
		293989 => x"FF",
		295013 => x"FF",
		296037 => x"FF",
		297061 => x"FF",
		298085 => x"FF",
		299109 => x"FF",
		300133 => x"FF",
		301157 => x"FF",
		302181 => x"FF",
		303205 => x"FF",
		304229 => x"FF",
		305253 => x"FF",
		306277 => x"FF",
		307301 => x"FF",
		308325 => x"FF",
		309349 => x"FF",
		310373 => x"FF",
		311397 => x"FF",
		312421 => x"FF",
		313445 => x"FF",
		314469 => x"FF",
		315493 => x"FF",
		316517 => x"FF",
		317541 => x"FF",
		318565 => x"FF",
		319589 => x"FF",
		320613 => x"FF",
		321637 => x"FF",
		322661 => x"FF",
		323685 => x"FF",
		324709 => x"FF",
		325733 => x"FF",
		326757 => x"FF",
		327781 => x"FF",
		328805 => x"FF",
		329829 => x"FF",
		330853 => x"FF",
		331877 => x"FF",
		332901 => x"FF",
		333925 => x"FF",
		334949 => x"FF",
		335973 => x"FF",
		336997 => x"FF",
		338021 => x"FF",
		339045 => x"FF",
		340069 => x"FF",
		341093 => x"FF",
		342117 => x"FF",
		343141 => x"FF",
		344165 => x"FF",
		345189 => x"FF",
		346213 => x"FF",
		347237 => x"FF",
		348261 => x"FF",
		349285 => x"FF",
		350309 => x"FF",
		351333 => x"FF",
		352357 => x"FF",
		353381 => x"FF",
		354405 => x"FF",
		355429 => x"FF",
		356453 => x"FF",
		357477 => x"FF",
		358501 => x"FF",
		359525 => x"FF",
		360549 => x"FF",
		361573 => x"FF",
		362597 => x"FF",
		363621 => x"FF",
		364645 => x"FF",
		365669 => x"FF",
		366693 => x"FF",
		367717 => x"FF",
		368741 => x"FF",
		369765 => x"FF",
		370789 => x"FF",
		371813 => x"FF",
		372837 => x"FF",
		373861 => x"FF",
		374885 => x"FF",
		375909 => x"FF",
		376933 => x"FF",
		377957 => x"FF",
		378981 => x"FF",
		380005 => x"FF",
		381029 => x"FF",
		382053 => x"FF",
		383077 => x"FF",
		384101 => x"FF",
		385125 => x"FF",
		386149 => x"FF",
		387173 => x"FF",
		388197 => x"FF",
		389221 => x"FF",
		390245 => x"FF",
		391269 => x"FF",
		392293 => x"FF",
		393317 => x"FF",
		394341 => x"FF",
		395365 => x"FF",
		396389 => x"FF",
		397413 => x"FF",
		398437 => x"FF",
		399461 => x"FF",
		400485 => x"FF",
		401509 => x"FF",
		402533 => x"FF",
		403557 => x"FF",
		404581 => x"FF",
		405605 => x"FF",
		406629 => x"FF",
		407653 => x"FF",
		408677 => x"FF",
		409701 => x"FF",
		410725 => x"FF",
		411749 => x"FF",
		412773 => x"FF",
		413797 => x"FF",
		414821 => x"FF",
		415845 => x"FF",
		416869 => x"FF",
		417893 => x"FF",
		418917 => x"FF",
		419941 => x"FF",
		420965 => x"FF",
		421989 => x"FF",
		423013 => x"FF",
		424037 => x"FF",
		425061 => x"FF",
		426085 => x"FF",
		427109 => x"FF",
		428133 => x"FF",
		429157 => x"FF",
		430181 => x"FF",
		431205 => x"FF",
		432229 => x"FF",
		433253 => x"FF",
		434277 => x"FF",
		435301 => x"FF",
		436325 => x"FF",
		437349 => x"FF",
		438373 => x"FF",
		439397 => x"FF",
		440421 => x"FF",
		441445 => x"FF",
		442469 => x"FF",
		443493 => x"FF",
		444517 => x"FF",
		445541 => x"FF",
		446565 => x"FF",
		447589 => x"FF",
		448613 => x"FF",
		449637 => x"FF",
		450661 => x"FF",
		451685 => x"FF",
		452709 => x"FF",
		453733 => x"FF",
		454757 => x"FF",
		455781 => x"FF",
		456805 => x"FF",
		457829 => x"FF",
		458853 => x"FF",
		459877 => x"FF",
		460901 => x"FF",
		461925 => x"FF",
		462949 => x"FF",
		463973 => x"FF",
		464997 => x"FF",
		466021 => x"FF",
		467045 => x"FF",
		468069 => x"FF",
		469093 => x"FF",
		19558 => x"FF",
		20582 => x"FF",
		21606 => x"FF",
		22630 => x"FF",
		23654 => x"FF",
		24678 => x"FF",
		25702 => x"FF",
		26726 => x"FF",
		27750 => x"FF",
		28774 => x"FF",
		29798 => x"FF",
		30822 => x"FF",
		31846 => x"FF",
		32870 => x"FF",
		33894 => x"FF",
		34918 => x"FF",
		35942 => x"FF",
		36966 => x"FF",
		37990 => x"FF",
		39014 => x"FF",
		40038 => x"FF",
		41062 => x"FF",
		42086 => x"FF",
		43110 => x"FF",
		44134 => x"FF",
		45158 => x"FF",
		46182 => x"FF",
		47206 => x"FF",
		48230 => x"FF",
		49254 => x"FF",
		50278 => x"FF",
		51302 => x"FF",
		52326 => x"FF",
		53350 => x"FF",
		54374 => x"FF",
		55398 => x"FF",
		56422 => x"FF",
		57446 => x"FF",
		58470 => x"FF",
		59494 => x"FF",
		60518 => x"FF",
		61542 => x"FF",
		62566 => x"FF",
		63590 => x"FF",
		64614 => x"FF",
		65638 => x"FF",
		66662 => x"FF",
		67686 => x"FF",
		68710 => x"FF",
		69734 => x"FF",
		70758 => x"FF",
		71782 => x"FF",
		72806 => x"FF",
		73830 => x"FF",
		74854 => x"FF",
		75878 => x"FF",
		76902 => x"FF",
		77926 => x"FF",
		78950 => x"FF",
		79974 => x"FF",
		80998 => x"FF",
		82022 => x"FF",
		83046 => x"FF",
		84070 => x"FF",
		85094 => x"FF",
		86118 => x"FF",
		87142 => x"FF",
		88166 => x"FF",
		89190 => x"FF",
		90214 => x"FF",
		91238 => x"FF",
		92262 => x"FF",
		93286 => x"FF",
		94310 => x"FF",
		95334 => x"FF",
		96358 => x"FF",
		97382 => x"FF",
		98406 => x"FF",
		99430 => x"FF",
		100454 => x"FF",
		101478 => x"FF",
		102502 => x"FF",
		103526 => x"FF",
		104550 => x"FF",
		105574 => x"FF",
		106598 => x"FF",
		107622 => x"FF",
		108646 => x"FF",
		109670 => x"FF",
		110694 => x"FF",
		111718 => x"FF",
		112742 => x"FF",
		113766 => x"FF",
		114790 => x"FF",
		115814 => x"FF",
		116838 => x"FF",
		117862 => x"FF",
		118886 => x"FF",
		119910 => x"FF",
		120934 => x"FF",
		121958 => x"FF",
		122982 => x"FF",
		124006 => x"FF",
		125030 => x"FF",
		126054 => x"FF",
		127078 => x"FF",
		128102 => x"FF",
		129126 => x"FF",
		130150 => x"FF",
		131174 => x"FF",
		132198 => x"FF",
		133222 => x"FF",
		134246 => x"FF",
		135270 => x"FF",
		136294 => x"FF",
		137318 => x"FF",
		138342 => x"FF",
		139366 => x"FF",
		140390 => x"FF",
		141414 => x"FF",
		142438 => x"FF",
		143462 => x"FF",
		144486 => x"FF",
		145510 => x"FF",
		146534 => x"FF",
		147558 => x"FF",
		148582 => x"FF",
		149606 => x"FF",
		150630 => x"FF",
		151654 => x"FF",
		152678 => x"FF",
		153702 => x"FF",
		154726 => x"FF",
		155750 => x"FF",
		156774 => x"FF",
		157798 => x"FF",
		158822 => x"FF",
		159846 => x"FF",
		160870 => x"FF",
		161894 => x"FF",
		162918 => x"FF",
		163942 => x"FF",
		164966 => x"FF",
		165990 => x"FF",
		167014 => x"FF",
		168038 => x"FF",
		169062 => x"FF",
		170086 => x"FF",
		171110 => x"FF",
		172134 => x"FF",
		173158 => x"FF",
		174182 => x"FF",
		175206 => x"FF",
		176230 => x"FF",
		177254 => x"FF",
		178278 => x"FF",
		179302 => x"FF",
		180326 => x"FF",
		181350 => x"FF",
		182374 => x"FF",
		183398 => x"FF",
		184422 => x"FF",
		185446 => x"FF",
		186470 => x"FF",
		187494 => x"FF",
		188518 => x"FF",
		189542 => x"FF",
		190566 => x"FF",
		191590 => x"FF",
		192614 => x"FF",
		193638 => x"FF",
		194662 => x"FF",
		195686 => x"FF",
		196710 => x"FF",
		197734 => x"FF",
		198758 => x"FF",
		199782 => x"FF",
		200806 => x"FF",
		201830 => x"FF",
		202854 => x"FF",
		203878 => x"FF",
		204902 => x"FF",
		205926 => x"FF",
		206950 => x"FF",
		207974 => x"FF",
		208998 => x"FF",
		210022 => x"FF",
		211046 => x"FF",
		212070 => x"FF",
		213094 => x"FF",
		214118 => x"FF",
		215142 => x"FF",
		216166 => x"FF",
		217190 => x"FF",
		218214 => x"FF",
		219238 => x"FF",
		220262 => x"FF",
		221286 => x"FF",
		222310 => x"FF",
		223334 => x"FF",
		224358 => x"FF",
		225382 => x"FF",
		226406 => x"FF",
		227430 => x"FF",
		228454 => x"FF",
		229478 => x"FF",
		230502 => x"FF",
		231526 => x"FF",
		232550 => x"FF",
		233574 => x"FF",
		234598 => x"FF",
		235622 => x"FF",
		236646 => x"FF",
		237670 => x"FF",
		238694 => x"FF",
		239718 => x"FF",
		240742 => x"FF",
		241766 => x"FF",
		242790 => x"FF",
		243814 => x"FF",
		244838 => x"FF",
		245862 => x"FF",
		246886 => x"FF",
		247910 => x"FF",
		248934 => x"FF",
		249958 => x"FF",
		250982 => x"FF",
		252006 => x"FF",
		253030 => x"FF",
		254054 => x"FF",
		255078 => x"FF",
		256102 => x"FF",
		257126 => x"FF",
		258150 => x"FF",
		259174 => x"FF",
		260198 => x"FF",
		261222 => x"FF",
		262246 => x"FF",
		263270 => x"FF",
		264294 => x"FF",
		265318 => x"FF",
		266342 => x"FF",
		267366 => x"FF",
		268390 => x"FF",
		269414 => x"FF",
		270438 => x"FF",
		271462 => x"FF",
		272486 => x"FF",
		273510 => x"FF",
		274534 => x"FF",
		275558 => x"FF",
		276582 => x"FF",
		277606 => x"FF",
		278630 => x"FF",
		279654 => x"FF",
		280678 => x"FF",
		281702 => x"FF",
		282726 => x"FF",
		283750 => x"FF",
		284774 => x"FF",
		285798 => x"FF",
		286822 => x"FF",
		287846 => x"FF",
		288870 => x"FF",
		289894 => x"FF",
		290918 => x"FF",
		291942 => x"FF",
		292966 => x"FF",
		293990 => x"FF",
		295014 => x"FF",
		296038 => x"FF",
		297062 => x"FF",
		298086 => x"FF",
		299110 => x"FF",
		300134 => x"FF",
		301158 => x"FF",
		302182 => x"FF",
		303206 => x"FF",
		304230 => x"FF",
		305254 => x"FF",
		306278 => x"FF",
		307302 => x"FF",
		308326 => x"FF",
		309350 => x"FF",
		310374 => x"FF",
		311398 => x"FF",
		312422 => x"FF",
		313446 => x"FF",
		314470 => x"FF",
		315494 => x"FF",
		316518 => x"FF",
		317542 => x"FF",
		318566 => x"FF",
		319590 => x"FF",
		320614 => x"FF",
		321638 => x"FF",
		322662 => x"FF",
		323686 => x"FF",
		324710 => x"FF",
		325734 => x"FF",
		326758 => x"FF",
		327782 => x"FF",
		328806 => x"FF",
		329830 => x"FF",
		330854 => x"FF",
		331878 => x"FF",
		332902 => x"FF",
		333926 => x"FF",
		334950 => x"FF",
		335974 => x"FF",
		336998 => x"FF",
		338022 => x"FF",
		339046 => x"FF",
		340070 => x"FF",
		341094 => x"FF",
		342118 => x"FF",
		343142 => x"FF",
		344166 => x"FF",
		345190 => x"FF",
		346214 => x"FF",
		347238 => x"FF",
		348262 => x"FF",
		349286 => x"FF",
		350310 => x"FF",
		351334 => x"FF",
		352358 => x"FF",
		353382 => x"FF",
		354406 => x"FF",
		355430 => x"FF",
		356454 => x"FF",
		357478 => x"FF",
		358502 => x"FF",
		359526 => x"FF",
		360550 => x"FF",
		361574 => x"FF",
		362598 => x"FF",
		363622 => x"FF",
		364646 => x"FF",
		365670 => x"FF",
		366694 => x"FF",
		367718 => x"FF",
		368742 => x"FF",
		369766 => x"FF",
		370790 => x"FF",
		371814 => x"FF",
		372838 => x"FF",
		373862 => x"FF",
		374886 => x"FF",
		375910 => x"FF",
		376934 => x"FF",
		377958 => x"FF",
		378982 => x"FF",
		380006 => x"FF",
		381030 => x"FF",
		382054 => x"FF",
		383078 => x"FF",
		384102 => x"FF",
		385126 => x"FF",
		386150 => x"FF",
		387174 => x"FF",
		388198 => x"FF",
		389222 => x"FF",
		390246 => x"FF",
		391270 => x"FF",
		392294 => x"FF",
		393318 => x"FF",
		394342 => x"FF",
		395366 => x"FF",
		396390 => x"FF",
		397414 => x"FF",
		398438 => x"FF",
		399462 => x"FF",
		400486 => x"FF",
		401510 => x"FF",
		402534 => x"FF",
		403558 => x"FF",
		404582 => x"FF",
		405606 => x"FF",
		406630 => x"FF",
		407654 => x"FF",
		408678 => x"FF",
		409702 => x"FF",
		410726 => x"FF",
		411750 => x"FF",
		412774 => x"FF",
		413798 => x"FF",
		414822 => x"FF",
		415846 => x"FF",
		416870 => x"FF",
		417894 => x"FF",
		418918 => x"FF",
		419942 => x"FF",
		420966 => x"FF",
		421990 => x"FF",
		423014 => x"FF",
		424038 => x"FF",
		425062 => x"FF",
		426086 => x"FF",
		427110 => x"FF",
		428134 => x"FF",
		429158 => x"FF",
		430182 => x"FF",
		431206 => x"FF",
		432230 => x"FF",
		433254 => x"FF",
		434278 => x"FF",
		435302 => x"FF",
		436326 => x"FF",
		437350 => x"FF",
		438374 => x"FF",
		439398 => x"FF",
		440422 => x"FF",
		441446 => x"FF",
		442470 => x"FF",
		443494 => x"FF",
		444518 => x"FF",
		445542 => x"FF",
		446566 => x"FF",
		447590 => x"FF",
		448614 => x"FF",
		449638 => x"FF",
		450662 => x"FF",
		451686 => x"FF",
		452710 => x"FF",
		453734 => x"FF",
		454758 => x"FF",
		455782 => x"FF",
		456806 => x"FF",
		457830 => x"FF",
		458854 => x"FF",
		459878 => x"FF",
		460902 => x"FF",
		461926 => x"FF",
		462950 => x"FF",
		463974 => x"FF",
		464998 => x"FF",
		466022 => x"FF",
		467046 => x"FF",
		468070 => x"FF",
		469094 => x"FF",
		19559 => x"FF",
		20583 => x"FF",
		21607 => x"FF",
		22631 => x"FF",
		23655 => x"FF",
		24679 => x"FF",
		25703 => x"FF",
		26727 => x"FF",
		27751 => x"FF",
		28775 => x"FF",
		29799 => x"FF",
		30823 => x"FF",
		31847 => x"FF",
		32871 => x"FF",
		33895 => x"FF",
		34919 => x"FF",
		35943 => x"FF",
		36967 => x"FF",
		37991 => x"FF",
		39015 => x"FF",
		40039 => x"FF",
		41063 => x"FF",
		42087 => x"FF",
		43111 => x"FF",
		44135 => x"FF",
		45159 => x"FF",
		46183 => x"FF",
		47207 => x"FF",
		48231 => x"FF",
		49255 => x"FF",
		50279 => x"FF",
		51303 => x"FF",
		52327 => x"FF",
		53351 => x"FF",
		54375 => x"FF",
		55399 => x"FF",
		56423 => x"FF",
		57447 => x"FF",
		58471 => x"FF",
		59495 => x"FF",
		60519 => x"FF",
		61543 => x"FF",
		62567 => x"FF",
		63591 => x"FF",
		64615 => x"FF",
		65639 => x"FF",
		66663 => x"FF",
		67687 => x"FF",
		68711 => x"FF",
		69735 => x"FF",
		70759 => x"FF",
		71783 => x"FF",
		72807 => x"FF",
		73831 => x"FF",
		74855 => x"FF",
		75879 => x"FF",
		76903 => x"FF",
		77927 => x"FF",
		78951 => x"FF",
		79975 => x"FF",
		80999 => x"FF",
		82023 => x"FF",
		83047 => x"FF",
		84071 => x"FF",
		85095 => x"FF",
		86119 => x"FF",
		87143 => x"FF",
		88167 => x"FF",
		89191 => x"FF",
		90215 => x"FF",
		91239 => x"FF",
		92263 => x"FF",
		93287 => x"FF",
		94311 => x"FF",
		95335 => x"FF",
		96359 => x"FF",
		97383 => x"FF",
		98407 => x"FF",
		99431 => x"FF",
		100455 => x"FF",
		101479 => x"FF",
		102503 => x"FF",
		103527 => x"FF",
		104551 => x"FF",
		105575 => x"FF",
		106599 => x"FF",
		107623 => x"FF",
		108647 => x"FF",
		109671 => x"FF",
		110695 => x"FF",
		111719 => x"FF",
		112743 => x"FF",
		113767 => x"FF",
		114791 => x"FF",
		115815 => x"FF",
		116839 => x"FF",
		117863 => x"FF",
		118887 => x"FF",
		119911 => x"FF",
		120935 => x"FF",
		121959 => x"FF",
		122983 => x"FF",
		124007 => x"FF",
		125031 => x"FF",
		126055 => x"FF",
		127079 => x"FF",
		128103 => x"FF",
		129127 => x"FF",
		130151 => x"FF",
		131175 => x"FF",
		132199 => x"FF",
		133223 => x"FF",
		134247 => x"FF",
		135271 => x"FF",
		136295 => x"FF",
		137319 => x"FF",
		138343 => x"FF",
		139367 => x"FF",
		140391 => x"FF",
		141415 => x"FF",
		142439 => x"FF",
		143463 => x"FF",
		144487 => x"FF",
		145511 => x"FF",
		146535 => x"FF",
		147559 => x"FF",
		148583 => x"FF",
		149607 => x"FF",
		150631 => x"FF",
		151655 => x"FF",
		152679 => x"FF",
		153703 => x"FF",
		154727 => x"FF",
		155751 => x"FF",
		156775 => x"FF",
		157799 => x"FF",
		158823 => x"FF",
		159847 => x"FF",
		160871 => x"FF",
		161895 => x"FF",
		162919 => x"FF",
		163943 => x"FF",
		164967 => x"FF",
		165991 => x"FF",
		167015 => x"FF",
		168039 => x"FF",
		169063 => x"FF",
		170087 => x"FF",
		171111 => x"FF",
		172135 => x"FF",
		173159 => x"FF",
		174183 => x"FF",
		175207 => x"FF",
		176231 => x"FF",
		177255 => x"FF",
		178279 => x"FF",
		179303 => x"FF",
		180327 => x"FF",
		181351 => x"FF",
		182375 => x"FF",
		183399 => x"FF",
		184423 => x"FF",
		185447 => x"FF",
		186471 => x"FF",
		187495 => x"FF",
		188519 => x"FF",
		189543 => x"FF",
		190567 => x"FF",
		191591 => x"FF",
		192615 => x"FF",
		193639 => x"FF",
		194663 => x"FF",
		195687 => x"FF",
		196711 => x"FF",
		197735 => x"FF",
		198759 => x"FF",
		199783 => x"FF",
		200807 => x"FF",
		201831 => x"FF",
		202855 => x"FF",
		203879 => x"FF",
		204903 => x"FF",
		205927 => x"FF",
		206951 => x"FF",
		207975 => x"FF",
		208999 => x"FF",
		210023 => x"FF",
		211047 => x"FF",
		212071 => x"FF",
		213095 => x"FF",
		214119 => x"FF",
		215143 => x"FF",
		216167 => x"FF",
		217191 => x"FF",
		218215 => x"FF",
		219239 => x"FF",
		220263 => x"FF",
		221287 => x"FF",
		222311 => x"FF",
		223335 => x"FF",
		224359 => x"FF",
		225383 => x"FF",
		226407 => x"FF",
		227431 => x"FF",
		228455 => x"FF",
		229479 => x"FF",
		230503 => x"FF",
		231527 => x"FF",
		232551 => x"FF",
		233575 => x"FF",
		234599 => x"FF",
		235623 => x"FF",
		236647 => x"FF",
		237671 => x"FF",
		238695 => x"FF",
		239719 => x"FF",
		240743 => x"FF",
		241767 => x"FF",
		242791 => x"FF",
		243815 => x"FF",
		244839 => x"FF",
		245863 => x"FF",
		246887 => x"FF",
		247911 => x"FF",
		248935 => x"FF",
		249959 => x"FF",
		250983 => x"FF",
		252007 => x"FF",
		253031 => x"FF",
		254055 => x"FF",
		255079 => x"FF",
		256103 => x"FF",
		257127 => x"FF",
		258151 => x"FF",
		259175 => x"FF",
		260199 => x"FF",
		261223 => x"FF",
		262247 => x"FF",
		263271 => x"FF",
		264295 => x"FF",
		265319 => x"FF",
		266343 => x"FF",
		267367 => x"FF",
		268391 => x"FF",
		269415 => x"FF",
		270439 => x"FF",
		271463 => x"FF",
		272487 => x"FF",
		273511 => x"FF",
		274535 => x"FF",
		275559 => x"FF",
		276583 => x"FF",
		277607 => x"FF",
		278631 => x"FF",
		279655 => x"FF",
		280679 => x"FF",
		281703 => x"FF",
		282727 => x"FF",
		283751 => x"FF",
		284775 => x"FF",
		285799 => x"FF",
		286823 => x"FF",
		287847 => x"FF",
		288871 => x"FF",
		289895 => x"FF",
		290919 => x"FF",
		291943 => x"FF",
		292967 => x"FF",
		293991 => x"FF",
		295015 => x"FF",
		296039 => x"FF",
		297063 => x"FF",
		298087 => x"FF",
		299111 => x"FF",
		300135 => x"FF",
		301159 => x"FF",
		302183 => x"FF",
		303207 => x"FF",
		304231 => x"FF",
		305255 => x"FF",
		306279 => x"FF",
		307303 => x"FF",
		308327 => x"FF",
		309351 => x"FF",
		310375 => x"FF",
		311399 => x"FF",
		312423 => x"FF",
		313447 => x"FF",
		314471 => x"FF",
		315495 => x"FF",
		316519 => x"FF",
		317543 => x"FF",
		318567 => x"FF",
		319591 => x"FF",
		320615 => x"FF",
		321639 => x"FF",
		322663 => x"FF",
		323687 => x"FF",
		324711 => x"FF",
		325735 => x"FF",
		326759 => x"FF",
		327783 => x"FF",
		328807 => x"FF",
		329831 => x"FF",
		330855 => x"FF",
		331879 => x"FF",
		332903 => x"FF",
		333927 => x"FF",
		334951 => x"FF",
		335975 => x"FF",
		336999 => x"FF",
		338023 => x"FF",
		339047 => x"FF",
		340071 => x"FF",
		341095 => x"FF",
		342119 => x"FF",
		343143 => x"FF",
		344167 => x"FF",
		345191 => x"FF",
		346215 => x"FF",
		347239 => x"FF",
		348263 => x"FF",
		349287 => x"FF",
		350311 => x"FF",
		351335 => x"FF",
		352359 => x"FF",
		353383 => x"FF",
		354407 => x"FF",
		355431 => x"FF",
		356455 => x"FF",
		357479 => x"FF",
		358503 => x"FF",
		359527 => x"FF",
		360551 => x"FF",
		361575 => x"FF",
		362599 => x"FF",
		363623 => x"FF",
		364647 => x"FF",
		365671 => x"FF",
		366695 => x"FF",
		367719 => x"FF",
		368743 => x"FF",
		369767 => x"FF",
		370791 => x"FF",
		371815 => x"FF",
		372839 => x"FF",
		373863 => x"FF",
		374887 => x"FF",
		375911 => x"FF",
		376935 => x"FF",
		377959 => x"FF",
		378983 => x"FF",
		380007 => x"FF",
		381031 => x"FF",
		382055 => x"FF",
		383079 => x"FF",
		384103 => x"FF",
		385127 => x"FF",
		386151 => x"FF",
		387175 => x"FF",
		388199 => x"FF",
		389223 => x"FF",
		390247 => x"FF",
		391271 => x"FF",
		392295 => x"FF",
		393319 => x"FF",
		394343 => x"FF",
		395367 => x"FF",
		396391 => x"FF",
		397415 => x"FF",
		398439 => x"FF",
		399463 => x"FF",
		400487 => x"FF",
		401511 => x"FF",
		402535 => x"FF",
		403559 => x"FF",
		404583 => x"FF",
		405607 => x"FF",
		406631 => x"FF",
		407655 => x"FF",
		408679 => x"FF",
		409703 => x"FF",
		410727 => x"FF",
		411751 => x"FF",
		412775 => x"FF",
		413799 => x"FF",
		414823 => x"FF",
		415847 => x"FF",
		416871 => x"FF",
		417895 => x"FF",
		418919 => x"FF",
		419943 => x"FF",
		420967 => x"FF",
		421991 => x"FF",
		423015 => x"FF",
		424039 => x"FF",
		425063 => x"FF",
		426087 => x"FF",
		427111 => x"FF",
		428135 => x"FF",
		429159 => x"FF",
		430183 => x"FF",
		431207 => x"FF",
		432231 => x"FF",
		433255 => x"FF",
		434279 => x"FF",
		435303 => x"FF",
		436327 => x"FF",
		437351 => x"FF",
		438375 => x"FF",
		439399 => x"FF",
		440423 => x"FF",
		441447 => x"FF",
		442471 => x"FF",
		443495 => x"FF",
		444519 => x"FF",
		445543 => x"FF",
		446567 => x"FF",
		447591 => x"FF",
		448615 => x"FF",
		449639 => x"FF",
		450663 => x"FF",
		451687 => x"FF",
		452711 => x"FF",
		453735 => x"FF",
		454759 => x"FF",
		455783 => x"FF",
		456807 => x"FF",
		457831 => x"FF",
		458855 => x"FF",
		459879 => x"FF",
		460903 => x"FF",
		461927 => x"FF",
		462951 => x"FF",
		463975 => x"FF",
		464999 => x"FF",
		466023 => x"FF",
		467047 => x"FF",
		468071 => x"FF",
		469095 => x"FF",
		19560 => x"FF",
		20584 => x"FF",
		21608 => x"FF",
		22632 => x"FF",
		23656 => x"FF",
		168040 => x"FF",
		169064 => x"FF",
		170088 => x"FF",
		171112 => x"FF",
		172136 => x"FF",
		316520 => x"FF",
		317544 => x"FF",
		318568 => x"FF",
		319592 => x"FF",
		320616 => x"FF",
		465000 => x"FF",
		466024 => x"FF",
		467048 => x"FF",
		468072 => x"FF",
		469096 => x"FF",
		19561 => x"FF",
		20585 => x"FF",
		21609 => x"FF",
		22633 => x"FF",
		23657 => x"FF",
		168041 => x"FF",
		169065 => x"FF",
		170089 => x"FF",
		171113 => x"FF",
		172137 => x"FF",
		316521 => x"FF",
		317545 => x"FF",
		318569 => x"FF",
		319593 => x"FF",
		320617 => x"FF",
		465001 => x"FF",
		466025 => x"FF",
		467049 => x"FF",
		468073 => x"FF",
		469097 => x"FF",
		19562 => x"FF",
		20586 => x"FF",
		21610 => x"FF",
		22634 => x"FF",
		23658 => x"FF",
		168042 => x"FF",
		169066 => x"FF",
		170090 => x"FF",
		171114 => x"FF",
		172138 => x"FF",
		316522 => x"FF",
		317546 => x"FF",
		318570 => x"FF",
		319594 => x"FF",
		320618 => x"FF",
		465002 => x"FF",
		466026 => x"FF",
		467050 => x"FF",
		468074 => x"FF",
		469098 => x"FF",
		19563 => x"FF",
		20587 => x"FF",
		21611 => x"FF",
		22635 => x"FF",
		23659 => x"FF",
		168043 => x"FF",
		169067 => x"FF",
		170091 => x"FF",
		171115 => x"FF",
		172139 => x"FF",
		316523 => x"FF",
		317547 => x"FF",
		318571 => x"FF",
		319595 => x"FF",
		320619 => x"FF",
		465003 => x"FF",
		466027 => x"FF",
		467051 => x"FF",
		468075 => x"FF",
		469099 => x"FF",
		19564 => x"FF",
		20588 => x"FF",
		21612 => x"FF",
		22636 => x"FF",
		23660 => x"FF",
		168044 => x"FF",
		169068 => x"FF",
		170092 => x"FF",
		171116 => x"FF",
		172140 => x"FF",
		316524 => x"FF",
		317548 => x"FF",
		318572 => x"FF",
		319596 => x"FF",
		320620 => x"FF",
		465004 => x"FF",
		466028 => x"FF",
		467052 => x"FF",
		468076 => x"FF",
		469100 => x"FF",
		19565 => x"FF",
		20589 => x"FF",
		21613 => x"FF",
		22637 => x"FF",
		23661 => x"FF",
		168045 => x"FF",
		169069 => x"FF",
		170093 => x"FF",
		171117 => x"FF",
		172141 => x"FF",
		316525 => x"FF",
		317549 => x"FF",
		318573 => x"FF",
		319597 => x"FF",
		320621 => x"FF",
		465005 => x"FF",
		466029 => x"FF",
		467053 => x"FF",
		468077 => x"FF",
		469101 => x"FF",
		19566 => x"FF",
		20590 => x"FF",
		21614 => x"FF",
		22638 => x"FF",
		23662 => x"FF",
		168046 => x"FF",
		169070 => x"FF",
		170094 => x"FF",
		171118 => x"FF",
		172142 => x"FF",
		316526 => x"FF",
		317550 => x"FF",
		318574 => x"FF",
		319598 => x"FF",
		320622 => x"FF",
		465006 => x"FF",
		466030 => x"FF",
		467054 => x"FF",
		468078 => x"FF",
		469102 => x"FF",
		19567 => x"FF",
		20591 => x"FF",
		21615 => x"FF",
		22639 => x"FF",
		23663 => x"FF",
		168047 => x"FF",
		169071 => x"FF",
		170095 => x"FF",
		171119 => x"FF",
		172143 => x"FF",
		316527 => x"FF",
		317551 => x"FF",
		318575 => x"FF",
		319599 => x"FF",
		320623 => x"FF",
		465007 => x"FF",
		466031 => x"FF",
		467055 => x"FF",
		468079 => x"FF",
		469103 => x"FF",
		19568 => x"FF",
		20592 => x"FF",
		21616 => x"FF",
		22640 => x"FF",
		23664 => x"FF",
		168048 => x"FF",
		169072 => x"FF",
		170096 => x"FF",
		171120 => x"FF",
		172144 => x"FF",
		316528 => x"FF",
		317552 => x"FF",
		318576 => x"FF",
		319600 => x"FF",
		320624 => x"FF",
		465008 => x"FF",
		466032 => x"FF",
		467056 => x"FF",
		468080 => x"FF",
		469104 => x"FF",
		19569 => x"FF",
		20593 => x"FF",
		21617 => x"FF",
		22641 => x"FF",
		23665 => x"FF",
		168049 => x"FF",
		169073 => x"FF",
		170097 => x"FF",
		171121 => x"FF",
		172145 => x"FF",
		316529 => x"FF",
		317553 => x"FF",
		318577 => x"FF",
		319601 => x"FF",
		320625 => x"FF",
		465009 => x"FF",
		466033 => x"FF",
		467057 => x"FF",
		468081 => x"FF",
		469105 => x"FF",
		19570 => x"FF",
		20594 => x"FF",
		21618 => x"FF",
		22642 => x"FF",
		23666 => x"FF",
		168050 => x"FF",
		169074 => x"FF",
		170098 => x"FF",
		171122 => x"FF",
		172146 => x"FF",
		316530 => x"FF",
		317554 => x"FF",
		318578 => x"FF",
		319602 => x"FF",
		320626 => x"FF",
		465010 => x"FF",
		466034 => x"FF",
		467058 => x"FF",
		468082 => x"FF",
		469106 => x"FF",
		19571 => x"FF",
		20595 => x"FF",
		21619 => x"FF",
		22643 => x"FF",
		23667 => x"FF",
		168051 => x"FF",
		169075 => x"FF",
		170099 => x"FF",
		171123 => x"FF",
		172147 => x"FF",
		316531 => x"FF",
		317555 => x"FF",
		318579 => x"FF",
		319603 => x"FF",
		320627 => x"FF",
		465011 => x"FF",
		466035 => x"FF",
		467059 => x"FF",
		468083 => x"FF",
		469107 => x"FF",
		19572 => x"FF",
		20596 => x"FF",
		21620 => x"FF",
		22644 => x"FF",
		23668 => x"FF",
		168052 => x"FF",
		169076 => x"FF",
		170100 => x"FF",
		171124 => x"FF",
		172148 => x"FF",
		316532 => x"FF",
		317556 => x"FF",
		318580 => x"FF",
		319604 => x"FF",
		320628 => x"FF",
		465012 => x"FF",
		466036 => x"FF",
		467060 => x"FF",
		468084 => x"FF",
		469108 => x"FF",
		19573 => x"FF",
		20597 => x"FF",
		21621 => x"FF",
		22645 => x"FF",
		23669 => x"FF",
		168053 => x"FF",
		169077 => x"FF",
		170101 => x"FF",
		171125 => x"FF",
		172149 => x"FF",
		316533 => x"FF",
		317557 => x"FF",
		318581 => x"FF",
		319605 => x"FF",
		320629 => x"FF",
		465013 => x"FF",
		466037 => x"FF",
		467061 => x"FF",
		468085 => x"FF",
		469109 => x"FF",
		19574 => x"FF",
		20598 => x"FF",
		21622 => x"FF",
		22646 => x"FF",
		23670 => x"FF",
		168054 => x"FF",
		169078 => x"FF",
		170102 => x"FF",
		171126 => x"FF",
		172150 => x"FF",
		316534 => x"FF",
		317558 => x"FF",
		318582 => x"FF",
		319606 => x"FF",
		320630 => x"FF",
		465014 => x"FF",
		466038 => x"FF",
		467062 => x"FF",
		468086 => x"FF",
		469110 => x"FF",
		19575 => x"FF",
		20599 => x"FF",
		21623 => x"FF",
		22647 => x"FF",
		23671 => x"FF",
		168055 => x"FF",
		169079 => x"FF",
		170103 => x"FF",
		171127 => x"FF",
		172151 => x"FF",
		316535 => x"FF",
		317559 => x"FF",
		318583 => x"FF",
		319607 => x"FF",
		320631 => x"FF",
		465015 => x"FF",
		466039 => x"FF",
		467063 => x"FF",
		468087 => x"FF",
		469111 => x"FF",
		19576 => x"FF",
		20600 => x"FF",
		21624 => x"FF",
		22648 => x"FF",
		23672 => x"FF",
		168056 => x"FF",
		169080 => x"FF",
		170104 => x"FF",
		171128 => x"FF",
		172152 => x"FF",
		316536 => x"FF",
		317560 => x"FF",
		318584 => x"FF",
		319608 => x"FF",
		320632 => x"FF",
		465016 => x"FF",
		466040 => x"FF",
		467064 => x"FF",
		468088 => x"FF",
		469112 => x"FF",
		19577 => x"FF",
		20601 => x"FF",
		21625 => x"FF",
		22649 => x"FF",
		23673 => x"FF",
		168057 => x"FF",
		169081 => x"FF",
		170105 => x"FF",
		171129 => x"FF",
		172153 => x"FF",
		316537 => x"FF",
		317561 => x"FF",
		318585 => x"FF",
		319609 => x"FF",
		320633 => x"FF",
		465017 => x"FF",
		466041 => x"FF",
		467065 => x"FF",
		468089 => x"FF",
		469113 => x"FF",
		19578 => x"FF",
		20602 => x"FF",
		21626 => x"FF",
		22650 => x"FF",
		23674 => x"FF",
		168058 => x"FF",
		169082 => x"FF",
		170106 => x"FF",
		171130 => x"FF",
		172154 => x"FF",
		316538 => x"FF",
		317562 => x"FF",
		318586 => x"FF",
		319610 => x"FF",
		320634 => x"FF",
		465018 => x"FF",
		466042 => x"FF",
		467066 => x"FF",
		468090 => x"FF",
		469114 => x"FF",
		19579 => x"FF",
		20603 => x"FF",
		21627 => x"FF",
		22651 => x"FF",
		23675 => x"FF",
		168059 => x"FF",
		169083 => x"FF",
		170107 => x"FF",
		171131 => x"FF",
		172155 => x"FF",
		316539 => x"FF",
		317563 => x"FF",
		318587 => x"FF",
		319611 => x"FF",
		320635 => x"FF",
		465019 => x"FF",
		466043 => x"FF",
		467067 => x"FF",
		468091 => x"FF",
		469115 => x"FF",
		19580 => x"FF",
		20604 => x"FF",
		21628 => x"FF",
		22652 => x"FF",
		23676 => x"FF",
		168060 => x"FF",
		169084 => x"FF",
		170108 => x"FF",
		171132 => x"FF",
		172156 => x"FF",
		316540 => x"FF",
		317564 => x"FF",
		318588 => x"FF",
		319612 => x"FF",
		320636 => x"FF",
		465020 => x"FF",
		466044 => x"FF",
		467068 => x"FF",
		468092 => x"FF",
		469116 => x"FF",
		19581 => x"FF",
		20605 => x"FF",
		21629 => x"FF",
		22653 => x"FF",
		23677 => x"FF",
		168061 => x"FF",
		169085 => x"FF",
		170109 => x"FF",
		171133 => x"FF",
		172157 => x"FF",
		316541 => x"FF",
		317565 => x"FF",
		318589 => x"FF",
		319613 => x"FF",
		320637 => x"FF",
		465021 => x"FF",
		466045 => x"FF",
		467069 => x"FF",
		468093 => x"FF",
		469117 => x"FF",
		19582 => x"FF",
		20606 => x"FF",
		21630 => x"FF",
		22654 => x"FF",
		23678 => x"FF",
		168062 => x"FF",
		169086 => x"FF",
		170110 => x"FF",
		171134 => x"FF",
		172158 => x"FF",
		316542 => x"FF",
		317566 => x"FF",
		318590 => x"FF",
		319614 => x"FF",
		320638 => x"FF",
		465022 => x"FF",
		466046 => x"FF",
		467070 => x"FF",
		468094 => x"FF",
		469118 => x"FF",
		19583 => x"FF",
		20607 => x"FF",
		21631 => x"FF",
		22655 => x"FF",
		23679 => x"FF",
		168063 => x"FF",
		169087 => x"FF",
		170111 => x"FF",
		171135 => x"FF",
		172159 => x"FF",
		316543 => x"FF",
		317567 => x"FF",
		318591 => x"FF",
		319615 => x"FF",
		320639 => x"FF",
		465023 => x"FF",
		466047 => x"FF",
		467071 => x"FF",
		468095 => x"FF",
		469119 => x"FF",
		19584 => x"FF",
		20608 => x"FF",
		21632 => x"FF",
		22656 => x"FF",
		23680 => x"FF",
		168064 => x"FF",
		169088 => x"FF",
		170112 => x"FF",
		171136 => x"FF",
		172160 => x"FF",
		316544 => x"FF",
		317568 => x"FF",
		318592 => x"FF",
		319616 => x"FF",
		320640 => x"FF",
		465024 => x"FF",
		466048 => x"FF",
		467072 => x"FF",
		468096 => x"FF",
		469120 => x"FF",
		19585 => x"FF",
		20609 => x"FF",
		21633 => x"FF",
		22657 => x"FF",
		23681 => x"FF",
		168065 => x"FF",
		169089 => x"FF",
		170113 => x"FF",
		171137 => x"FF",
		172161 => x"FF",
		316545 => x"FF",
		317569 => x"FF",
		318593 => x"FF",
		319617 => x"FF",
		320641 => x"FF",
		465025 => x"FF",
		466049 => x"FF",
		467073 => x"FF",
		468097 => x"FF",
		469121 => x"FF",
		19586 => x"FF",
		20610 => x"FF",
		21634 => x"FF",
		22658 => x"FF",
		23682 => x"FF",
		168066 => x"FF",
		169090 => x"FF",
		170114 => x"FF",
		171138 => x"FF",
		172162 => x"FF",
		316546 => x"FF",
		317570 => x"FF",
		318594 => x"FF",
		319618 => x"FF",
		320642 => x"FF",
		465026 => x"FF",
		466050 => x"FF",
		467074 => x"FF",
		468098 => x"FF",
		469122 => x"FF",
		19587 => x"FF",
		20611 => x"FF",
		21635 => x"FF",
		22659 => x"FF",
		23683 => x"FF",
		168067 => x"FF",
		169091 => x"FF",
		170115 => x"FF",
		171139 => x"FF",
		172163 => x"FF",
		316547 => x"FF",
		317571 => x"FF",
		318595 => x"FF",
		319619 => x"FF",
		320643 => x"FF",
		465027 => x"FF",
		466051 => x"FF",
		467075 => x"FF",
		468099 => x"FF",
		469123 => x"FF",
		19588 => x"FF",
		20612 => x"FF",
		21636 => x"FF",
		22660 => x"FF",
		23684 => x"FF",
		168068 => x"FF",
		169092 => x"FF",
		170116 => x"FF",
		171140 => x"FF",
		172164 => x"FF",
		316548 => x"FF",
		317572 => x"FF",
		318596 => x"FF",
		319620 => x"FF",
		320644 => x"FF",
		465028 => x"FF",
		466052 => x"FF",
		467076 => x"FF",
		468100 => x"FF",
		469124 => x"FF",
		19589 => x"FF",
		20613 => x"FF",
		21637 => x"FF",
		22661 => x"FF",
		23685 => x"FF",
		168069 => x"FF",
		169093 => x"FF",
		170117 => x"FF",
		171141 => x"FF",
		172165 => x"FF",
		316549 => x"FF",
		317573 => x"FF",
		318597 => x"FF",
		319621 => x"FF",
		320645 => x"FF",
		465029 => x"FF",
		466053 => x"FF",
		467077 => x"FF",
		468101 => x"FF",
		469125 => x"FF",
		19590 => x"FF",
		20614 => x"FF",
		21638 => x"FF",
		22662 => x"FF",
		23686 => x"FF",
		168070 => x"FF",
		169094 => x"FF",
		170118 => x"FF",
		171142 => x"FF",
		172166 => x"FF",
		316550 => x"FF",
		317574 => x"FF",
		318598 => x"FF",
		319622 => x"FF",
		320646 => x"FF",
		465030 => x"FF",
		466054 => x"FF",
		467078 => x"FF",
		468102 => x"FF",
		469126 => x"FF",
		19591 => x"FF",
		20615 => x"FF",
		21639 => x"FF",
		22663 => x"FF",
		23687 => x"FF",
		168071 => x"FF",
		169095 => x"FF",
		170119 => x"FF",
		171143 => x"FF",
		172167 => x"FF",
		316551 => x"FF",
		317575 => x"FF",
		318599 => x"FF",
		319623 => x"FF",
		320647 => x"FF",
		465031 => x"FF",
		466055 => x"FF",
		467079 => x"FF",
		468103 => x"FF",
		469127 => x"FF",
		19592 => x"FF",
		20616 => x"FF",
		21640 => x"FF",
		22664 => x"FF",
		23688 => x"FF",
		168072 => x"FF",
		169096 => x"FF",
		170120 => x"FF",
		171144 => x"FF",
		172168 => x"FF",
		316552 => x"FF",
		317576 => x"FF",
		318600 => x"FF",
		319624 => x"FF",
		320648 => x"FF",
		465032 => x"FF",
		466056 => x"FF",
		467080 => x"FF",
		468104 => x"FF",
		469128 => x"FF",
		19593 => x"FF",
		20617 => x"FF",
		21641 => x"FF",
		22665 => x"FF",
		23689 => x"FF",
		168073 => x"FF",
		169097 => x"FF",
		170121 => x"FF",
		171145 => x"FF",
		172169 => x"FF",
		316553 => x"FF",
		317577 => x"FF",
		318601 => x"FF",
		319625 => x"FF",
		320649 => x"FF",
		465033 => x"FF",
		466057 => x"FF",
		467081 => x"FF",
		468105 => x"FF",
		469129 => x"FF",
		19594 => x"FF",
		20618 => x"FF",
		21642 => x"FF",
		22666 => x"FF",
		23690 => x"FF",
		168074 => x"FF",
		169098 => x"FF",
		170122 => x"FF",
		171146 => x"FF",
		172170 => x"FF",
		316554 => x"FF",
		317578 => x"FF",
		318602 => x"FF",
		319626 => x"FF",
		320650 => x"FF",
		465034 => x"FF",
		466058 => x"FF",
		467082 => x"FF",
		468106 => x"FF",
		469130 => x"FF",
		19595 => x"FF",
		20619 => x"FF",
		21643 => x"FF",
		22667 => x"FF",
		23691 => x"FF",
		168075 => x"FF",
		169099 => x"FF",
		170123 => x"FF",
		171147 => x"FF",
		172171 => x"FF",
		316555 => x"FF",
		317579 => x"FF",
		318603 => x"FF",
		319627 => x"FF",
		320651 => x"FF",
		465035 => x"FF",
		466059 => x"FF",
		467083 => x"FF",
		468107 => x"FF",
		469131 => x"FF",
		19596 => x"FF",
		20620 => x"FF",
		21644 => x"FF",
		22668 => x"FF",
		23692 => x"FF",
		168076 => x"FF",
		169100 => x"FF",
		170124 => x"FF",
		171148 => x"FF",
		172172 => x"FF",
		316556 => x"FF",
		317580 => x"FF",
		318604 => x"FF",
		319628 => x"FF",
		320652 => x"FF",
		465036 => x"FF",
		466060 => x"FF",
		467084 => x"FF",
		468108 => x"FF",
		469132 => x"FF",
		19597 => x"FF",
		20621 => x"FF",
		21645 => x"FF",
		22669 => x"FF",
		23693 => x"FF",
		168077 => x"FF",
		169101 => x"FF",
		170125 => x"FF",
		171149 => x"FF",
		172173 => x"FF",
		316557 => x"FF",
		317581 => x"FF",
		318605 => x"FF",
		319629 => x"FF",
		320653 => x"FF",
		465037 => x"FF",
		466061 => x"FF",
		467085 => x"FF",
		468109 => x"FF",
		469133 => x"FF",
		19598 => x"FF",
		20622 => x"FF",
		21646 => x"FF",
		22670 => x"FF",
		23694 => x"FF",
		168078 => x"FF",
		169102 => x"FF",
		170126 => x"FF",
		171150 => x"FF",
		172174 => x"FF",
		316558 => x"FF",
		317582 => x"FF",
		318606 => x"FF",
		319630 => x"FF",
		320654 => x"FF",
		465038 => x"FF",
		466062 => x"FF",
		467086 => x"FF",
		468110 => x"FF",
		469134 => x"FF",
		19599 => x"FF",
		20623 => x"FF",
		21647 => x"FF",
		22671 => x"FF",
		23695 => x"FF",
		168079 => x"FF",
		169103 => x"FF",
		170127 => x"FF",
		171151 => x"FF",
		172175 => x"FF",
		316559 => x"FF",
		317583 => x"FF",
		318607 => x"FF",
		319631 => x"FF",
		320655 => x"FF",
		465039 => x"FF",
		466063 => x"FF",
		467087 => x"FF",
		468111 => x"FF",
		469135 => x"FF",
		19600 => x"FF",
		20624 => x"FF",
		21648 => x"FF",
		22672 => x"FF",
		23696 => x"FF",
		168080 => x"FF",
		169104 => x"FF",
		170128 => x"FF",
		171152 => x"FF",
		172176 => x"FF",
		316560 => x"FF",
		317584 => x"FF",
		318608 => x"FF",
		319632 => x"FF",
		320656 => x"FF",
		465040 => x"FF",
		466064 => x"FF",
		467088 => x"FF",
		468112 => x"FF",
		469136 => x"FF",
		19601 => x"FF",
		20625 => x"FF",
		21649 => x"FF",
		22673 => x"FF",
		23697 => x"FF",
		168081 => x"FF",
		169105 => x"FF",
		170129 => x"FF",
		171153 => x"FF",
		172177 => x"FF",
		316561 => x"FF",
		317585 => x"FF",
		318609 => x"FF",
		319633 => x"FF",
		320657 => x"FF",
		465041 => x"FF",
		466065 => x"FF",
		467089 => x"FF",
		468113 => x"FF",
		469137 => x"FF",
		19602 => x"FF",
		20626 => x"FF",
		21650 => x"FF",
		22674 => x"FF",
		23698 => x"FF",
		168082 => x"FF",
		169106 => x"FF",
		170130 => x"FF",
		171154 => x"FF",
		172178 => x"FF",
		316562 => x"FF",
		317586 => x"FF",
		318610 => x"FF",
		319634 => x"FF",
		320658 => x"FF",
		465042 => x"FF",
		466066 => x"FF",
		467090 => x"FF",
		468114 => x"FF",
		469138 => x"FF",
		19603 => x"FF",
		20627 => x"FF",
		21651 => x"FF",
		22675 => x"FF",
		23699 => x"FF",
		168083 => x"FF",
		169107 => x"FF",
		170131 => x"FF",
		171155 => x"FF",
		172179 => x"FF",
		316563 => x"FF",
		317587 => x"FF",
		318611 => x"FF",
		319635 => x"FF",
		320659 => x"FF",
		465043 => x"FF",
		466067 => x"FF",
		467091 => x"FF",
		468115 => x"FF",
		469139 => x"FF",
		19604 => x"FF",
		20628 => x"FF",
		21652 => x"FF",
		22676 => x"FF",
		23700 => x"FF",
		168084 => x"FF",
		169108 => x"FF",
		170132 => x"FF",
		171156 => x"FF",
		172180 => x"FF",
		316564 => x"FF",
		317588 => x"FF",
		318612 => x"FF",
		319636 => x"FF",
		320660 => x"FF",
		465044 => x"FF",
		466068 => x"FF",
		467092 => x"FF",
		468116 => x"FF",
		469140 => x"FF",
		19605 => x"FF",
		20629 => x"FF",
		21653 => x"FF",
		22677 => x"FF",
		23701 => x"FF",
		168085 => x"FF",
		169109 => x"FF",
		170133 => x"FF",
		171157 => x"FF",
		172181 => x"FF",
		316565 => x"FF",
		317589 => x"FF",
		318613 => x"FF",
		319637 => x"FF",
		320661 => x"FF",
		465045 => x"FF",
		466069 => x"FF",
		467093 => x"FF",
		468117 => x"FF",
		469141 => x"FF",
		19606 => x"FF",
		20630 => x"FF",
		21654 => x"FF",
		22678 => x"FF",
		23702 => x"FF",
		168086 => x"FF",
		169110 => x"FF",
		170134 => x"FF",
		171158 => x"FF",
		172182 => x"FF",
		316566 => x"FF",
		317590 => x"FF",
		318614 => x"FF",
		319638 => x"FF",
		320662 => x"FF",
		465046 => x"FF",
		466070 => x"FF",
		467094 => x"FF",
		468118 => x"FF",
		469142 => x"FF",
		19607 => x"FF",
		20631 => x"FF",
		21655 => x"FF",
		22679 => x"FF",
		23703 => x"FF",
		168087 => x"FF",
		169111 => x"FF",
		170135 => x"FF",
		171159 => x"FF",
		172183 => x"FF",
		316567 => x"FF",
		317591 => x"FF",
		318615 => x"FF",
		319639 => x"FF",
		320663 => x"FF",
		465047 => x"FF",
		466071 => x"FF",
		467095 => x"FF",
		468119 => x"FF",
		469143 => x"FF",
		19608 => x"FF",
		20632 => x"FF",
		21656 => x"FF",
		22680 => x"FF",
		23704 => x"FF",
		168088 => x"FF",
		169112 => x"FF",
		170136 => x"FF",
		171160 => x"FF",
		172184 => x"FF",
		316568 => x"FF",
		317592 => x"FF",
		318616 => x"FF",
		319640 => x"FF",
		320664 => x"FF",
		465048 => x"FF",
		466072 => x"FF",
		467096 => x"FF",
		468120 => x"FF",
		469144 => x"FF",
		19609 => x"FF",
		20633 => x"FF",
		21657 => x"FF",
		22681 => x"FF",
		23705 => x"FF",
		168089 => x"FF",
		169113 => x"FF",
		170137 => x"FF",
		171161 => x"FF",
		172185 => x"FF",
		316569 => x"FF",
		317593 => x"FF",
		318617 => x"FF",
		319641 => x"FF",
		320665 => x"FF",
		465049 => x"FF",
		466073 => x"FF",
		467097 => x"FF",
		468121 => x"FF",
		469145 => x"FF",
		19610 => x"FF",
		20634 => x"FF",
		21658 => x"FF",
		22682 => x"FF",
		23706 => x"FF",
		168090 => x"FF",
		169114 => x"FF",
		170138 => x"FF",
		171162 => x"FF",
		172186 => x"FF",
		316570 => x"FF",
		317594 => x"FF",
		318618 => x"FF",
		319642 => x"FF",
		320666 => x"FF",
		465050 => x"FF",
		466074 => x"FF",
		467098 => x"FF",
		468122 => x"FF",
		469146 => x"FF",
		19611 => x"FF",
		20635 => x"FF",
		21659 => x"FF",
		22683 => x"FF",
		23707 => x"FF",
		168091 => x"FF",
		169115 => x"FF",
		170139 => x"FF",
		171163 => x"FF",
		172187 => x"FF",
		316571 => x"FF",
		317595 => x"FF",
		318619 => x"FF",
		319643 => x"FF",
		320667 => x"FF",
		465051 => x"FF",
		466075 => x"FF",
		467099 => x"FF",
		468123 => x"FF",
		469147 => x"FF",
		19612 => x"FF",
		20636 => x"FF",
		21660 => x"FF",
		22684 => x"FF",
		23708 => x"FF",
		168092 => x"FF",
		169116 => x"FF",
		170140 => x"FF",
		171164 => x"FF",
		172188 => x"FF",
		316572 => x"FF",
		317596 => x"FF",
		318620 => x"FF",
		319644 => x"FF",
		320668 => x"FF",
		465052 => x"FF",
		466076 => x"FF",
		467100 => x"FF",
		468124 => x"FF",
		469148 => x"FF",
		19613 => x"FF",
		20637 => x"FF",
		21661 => x"FF",
		22685 => x"FF",
		23709 => x"FF",
		168093 => x"FF",
		169117 => x"FF",
		170141 => x"FF",
		171165 => x"FF",
		172189 => x"FF",
		316573 => x"FF",
		317597 => x"FF",
		318621 => x"FF",
		319645 => x"FF",
		320669 => x"FF",
		465053 => x"FF",
		466077 => x"FF",
		467101 => x"FF",
		468125 => x"FF",
		469149 => x"FF",
		19614 => x"FF",
		20638 => x"FF",
		21662 => x"FF",
		22686 => x"FF",
		23710 => x"FF",
		168094 => x"FF",
		169118 => x"FF",
		170142 => x"FF",
		171166 => x"FF",
		172190 => x"FF",
		316574 => x"FF",
		317598 => x"FF",
		318622 => x"FF",
		319646 => x"FF",
		320670 => x"FF",
		465054 => x"FF",
		466078 => x"FF",
		467102 => x"FF",
		468126 => x"FF",
		469150 => x"FF",
		19615 => x"FF",
		20639 => x"FF",
		21663 => x"FF",
		22687 => x"FF",
		23711 => x"FF",
		168095 => x"FF",
		169119 => x"FF",
		170143 => x"FF",
		171167 => x"FF",
		172191 => x"FF",
		316575 => x"FF",
		317599 => x"FF",
		318623 => x"FF",
		319647 => x"FF",
		320671 => x"FF",
		465055 => x"FF",
		466079 => x"FF",
		467103 => x"FF",
		468127 => x"FF",
		469151 => x"FF",
		19616 => x"FF",
		20640 => x"FF",
		21664 => x"FF",
		22688 => x"FF",
		23712 => x"FF",
		168096 => x"FF",
		169120 => x"FF",
		170144 => x"FF",
		171168 => x"FF",
		172192 => x"FF",
		316576 => x"FF",
		317600 => x"FF",
		318624 => x"FF",
		319648 => x"FF",
		320672 => x"FF",
		465056 => x"FF",
		466080 => x"FF",
		467104 => x"FF",
		468128 => x"FF",
		469152 => x"FF",
		19617 => x"FF",
		20641 => x"FF",
		21665 => x"FF",
		22689 => x"FF",
		23713 => x"FF",
		168097 => x"FF",
		169121 => x"FF",
		170145 => x"FF",
		171169 => x"FF",
		172193 => x"FF",
		316577 => x"FF",
		317601 => x"FF",
		318625 => x"FF",
		319649 => x"FF",
		320673 => x"FF",
		465057 => x"FF",
		466081 => x"FF",
		467105 => x"FF",
		468129 => x"FF",
		469153 => x"FF",
		19618 => x"FF",
		20642 => x"FF",
		21666 => x"FF",
		22690 => x"FF",
		23714 => x"FF",
		168098 => x"FF",
		169122 => x"FF",
		170146 => x"FF",
		171170 => x"FF",
		172194 => x"FF",
		316578 => x"FF",
		317602 => x"FF",
		318626 => x"FF",
		319650 => x"FF",
		320674 => x"FF",
		465058 => x"FF",
		466082 => x"FF",
		467106 => x"FF",
		468130 => x"FF",
		469154 => x"FF",
		19619 => x"FF",
		20643 => x"FF",
		21667 => x"FF",
		22691 => x"FF",
		23715 => x"FF",
		168099 => x"FF",
		169123 => x"FF",
		170147 => x"FF",
		171171 => x"FF",
		172195 => x"FF",
		316579 => x"FF",
		317603 => x"FF",
		318627 => x"FF",
		319651 => x"FF",
		320675 => x"FF",
		465059 => x"FF",
		466083 => x"FF",
		467107 => x"FF",
		468131 => x"FF",
		469155 => x"FF",
		19620 => x"FF",
		20644 => x"FF",
		21668 => x"FF",
		22692 => x"FF",
		23716 => x"FF",
		168100 => x"FF",
		169124 => x"FF",
		170148 => x"FF",
		171172 => x"FF",
		172196 => x"FF",
		316580 => x"FF",
		317604 => x"FF",
		318628 => x"FF",
		319652 => x"FF",
		320676 => x"FF",
		465060 => x"FF",
		466084 => x"FF",
		467108 => x"FF",
		468132 => x"FF",
		469156 => x"FF",
		19621 => x"FF",
		20645 => x"FF",
		21669 => x"FF",
		22693 => x"FF",
		23717 => x"FF",
		168101 => x"FF",
		169125 => x"FF",
		170149 => x"FF",
		171173 => x"FF",
		172197 => x"FF",
		316581 => x"FF",
		317605 => x"FF",
		318629 => x"FF",
		319653 => x"FF",
		320677 => x"FF",
		465061 => x"FF",
		466085 => x"FF",
		467109 => x"FF",
		468133 => x"FF",
		469157 => x"FF",
		19622 => x"FF",
		20646 => x"FF",
		21670 => x"FF",
		22694 => x"FF",
		23718 => x"FF",
		168102 => x"FF",
		169126 => x"FF",
		170150 => x"FF",
		171174 => x"FF",
		172198 => x"FF",
		316582 => x"FF",
		317606 => x"FF",
		318630 => x"FF",
		319654 => x"FF",
		320678 => x"FF",
		465062 => x"FF",
		466086 => x"FF",
		467110 => x"FF",
		468134 => x"FF",
		469158 => x"FF",
		19623 => x"FF",
		20647 => x"FF",
		21671 => x"FF",
		22695 => x"FF",
		23719 => x"FF",
		168103 => x"FF",
		169127 => x"FF",
		170151 => x"FF",
		171175 => x"FF",
		172199 => x"FF",
		316583 => x"FF",
		317607 => x"FF",
		318631 => x"FF",
		319655 => x"FF",
		320679 => x"FF",
		465063 => x"FF",
		466087 => x"FF",
		467111 => x"FF",
		468135 => x"FF",
		469159 => x"FF",
		19624 => x"FF",
		20648 => x"FF",
		21672 => x"FF",
		22696 => x"FF",
		23720 => x"FF",
		168104 => x"FF",
		169128 => x"FF",
		170152 => x"FF",
		171176 => x"FF",
		172200 => x"FF",
		316584 => x"FF",
		317608 => x"FF",
		318632 => x"FF",
		319656 => x"FF",
		320680 => x"FF",
		465064 => x"FF",
		466088 => x"FF",
		467112 => x"FF",
		468136 => x"FF",
		469160 => x"FF",
		19625 => x"FF",
		20649 => x"FF",
		21673 => x"FF",
		22697 => x"FF",
		23721 => x"FF",
		168105 => x"FF",
		169129 => x"FF",
		170153 => x"FF",
		171177 => x"FF",
		172201 => x"FF",
		316585 => x"FF",
		317609 => x"FF",
		318633 => x"FF",
		319657 => x"FF",
		320681 => x"FF",
		465065 => x"FF",
		466089 => x"FF",
		467113 => x"FF",
		468137 => x"FF",
		469161 => x"FF",
		19626 => x"FF",
		20650 => x"FF",
		21674 => x"FF",
		22698 => x"FF",
		23722 => x"FF",
		168106 => x"FF",
		169130 => x"FF",
		170154 => x"FF",
		171178 => x"FF",
		172202 => x"FF",
		316586 => x"FF",
		317610 => x"FF",
		318634 => x"FF",
		319658 => x"FF",
		320682 => x"FF",
		465066 => x"FF",
		466090 => x"FF",
		467114 => x"FF",
		468138 => x"FF",
		469162 => x"FF",
		19627 => x"FF",
		20651 => x"FF",
		21675 => x"FF",
		22699 => x"FF",
		23723 => x"FF",
		168107 => x"FF",
		169131 => x"FF",
		170155 => x"FF",
		171179 => x"FF",
		172203 => x"FF",
		316587 => x"FF",
		317611 => x"FF",
		318635 => x"FF",
		319659 => x"FF",
		320683 => x"FF",
		465067 => x"FF",
		466091 => x"FF",
		467115 => x"FF",
		468139 => x"FF",
		469163 => x"FF",
		19628 => x"FF",
		20652 => x"FF",
		21676 => x"FF",
		22700 => x"FF",
		23724 => x"FF",
		168108 => x"FF",
		169132 => x"FF",
		170156 => x"FF",
		171180 => x"FF",
		172204 => x"FF",
		316588 => x"FF",
		317612 => x"FF",
		318636 => x"FF",
		319660 => x"FF",
		320684 => x"FF",
		465068 => x"FF",
		466092 => x"FF",
		467116 => x"FF",
		468140 => x"FF",
		469164 => x"FF",
		19629 => x"FF",
		20653 => x"FF",
		21677 => x"FF",
		22701 => x"FF",
		23725 => x"FF",
		168109 => x"FF",
		169133 => x"FF",
		170157 => x"FF",
		171181 => x"FF",
		172205 => x"FF",
		316589 => x"FF",
		317613 => x"FF",
		318637 => x"FF",
		319661 => x"FF",
		320685 => x"FF",
		465069 => x"FF",
		466093 => x"FF",
		467117 => x"FF",
		468141 => x"FF",
		469165 => x"FF",
		19630 => x"FF",
		20654 => x"FF",
		21678 => x"FF",
		22702 => x"FF",
		23726 => x"FF",
		168110 => x"FF",
		169134 => x"FF",
		170158 => x"FF",
		171182 => x"FF",
		172206 => x"FF",
		316590 => x"FF",
		317614 => x"FF",
		318638 => x"FF",
		319662 => x"FF",
		320686 => x"FF",
		465070 => x"FF",
		466094 => x"FF",
		467118 => x"FF",
		468142 => x"FF",
		469166 => x"FF",
		19631 => x"FF",
		20655 => x"FF",
		21679 => x"FF",
		22703 => x"FF",
		23727 => x"FF",
		168111 => x"FF",
		169135 => x"FF",
		170159 => x"FF",
		171183 => x"FF",
		172207 => x"FF",
		316591 => x"FF",
		317615 => x"FF",
		318639 => x"FF",
		319663 => x"FF",
		320687 => x"FF",
		465071 => x"FF",
		466095 => x"FF",
		467119 => x"FF",
		468143 => x"FF",
		469167 => x"FF",
		19632 => x"FF",
		20656 => x"FF",
		21680 => x"FF",
		22704 => x"FF",
		23728 => x"FF",
		168112 => x"FF",
		169136 => x"FF",
		170160 => x"FF",
		171184 => x"FF",
		172208 => x"FF",
		316592 => x"FF",
		317616 => x"FF",
		318640 => x"FF",
		319664 => x"FF",
		320688 => x"FF",
		465072 => x"FF",
		466096 => x"FF",
		467120 => x"FF",
		468144 => x"FF",
		469168 => x"FF",
		19633 => x"FF",
		20657 => x"FF",
		21681 => x"FF",
		22705 => x"FF",
		23729 => x"FF",
		168113 => x"FF",
		169137 => x"FF",
		170161 => x"FF",
		171185 => x"FF",
		172209 => x"FF",
		316593 => x"FF",
		317617 => x"FF",
		318641 => x"FF",
		319665 => x"FF",
		320689 => x"FF",
		465073 => x"FF",
		466097 => x"FF",
		467121 => x"FF",
		468145 => x"FF",
		469169 => x"FF",
		19634 => x"FF",
		20658 => x"FF",
		21682 => x"FF",
		22706 => x"FF",
		23730 => x"FF",
		168114 => x"FF",
		169138 => x"FF",
		170162 => x"FF",
		171186 => x"FF",
		172210 => x"FF",
		316594 => x"FF",
		317618 => x"FF",
		318642 => x"FF",
		319666 => x"FF",
		320690 => x"FF",
		465074 => x"FF",
		466098 => x"FF",
		467122 => x"FF",
		468146 => x"FF",
		469170 => x"FF",
		19635 => x"FF",
		20659 => x"FF",
		21683 => x"FF",
		22707 => x"FF",
		23731 => x"FF",
		168115 => x"FF",
		169139 => x"FF",
		170163 => x"FF",
		171187 => x"FF",
		172211 => x"FF",
		316595 => x"FF",
		317619 => x"FF",
		318643 => x"FF",
		319667 => x"FF",
		320691 => x"FF",
		465075 => x"FF",
		466099 => x"FF",
		467123 => x"FF",
		468147 => x"FF",
		469171 => x"FF",
		19636 => x"FF",
		20660 => x"FF",
		21684 => x"FF",
		22708 => x"FF",
		23732 => x"FF",
		168116 => x"FF",
		169140 => x"FF",
		170164 => x"FF",
		171188 => x"FF",
		172212 => x"FF",
		316596 => x"FF",
		317620 => x"FF",
		318644 => x"FF",
		319668 => x"FF",
		320692 => x"FF",
		465076 => x"FF",
		466100 => x"FF",
		467124 => x"FF",
		468148 => x"FF",
		469172 => x"FF",
		19637 => x"FF",
		20661 => x"FF",
		21685 => x"FF",
		22709 => x"FF",
		23733 => x"FF",
		168117 => x"FF",
		169141 => x"FF",
		170165 => x"FF",
		171189 => x"FF",
		172213 => x"FF",
		316597 => x"FF",
		317621 => x"FF",
		318645 => x"FF",
		319669 => x"FF",
		320693 => x"FF",
		465077 => x"FF",
		466101 => x"FF",
		467125 => x"FF",
		468149 => x"FF",
		469173 => x"FF",
		19638 => x"FF",
		20662 => x"FF",
		21686 => x"FF",
		22710 => x"FF",
		23734 => x"FF",
		168118 => x"FF",
		169142 => x"FF",
		170166 => x"FF",
		171190 => x"FF",
		172214 => x"FF",
		316598 => x"FF",
		317622 => x"FF",
		318646 => x"FF",
		319670 => x"FF",
		320694 => x"FF",
		465078 => x"FF",
		466102 => x"FF",
		467126 => x"FF",
		468150 => x"FF",
		469174 => x"FF",
		19639 => x"FF",
		20663 => x"FF",
		21687 => x"FF",
		22711 => x"FF",
		23735 => x"FF",
		168119 => x"FF",
		169143 => x"FF",
		170167 => x"FF",
		171191 => x"FF",
		172215 => x"FF",
		316599 => x"FF",
		317623 => x"FF",
		318647 => x"FF",
		319671 => x"FF",
		320695 => x"FF",
		465079 => x"FF",
		466103 => x"FF",
		467127 => x"FF",
		468151 => x"FF",
		469175 => x"FF",
		19640 => x"FF",
		20664 => x"FF",
		21688 => x"FF",
		22712 => x"FF",
		23736 => x"FF",
		168120 => x"FF",
		169144 => x"FF",
		170168 => x"FF",
		171192 => x"FF",
		172216 => x"FF",
		316600 => x"FF",
		317624 => x"FF",
		318648 => x"FF",
		319672 => x"FF",
		320696 => x"FF",
		465080 => x"FF",
		466104 => x"FF",
		467128 => x"FF",
		468152 => x"FF",
		469176 => x"FF",
		19641 => x"FF",
		20665 => x"FF",
		21689 => x"FF",
		22713 => x"FF",
		23737 => x"FF",
		168121 => x"FF",
		169145 => x"FF",
		170169 => x"FF",
		171193 => x"FF",
		172217 => x"FF",
		316601 => x"FF",
		317625 => x"FF",
		318649 => x"FF",
		319673 => x"FF",
		320697 => x"FF",
		465081 => x"FF",
		466105 => x"FF",
		467129 => x"FF",
		468153 => x"FF",
		469177 => x"FF",
		19642 => x"FF",
		20666 => x"FF",
		21690 => x"FF",
		22714 => x"FF",
		23738 => x"FF",
		168122 => x"FF",
		169146 => x"FF",
		170170 => x"FF",
		171194 => x"FF",
		172218 => x"FF",
		316602 => x"FF",
		317626 => x"FF",
		318650 => x"FF",
		319674 => x"FF",
		320698 => x"FF",
		465082 => x"FF",
		466106 => x"FF",
		467130 => x"FF",
		468154 => x"FF",
		469178 => x"FF",
		19643 => x"FF",
		20667 => x"FF",
		21691 => x"FF",
		22715 => x"FF",
		23739 => x"FF",
		168123 => x"FF",
		169147 => x"FF",
		170171 => x"FF",
		171195 => x"FF",
		172219 => x"FF",
		316603 => x"FF",
		317627 => x"FF",
		318651 => x"FF",
		319675 => x"FF",
		320699 => x"FF",
		465083 => x"FF",
		466107 => x"FF",
		467131 => x"FF",
		468155 => x"FF",
		469179 => x"FF",
		19644 => x"FF",
		20668 => x"FF",
		21692 => x"FF",
		22716 => x"FF",
		23740 => x"FF",
		168124 => x"FF",
		169148 => x"FF",
		170172 => x"FF",
		171196 => x"FF",
		172220 => x"FF",
		316604 => x"FF",
		317628 => x"FF",
		318652 => x"FF",
		319676 => x"FF",
		320700 => x"FF",
		465084 => x"FF",
		466108 => x"FF",
		467132 => x"FF",
		468156 => x"FF",
		469180 => x"FF",
		19645 => x"FF",
		20669 => x"FF",
		21693 => x"FF",
		22717 => x"FF",
		23741 => x"FF",
		168125 => x"FF",
		169149 => x"FF",
		170173 => x"FF",
		171197 => x"FF",
		172221 => x"FF",
		316605 => x"FF",
		317629 => x"FF",
		318653 => x"FF",
		319677 => x"FF",
		320701 => x"FF",
		465085 => x"FF",
		466109 => x"FF",
		467133 => x"FF",
		468157 => x"FF",
		469181 => x"FF",
		19646 => x"FF",
		20670 => x"FF",
		21694 => x"FF",
		22718 => x"FF",
		23742 => x"FF",
		168126 => x"FF",
		169150 => x"FF",
		170174 => x"FF",
		171198 => x"FF",
		172222 => x"FF",
		316606 => x"FF",
		317630 => x"FF",
		318654 => x"FF",
		319678 => x"FF",
		320702 => x"FF",
		465086 => x"FF",
		466110 => x"FF",
		467134 => x"FF",
		468158 => x"FF",
		469182 => x"FF",
		19647 => x"FF",
		20671 => x"FF",
		21695 => x"FF",
		22719 => x"FF",
		23743 => x"FF",
		168127 => x"FF",
		169151 => x"FF",
		170175 => x"FF",
		171199 => x"FF",
		172223 => x"FF",
		316607 => x"FF",
		317631 => x"FF",
		318655 => x"FF",
		319679 => x"FF",
		320703 => x"FF",
		465087 => x"FF",
		466111 => x"FF",
		467135 => x"FF",
		468159 => x"FF",
		469183 => x"FF",
		19648 => x"FF",
		20672 => x"FF",
		21696 => x"FF",
		22720 => x"FF",
		23744 => x"FF",
		168128 => x"FF",
		169152 => x"FF",
		170176 => x"FF",
		171200 => x"FF",
		172224 => x"FF",
		316608 => x"FF",
		317632 => x"FF",
		318656 => x"FF",
		319680 => x"FF",
		320704 => x"FF",
		465088 => x"FF",
		466112 => x"FF",
		467136 => x"FF",
		468160 => x"FF",
		469184 => x"FF",
		19649 => x"FF",
		20673 => x"FF",
		21697 => x"FF",
		22721 => x"FF",
		23745 => x"FF",
		168129 => x"FF",
		169153 => x"FF",
		170177 => x"FF",
		171201 => x"FF",
		172225 => x"FF",
		316609 => x"FF",
		317633 => x"FF",
		318657 => x"FF",
		319681 => x"FF",
		320705 => x"FF",
		465089 => x"FF",
		466113 => x"FF",
		467137 => x"FF",
		468161 => x"FF",
		469185 => x"FF",
		19650 => x"FF",
		20674 => x"FF",
		21698 => x"FF",
		22722 => x"FF",
		23746 => x"FF",
		168130 => x"FF",
		169154 => x"FF",
		170178 => x"FF",
		171202 => x"FF",
		172226 => x"FF",
		316610 => x"FF",
		317634 => x"FF",
		318658 => x"FF",
		319682 => x"FF",
		320706 => x"FF",
		465090 => x"FF",
		466114 => x"FF",
		467138 => x"FF",
		468162 => x"FF",
		469186 => x"FF",
		19651 => x"FF",
		20675 => x"FF",
		21699 => x"FF",
		22723 => x"FF",
		23747 => x"FF",
		168131 => x"FF",
		169155 => x"FF",
		170179 => x"FF",
		171203 => x"FF",
		172227 => x"FF",
		316611 => x"FF",
		317635 => x"FF",
		318659 => x"FF",
		319683 => x"FF",
		320707 => x"FF",
		465091 => x"FF",
		466115 => x"FF",
		467139 => x"FF",
		468163 => x"FF",
		469187 => x"FF",
		19652 => x"FF",
		20676 => x"FF",
		21700 => x"FF",
		22724 => x"FF",
		23748 => x"FF",
		168132 => x"FF",
		169156 => x"FF",
		170180 => x"FF",
		171204 => x"FF",
		172228 => x"FF",
		316612 => x"FF",
		317636 => x"FF",
		318660 => x"FF",
		319684 => x"FF",
		320708 => x"FF",
		465092 => x"FF",
		466116 => x"FF",
		467140 => x"FF",
		468164 => x"FF",
		469188 => x"FF",
		19653 => x"FF",
		20677 => x"FF",
		21701 => x"FF",
		22725 => x"FF",
		23749 => x"FF",
		168133 => x"FF",
		169157 => x"FF",
		170181 => x"FF",
		171205 => x"FF",
		172229 => x"FF",
		316613 => x"FF",
		317637 => x"FF",
		318661 => x"FF",
		319685 => x"FF",
		320709 => x"FF",
		465093 => x"FF",
		466117 => x"FF",
		467141 => x"FF",
		468165 => x"FF",
		469189 => x"FF",
		19654 => x"FF",
		20678 => x"FF",
		21702 => x"FF",
		22726 => x"FF",
		23750 => x"FF",
		168134 => x"FF",
		169158 => x"FF",
		170182 => x"FF",
		171206 => x"FF",
		172230 => x"FF",
		316614 => x"FF",
		317638 => x"FF",
		318662 => x"FF",
		319686 => x"FF",
		320710 => x"FF",
		465094 => x"FF",
		466118 => x"FF",
		467142 => x"FF",
		468166 => x"FF",
		469190 => x"FF",
		19655 => x"FF",
		20679 => x"FF",
		21703 => x"FF",
		22727 => x"FF",
		23751 => x"FF",
		168135 => x"FF",
		169159 => x"FF",
		170183 => x"FF",
		171207 => x"FF",
		172231 => x"FF",
		316615 => x"FF",
		317639 => x"FF",
		318663 => x"FF",
		319687 => x"FF",
		320711 => x"FF",
		465095 => x"FF",
		466119 => x"FF",
		467143 => x"FF",
		468167 => x"FF",
		469191 => x"FF",
		19656 => x"FF",
		20680 => x"FF",
		21704 => x"FF",
		22728 => x"FF",
		23752 => x"FF",
		168136 => x"FF",
		169160 => x"FF",
		170184 => x"FF",
		171208 => x"FF",
		172232 => x"FF",
		316616 => x"FF",
		317640 => x"FF",
		318664 => x"FF",
		319688 => x"FF",
		320712 => x"FF",
		465096 => x"FF",
		466120 => x"FF",
		467144 => x"FF",
		468168 => x"FF",
		469192 => x"FF",
		19657 => x"FF",
		20681 => x"FF",
		21705 => x"FF",
		22729 => x"FF",
		23753 => x"FF",
		168137 => x"FF",
		169161 => x"FF",
		170185 => x"FF",
		171209 => x"FF",
		172233 => x"FF",
		316617 => x"FF",
		317641 => x"FF",
		318665 => x"FF",
		319689 => x"FF",
		320713 => x"FF",
		465097 => x"FF",
		466121 => x"FF",
		467145 => x"FF",
		468169 => x"FF",
		469193 => x"FF",
		19658 => x"FF",
		20682 => x"FF",
		21706 => x"FF",
		22730 => x"FF",
		23754 => x"FF",
		168138 => x"FF",
		169162 => x"FF",
		170186 => x"FF",
		171210 => x"FF",
		172234 => x"FF",
		316618 => x"FF",
		317642 => x"FF",
		318666 => x"FF",
		319690 => x"FF",
		320714 => x"FF",
		465098 => x"FF",
		466122 => x"FF",
		467146 => x"FF",
		468170 => x"FF",
		469194 => x"FF",
		19659 => x"FF",
		20683 => x"FF",
		21707 => x"FF",
		22731 => x"FF",
		23755 => x"FF",
		168139 => x"FF",
		169163 => x"FF",
		170187 => x"FF",
		171211 => x"FF",
		172235 => x"FF",
		316619 => x"FF",
		317643 => x"FF",
		318667 => x"FF",
		319691 => x"FF",
		320715 => x"FF",
		465099 => x"FF",
		466123 => x"FF",
		467147 => x"FF",
		468171 => x"FF",
		469195 => x"FF",
		19660 => x"FF",
		20684 => x"FF",
		21708 => x"FF",
		22732 => x"FF",
		23756 => x"FF",
		168140 => x"FF",
		169164 => x"FF",
		170188 => x"FF",
		171212 => x"FF",
		172236 => x"FF",
		316620 => x"FF",
		317644 => x"FF",
		318668 => x"FF",
		319692 => x"FF",
		320716 => x"FF",
		465100 => x"FF",
		466124 => x"FF",
		467148 => x"FF",
		468172 => x"FF",
		469196 => x"FF",
		19661 => x"FF",
		20685 => x"FF",
		21709 => x"FF",
		22733 => x"FF",
		23757 => x"FF",
		168141 => x"FF",
		169165 => x"FF",
		170189 => x"FF",
		171213 => x"FF",
		172237 => x"FF",
		316621 => x"FF",
		317645 => x"FF",
		318669 => x"FF",
		319693 => x"FF",
		320717 => x"FF",
		465101 => x"FF",
		466125 => x"FF",
		467149 => x"FF",
		468173 => x"FF",
		469197 => x"FF",
		19662 => x"FF",
		20686 => x"FF",
		21710 => x"FF",
		22734 => x"FF",
		23758 => x"FF",
		168142 => x"FF",
		169166 => x"FF",
		170190 => x"FF",
		171214 => x"FF",
		172238 => x"FF",
		316622 => x"FF",
		317646 => x"FF",
		318670 => x"FF",
		319694 => x"FF",
		320718 => x"FF",
		465102 => x"FF",
		466126 => x"FF",
		467150 => x"FF",
		468174 => x"FF",
		469198 => x"FF",
		19663 => x"FF",
		20687 => x"FF",
		21711 => x"FF",
		22735 => x"FF",
		23759 => x"FF",
		168143 => x"FF",
		169167 => x"FF",
		170191 => x"FF",
		171215 => x"FF",
		172239 => x"FF",
		316623 => x"FF",
		317647 => x"FF",
		318671 => x"FF",
		319695 => x"FF",
		320719 => x"FF",
		465103 => x"FF",
		466127 => x"FF",
		467151 => x"FF",
		468175 => x"FF",
		469199 => x"FF",
		19664 => x"FF",
		20688 => x"FF",
		21712 => x"FF",
		22736 => x"FF",
		23760 => x"FF",
		168144 => x"FF",
		169168 => x"FF",
		170192 => x"FF",
		171216 => x"FF",
		172240 => x"FF",
		316624 => x"FF",
		317648 => x"FF",
		318672 => x"FF",
		319696 => x"FF",
		320720 => x"FF",
		465104 => x"FF",
		466128 => x"FF",
		467152 => x"FF",
		468176 => x"FF",
		469200 => x"FF",
		19665 => x"FF",
		20689 => x"FF",
		21713 => x"FF",
		22737 => x"FF",
		23761 => x"FF",
		168145 => x"FF",
		169169 => x"FF",
		170193 => x"FF",
		171217 => x"FF",
		172241 => x"FF",
		316625 => x"FF",
		317649 => x"FF",
		318673 => x"FF",
		319697 => x"FF",
		320721 => x"FF",
		465105 => x"FF",
		466129 => x"FF",
		467153 => x"FF",
		468177 => x"FF",
		469201 => x"FF",
		19666 => x"FF",
		20690 => x"FF",
		21714 => x"FF",
		22738 => x"FF",
		23762 => x"FF",
		168146 => x"FF",
		169170 => x"FF",
		170194 => x"FF",
		171218 => x"FF",
		172242 => x"FF",
		316626 => x"FF",
		317650 => x"FF",
		318674 => x"FF",
		319698 => x"FF",
		320722 => x"FF",
		465106 => x"FF",
		466130 => x"FF",
		467154 => x"FF",
		468178 => x"FF",
		469202 => x"FF",
		19667 => x"FF",
		20691 => x"FF",
		21715 => x"FF",
		22739 => x"FF",
		23763 => x"FF",
		168147 => x"FF",
		169171 => x"FF",
		170195 => x"FF",
		171219 => x"FF",
		172243 => x"FF",
		316627 => x"FF",
		317651 => x"FF",
		318675 => x"FF",
		319699 => x"FF",
		320723 => x"FF",
		465107 => x"FF",
		466131 => x"FF",
		467155 => x"FF",
		468179 => x"FF",
		469203 => x"FF",
		19668 => x"FF",
		20692 => x"FF",
		21716 => x"FF",
		22740 => x"FF",
		23764 => x"FF",
		168148 => x"FF",
		169172 => x"FF",
		170196 => x"FF",
		171220 => x"FF",
		172244 => x"FF",
		316628 => x"FF",
		317652 => x"FF",
		318676 => x"FF",
		319700 => x"FF",
		320724 => x"FF",
		465108 => x"FF",
		466132 => x"FF",
		467156 => x"FF",
		468180 => x"FF",
		469204 => x"FF",
		19669 => x"FF",
		20693 => x"FF",
		21717 => x"FF",
		22741 => x"FF",
		23765 => x"FF",
		168149 => x"FF",
		169173 => x"FF",
		170197 => x"FF",
		171221 => x"FF",
		172245 => x"FF",
		316629 => x"FF",
		317653 => x"FF",
		318677 => x"FF",
		319701 => x"FF",
		320725 => x"FF",
		465109 => x"FF",
		466133 => x"FF",
		467157 => x"FF",
		468181 => x"FF",
		469205 => x"FF",
		19670 => x"FF",
		20694 => x"FF",
		21718 => x"FF",
		22742 => x"FF",
		23766 => x"FF",
		168150 => x"FF",
		169174 => x"FF",
		170198 => x"FF",
		171222 => x"FF",
		172246 => x"FF",
		316630 => x"FF",
		317654 => x"FF",
		318678 => x"FF",
		319702 => x"FF",
		320726 => x"FF",
		465110 => x"FF",
		466134 => x"FF",
		467158 => x"FF",
		468182 => x"FF",
		469206 => x"FF",
		19671 => x"FF",
		20695 => x"FF",
		21719 => x"FF",
		22743 => x"FF",
		23767 => x"FF",
		168151 => x"FF",
		169175 => x"FF",
		170199 => x"FF",
		171223 => x"FF",
		172247 => x"FF",
		316631 => x"FF",
		317655 => x"FF",
		318679 => x"FF",
		319703 => x"FF",
		320727 => x"FF",
		465111 => x"FF",
		466135 => x"FF",
		467159 => x"FF",
		468183 => x"FF",
		469207 => x"FF",
		19672 => x"FF",
		20696 => x"FF",
		21720 => x"FF",
		22744 => x"FF",
		23768 => x"FF",
		168152 => x"FF",
		169176 => x"FF",
		170200 => x"FF",
		171224 => x"FF",
		172248 => x"FF",
		316632 => x"FF",
		317656 => x"FF",
		318680 => x"FF",
		319704 => x"FF",
		320728 => x"FF",
		465112 => x"FF",
		466136 => x"FF",
		467160 => x"FF",
		468184 => x"FF",
		469208 => x"FF",
		19673 => x"FF",
		20697 => x"FF",
		21721 => x"FF",
		22745 => x"FF",
		23769 => x"FF",
		168153 => x"FF",
		169177 => x"FF",
		170201 => x"FF",
		171225 => x"FF",
		172249 => x"FF",
		316633 => x"FF",
		317657 => x"FF",
		318681 => x"FF",
		319705 => x"FF",
		320729 => x"FF",
		465113 => x"FF",
		466137 => x"FF",
		467161 => x"FF",
		468185 => x"FF",
		469209 => x"FF",
		19674 => x"FF",
		20698 => x"FF",
		21722 => x"FF",
		22746 => x"FF",
		23770 => x"FF",
		168154 => x"FF",
		169178 => x"FF",
		170202 => x"FF",
		171226 => x"FF",
		172250 => x"FF",
		316634 => x"FF",
		317658 => x"FF",
		318682 => x"FF",
		319706 => x"FF",
		320730 => x"FF",
		465114 => x"FF",
		466138 => x"FF",
		467162 => x"FF",
		468186 => x"FF",
		469210 => x"FF",
		19675 => x"FF",
		20699 => x"FF",
		21723 => x"FF",
		22747 => x"FF",
		23771 => x"FF",
		168155 => x"FF",
		169179 => x"FF",
		170203 => x"FF",
		171227 => x"FF",
		172251 => x"FF",
		316635 => x"FF",
		317659 => x"FF",
		318683 => x"FF",
		319707 => x"FF",
		320731 => x"FF",
		465115 => x"FF",
		466139 => x"FF",
		467163 => x"FF",
		468187 => x"FF",
		469211 => x"FF",
		19676 => x"FF",
		20700 => x"FF",
		21724 => x"FF",
		22748 => x"FF",
		23772 => x"FF",
		168156 => x"FF",
		169180 => x"FF",
		170204 => x"FF",
		171228 => x"FF",
		172252 => x"FF",
		316636 => x"FF",
		317660 => x"FF",
		318684 => x"FF",
		319708 => x"FF",
		320732 => x"FF",
		465116 => x"FF",
		466140 => x"FF",
		467164 => x"FF",
		468188 => x"FF",
		469212 => x"FF",
		19677 => x"FF",
		20701 => x"FF",
		21725 => x"FF",
		22749 => x"FF",
		23773 => x"FF",
		168157 => x"FF",
		169181 => x"FF",
		170205 => x"FF",
		171229 => x"FF",
		172253 => x"FF",
		316637 => x"FF",
		317661 => x"FF",
		318685 => x"FF",
		319709 => x"FF",
		320733 => x"FF",
		465117 => x"FF",
		466141 => x"FF",
		467165 => x"FF",
		468189 => x"FF",
		469213 => x"FF",
		19678 => x"FF",
		20702 => x"FF",
		21726 => x"FF",
		22750 => x"FF",
		23774 => x"FF",
		168158 => x"FF",
		169182 => x"FF",
		170206 => x"FF",
		171230 => x"FF",
		172254 => x"FF",
		316638 => x"FF",
		317662 => x"FF",
		318686 => x"FF",
		319710 => x"FF",
		320734 => x"FF",
		465118 => x"FF",
		466142 => x"FF",
		467166 => x"FF",
		468190 => x"FF",
		469214 => x"FF",
		19679 => x"FF",
		20703 => x"FF",
		21727 => x"FF",
		22751 => x"FF",
		23775 => x"FF",
		168159 => x"FF",
		169183 => x"FF",
		170207 => x"FF",
		171231 => x"FF",
		172255 => x"FF",
		316639 => x"FF",
		317663 => x"FF",
		318687 => x"FF",
		319711 => x"FF",
		320735 => x"FF",
		465119 => x"FF",
		466143 => x"FF",
		467167 => x"FF",
		468191 => x"FF",
		469215 => x"FF",
		19680 => x"FF",
		20704 => x"FF",
		21728 => x"FF",
		22752 => x"FF",
		23776 => x"FF",
		168160 => x"FF",
		169184 => x"FF",
		170208 => x"FF",
		171232 => x"FF",
		172256 => x"FF",
		316640 => x"FF",
		317664 => x"FF",
		318688 => x"FF",
		319712 => x"FF",
		320736 => x"FF",
		465120 => x"FF",
		466144 => x"FF",
		467168 => x"FF",
		468192 => x"FF",
		469216 => x"FF",
		19681 => x"FF",
		20705 => x"FF",
		21729 => x"FF",
		22753 => x"FF",
		23777 => x"FF",
		168161 => x"FF",
		169185 => x"FF",
		170209 => x"FF",
		171233 => x"FF",
		172257 => x"FF",
		316641 => x"FF",
		317665 => x"FF",
		318689 => x"FF",
		319713 => x"FF",
		320737 => x"FF",
		465121 => x"FF",
		466145 => x"FF",
		467169 => x"FF",
		468193 => x"FF",
		469217 => x"FF",
		19682 => x"FF",
		20706 => x"FF",
		21730 => x"FF",
		22754 => x"FF",
		23778 => x"FF",
		168162 => x"FF",
		169186 => x"FF",
		170210 => x"FF",
		171234 => x"FF",
		172258 => x"FF",
		316642 => x"FF",
		317666 => x"FF",
		318690 => x"FF",
		319714 => x"FF",
		320738 => x"FF",
		465122 => x"FF",
		466146 => x"FF",
		467170 => x"FF",
		468194 => x"FF",
		469218 => x"FF",
		19683 => x"FF",
		20707 => x"FF",
		21731 => x"FF",
		22755 => x"FF",
		23779 => x"FF",
		168163 => x"FF",
		169187 => x"FF",
		170211 => x"FF",
		171235 => x"FF",
		172259 => x"FF",
		316643 => x"FF",
		317667 => x"FF",
		318691 => x"FF",
		319715 => x"FF",
		320739 => x"FF",
		465123 => x"FF",
		466147 => x"FF",
		467171 => x"FF",
		468195 => x"FF",
		469219 => x"FF",
		19684 => x"FF",
		20708 => x"FF",
		21732 => x"FF",
		22756 => x"FF",
		23780 => x"FF",
		168164 => x"FF",
		169188 => x"FF",
		170212 => x"FF",
		171236 => x"FF",
		172260 => x"FF",
		316644 => x"FF",
		317668 => x"FF",
		318692 => x"FF",
		319716 => x"FF",
		320740 => x"FF",
		465124 => x"FF",
		466148 => x"FF",
		467172 => x"FF",
		468196 => x"FF",
		469220 => x"FF",
		19685 => x"FF",
		20709 => x"FF",
		21733 => x"FF",
		22757 => x"FF",
		23781 => x"FF",
		168165 => x"FF",
		169189 => x"FF",
		170213 => x"FF",
		171237 => x"FF",
		172261 => x"FF",
		316645 => x"FF",
		317669 => x"FF",
		318693 => x"FF",
		319717 => x"FF",
		320741 => x"FF",
		465125 => x"FF",
		466149 => x"FF",
		467173 => x"FF",
		468197 => x"FF",
		469221 => x"FF",
		19686 => x"FF",
		20710 => x"FF",
		21734 => x"FF",
		22758 => x"FF",
		23782 => x"FF",
		168166 => x"FF",
		169190 => x"FF",
		170214 => x"FF",
		171238 => x"FF",
		172262 => x"FF",
		316646 => x"FF",
		317670 => x"FF",
		318694 => x"FF",
		319718 => x"FF",
		320742 => x"FF",
		465126 => x"FF",
		466150 => x"FF",
		467174 => x"FF",
		468198 => x"FF",
		469222 => x"FF",
		19687 => x"FF",
		20711 => x"FF",
		21735 => x"FF",
		22759 => x"FF",
		23783 => x"FF",
		168167 => x"FF",
		169191 => x"FF",
		170215 => x"FF",
		171239 => x"FF",
		172263 => x"FF",
		316647 => x"FF",
		317671 => x"FF",
		318695 => x"FF",
		319719 => x"FF",
		320743 => x"FF",
		465127 => x"FF",
		466151 => x"FF",
		467175 => x"FF",
		468199 => x"FF",
		469223 => x"FF",
		19688 => x"FF",
		20712 => x"FF",
		21736 => x"FF",
		22760 => x"FF",
		23784 => x"FF",
		168168 => x"FF",
		169192 => x"FF",
		170216 => x"FF",
		171240 => x"FF",
		172264 => x"FF",
		316648 => x"FF",
		317672 => x"FF",
		318696 => x"FF",
		319720 => x"FF",
		320744 => x"FF",
		465128 => x"FF",
		466152 => x"FF",
		467176 => x"FF",
		468200 => x"FF",
		469224 => x"FF",
		19689 => x"FF",
		20713 => x"FF",
		21737 => x"FF",
		22761 => x"FF",
		23785 => x"FF",
		168169 => x"FF",
		169193 => x"FF",
		170217 => x"FF",
		171241 => x"FF",
		172265 => x"FF",
		316649 => x"FF",
		317673 => x"FF",
		318697 => x"FF",
		319721 => x"FF",
		320745 => x"FF",
		465129 => x"FF",
		466153 => x"FF",
		467177 => x"FF",
		468201 => x"FF",
		469225 => x"FF",
		19690 => x"FF",
		20714 => x"FF",
		21738 => x"FF",
		22762 => x"FF",
		23786 => x"FF",
		168170 => x"FF",
		169194 => x"FF",
		170218 => x"FF",
		171242 => x"FF",
		172266 => x"FF",
		316650 => x"FF",
		317674 => x"FF",
		318698 => x"FF",
		319722 => x"FF",
		320746 => x"FF",
		465130 => x"FF",
		466154 => x"FF",
		467178 => x"FF",
		468202 => x"FF",
		469226 => x"FF",
		19691 => x"FF",
		20715 => x"FF",
		21739 => x"FF",
		22763 => x"FF",
		23787 => x"FF",
		168171 => x"FF",
		169195 => x"FF",
		170219 => x"FF",
		171243 => x"FF",
		172267 => x"FF",
		316651 => x"FF",
		317675 => x"FF",
		318699 => x"FF",
		319723 => x"FF",
		320747 => x"FF",
		465131 => x"FF",
		466155 => x"FF",
		467179 => x"FF",
		468203 => x"FF",
		469227 => x"FF",
		19692 => x"FF",
		20716 => x"FF",
		21740 => x"FF",
		22764 => x"FF",
		23788 => x"FF",
		168172 => x"FF",
		169196 => x"FF",
		170220 => x"FF",
		171244 => x"FF",
		172268 => x"FF",
		316652 => x"FF",
		317676 => x"FF",
		318700 => x"FF",
		319724 => x"FF",
		320748 => x"FF",
		465132 => x"FF",
		466156 => x"FF",
		467180 => x"FF",
		468204 => x"FF",
		469228 => x"FF",
		19693 => x"FF",
		20717 => x"FF",
		21741 => x"FF",
		22765 => x"FF",
		23789 => x"FF",
		168173 => x"FF",
		169197 => x"FF",
		170221 => x"FF",
		171245 => x"FF",
		172269 => x"FF",
		316653 => x"FF",
		317677 => x"FF",
		318701 => x"FF",
		319725 => x"FF",
		320749 => x"FF",
		465133 => x"FF",
		466157 => x"FF",
		467181 => x"FF",
		468205 => x"FF",
		469229 => x"FF",
		19694 => x"FF",
		20718 => x"FF",
		21742 => x"FF",
		22766 => x"FF",
		23790 => x"FF",
		168174 => x"FF",
		169198 => x"FF",
		170222 => x"FF",
		171246 => x"FF",
		172270 => x"FF",
		316654 => x"FF",
		317678 => x"FF",
		318702 => x"FF",
		319726 => x"FF",
		320750 => x"FF",
		465134 => x"FF",
		466158 => x"FF",
		467182 => x"FF",
		468206 => x"FF",
		469230 => x"FF",
		19695 => x"FF",
		20719 => x"FF",
		21743 => x"FF",
		22767 => x"FF",
		23791 => x"FF",
		168175 => x"FF",
		169199 => x"FF",
		170223 => x"FF",
		171247 => x"FF",
		172271 => x"FF",
		316655 => x"FF",
		317679 => x"FF",
		318703 => x"FF",
		319727 => x"FF",
		320751 => x"FF",
		465135 => x"FF",
		466159 => x"FF",
		467183 => x"FF",
		468207 => x"FF",
		469231 => x"FF",
		19696 => x"FF",
		20720 => x"FF",
		21744 => x"FF",
		22768 => x"FF",
		23792 => x"FF",
		168176 => x"FF",
		169200 => x"FF",
		170224 => x"FF",
		171248 => x"FF",
		172272 => x"FF",
		316656 => x"FF",
		317680 => x"FF",
		318704 => x"FF",
		319728 => x"FF",
		320752 => x"FF",
		465136 => x"FF",
		466160 => x"FF",
		467184 => x"FF",
		468208 => x"FF",
		469232 => x"FF",
		19697 => x"FF",
		20721 => x"FF",
		21745 => x"FF",
		22769 => x"FF",
		23793 => x"FF",
		168177 => x"FF",
		169201 => x"FF",
		170225 => x"FF",
		171249 => x"FF",
		172273 => x"FF",
		316657 => x"FF",
		317681 => x"FF",
		318705 => x"FF",
		319729 => x"FF",
		320753 => x"FF",
		465137 => x"FF",
		466161 => x"FF",
		467185 => x"FF",
		468209 => x"FF",
		469233 => x"FF",
		19698 => x"FF",
		20722 => x"FF",
		21746 => x"FF",
		22770 => x"FF",
		23794 => x"FF",
		168178 => x"FF",
		169202 => x"FF",
		170226 => x"FF",
		171250 => x"FF",
		172274 => x"FF",
		316658 => x"FF",
		317682 => x"FF",
		318706 => x"FF",
		319730 => x"FF",
		320754 => x"FF",
		465138 => x"FF",
		466162 => x"FF",
		467186 => x"FF",
		468210 => x"FF",
		469234 => x"FF",
		19699 => x"FF",
		20723 => x"FF",
		21747 => x"FF",
		22771 => x"FF",
		23795 => x"FF",
		168179 => x"FF",
		169203 => x"FF",
		170227 => x"FF",
		171251 => x"FF",
		172275 => x"FF",
		316659 => x"FF",
		317683 => x"FF",
		318707 => x"FF",
		319731 => x"FF",
		320755 => x"FF",
		465139 => x"FF",
		466163 => x"FF",
		467187 => x"FF",
		468211 => x"FF",
		469235 => x"FF",
		19700 => x"FF",
		20724 => x"FF",
		21748 => x"FF",
		22772 => x"FF",
		23796 => x"FF",
		24820 => x"FF",
		25844 => x"FF",
		26868 => x"FF",
		27892 => x"FF",
		28916 => x"FF",
		29940 => x"FF",
		30964 => x"FF",
		31988 => x"FF",
		33012 => x"FF",
		34036 => x"FF",
		35060 => x"FF",
		36084 => x"FF",
		37108 => x"FF",
		38132 => x"FF",
		39156 => x"FF",
		40180 => x"FF",
		41204 => x"FF",
		42228 => x"FF",
		43252 => x"FF",
		44276 => x"FF",
		45300 => x"FF",
		46324 => x"FF",
		47348 => x"FF",
		48372 => x"FF",
		49396 => x"FF",
		50420 => x"FF",
		51444 => x"FF",
		52468 => x"FF",
		53492 => x"FF",
		54516 => x"FF",
		55540 => x"FF",
		56564 => x"FF",
		57588 => x"FF",
		58612 => x"FF",
		59636 => x"FF",
		60660 => x"FF",
		61684 => x"FF",
		62708 => x"FF",
		63732 => x"FF",
		64756 => x"FF",
		65780 => x"FF",
		66804 => x"FF",
		67828 => x"FF",
		68852 => x"FF",
		69876 => x"FF",
		70900 => x"FF",
		71924 => x"FF",
		72948 => x"FF",
		73972 => x"FF",
		74996 => x"FF",
		76020 => x"FF",
		77044 => x"FF",
		78068 => x"FF",
		79092 => x"FF",
		80116 => x"FF",
		81140 => x"FF",
		82164 => x"FF",
		83188 => x"FF",
		84212 => x"FF",
		85236 => x"FF",
		86260 => x"FF",
		87284 => x"FF",
		88308 => x"FF",
		89332 => x"FF",
		90356 => x"FF",
		91380 => x"FF",
		92404 => x"FF",
		93428 => x"FF",
		94452 => x"FF",
		95476 => x"FF",
		96500 => x"FF",
		97524 => x"FF",
		98548 => x"FF",
		99572 => x"FF",
		100596 => x"FF",
		101620 => x"FF",
		102644 => x"FF",
		103668 => x"FF",
		104692 => x"FF",
		105716 => x"FF",
		106740 => x"FF",
		107764 => x"FF",
		108788 => x"FF",
		109812 => x"FF",
		110836 => x"FF",
		111860 => x"FF",
		112884 => x"FF",
		113908 => x"FF",
		114932 => x"FF",
		115956 => x"FF",
		116980 => x"FF",
		118004 => x"FF",
		119028 => x"FF",
		120052 => x"FF",
		121076 => x"FF",
		122100 => x"FF",
		123124 => x"FF",
		124148 => x"FF",
		125172 => x"FF",
		126196 => x"FF",
		127220 => x"FF",
		128244 => x"FF",
		129268 => x"FF",
		130292 => x"FF",
		131316 => x"FF",
		132340 => x"FF",
		133364 => x"FF",
		134388 => x"FF",
		135412 => x"FF",
		136436 => x"FF",
		137460 => x"FF",
		138484 => x"FF",
		139508 => x"FF",
		140532 => x"FF",
		141556 => x"FF",
		142580 => x"FF",
		143604 => x"FF",
		144628 => x"FF",
		145652 => x"FF",
		146676 => x"FF",
		147700 => x"FF",
		148724 => x"FF",
		149748 => x"FF",
		150772 => x"FF",
		151796 => x"FF",
		152820 => x"FF",
		153844 => x"FF",
		154868 => x"FF",
		155892 => x"FF",
		156916 => x"FF",
		157940 => x"FF",
		158964 => x"FF",
		159988 => x"FF",
		161012 => x"FF",
		162036 => x"FF",
		163060 => x"FF",
		164084 => x"FF",
		165108 => x"FF",
		166132 => x"FF",
		167156 => x"FF",
		168180 => x"FF",
		169204 => x"FF",
		170228 => x"FF",
		171252 => x"FF",
		172276 => x"FF",
		173300 => x"FF",
		174324 => x"FF",
		175348 => x"FF",
		176372 => x"FF",
		177396 => x"FF",
		178420 => x"FF",
		179444 => x"FF",
		180468 => x"FF",
		181492 => x"FF",
		182516 => x"FF",
		183540 => x"FF",
		184564 => x"FF",
		185588 => x"FF",
		186612 => x"FF",
		187636 => x"FF",
		188660 => x"FF",
		189684 => x"FF",
		190708 => x"FF",
		191732 => x"FF",
		192756 => x"FF",
		193780 => x"FF",
		194804 => x"FF",
		195828 => x"FF",
		196852 => x"FF",
		197876 => x"FF",
		198900 => x"FF",
		199924 => x"FF",
		200948 => x"FF",
		201972 => x"FF",
		202996 => x"FF",
		204020 => x"FF",
		205044 => x"FF",
		206068 => x"FF",
		207092 => x"FF",
		208116 => x"FF",
		209140 => x"FF",
		210164 => x"FF",
		211188 => x"FF",
		212212 => x"FF",
		213236 => x"FF",
		214260 => x"FF",
		215284 => x"FF",
		216308 => x"FF",
		217332 => x"FF",
		218356 => x"FF",
		219380 => x"FF",
		220404 => x"FF",
		221428 => x"FF",
		222452 => x"FF",
		223476 => x"FF",
		224500 => x"FF",
		225524 => x"FF",
		226548 => x"FF",
		227572 => x"FF",
		228596 => x"FF",
		229620 => x"FF",
		230644 => x"FF",
		231668 => x"FF",
		232692 => x"FF",
		233716 => x"FF",
		234740 => x"FF",
		235764 => x"FF",
		236788 => x"FF",
		237812 => x"FF",
		238836 => x"FF",
		239860 => x"FF",
		240884 => x"FF",
		241908 => x"FF",
		242932 => x"FF",
		243956 => x"FF",
		244980 => x"FF",
		246004 => x"FF",
		247028 => x"FF",
		248052 => x"FF",
		249076 => x"FF",
		250100 => x"FF",
		251124 => x"FF",
		252148 => x"FF",
		253172 => x"FF",
		254196 => x"FF",
		255220 => x"FF",
		256244 => x"FF",
		257268 => x"FF",
		258292 => x"FF",
		259316 => x"FF",
		260340 => x"FF",
		261364 => x"FF",
		262388 => x"FF",
		263412 => x"FF",
		264436 => x"FF",
		265460 => x"FF",
		266484 => x"FF",
		267508 => x"FF",
		268532 => x"FF",
		269556 => x"FF",
		270580 => x"FF",
		271604 => x"FF",
		272628 => x"FF",
		273652 => x"FF",
		274676 => x"FF",
		275700 => x"FF",
		276724 => x"FF",
		277748 => x"FF",
		278772 => x"FF",
		279796 => x"FF",
		280820 => x"FF",
		281844 => x"FF",
		282868 => x"FF",
		283892 => x"FF",
		284916 => x"FF",
		285940 => x"FF",
		286964 => x"FF",
		287988 => x"FF",
		289012 => x"FF",
		290036 => x"FF",
		291060 => x"FF",
		292084 => x"FF",
		293108 => x"FF",
		294132 => x"FF",
		295156 => x"FF",
		296180 => x"FF",
		297204 => x"FF",
		298228 => x"FF",
		299252 => x"FF",
		300276 => x"FF",
		301300 => x"FF",
		302324 => x"FF",
		303348 => x"FF",
		304372 => x"FF",
		305396 => x"FF",
		306420 => x"FF",
		307444 => x"FF",
		308468 => x"FF",
		309492 => x"FF",
		310516 => x"FF",
		311540 => x"FF",
		312564 => x"FF",
		313588 => x"FF",
		314612 => x"FF",
		315636 => x"FF",
		316660 => x"FF",
		317684 => x"FF",
		318708 => x"FF",
		319732 => x"FF",
		320756 => x"FF",
		321780 => x"FF",
		322804 => x"FF",
		323828 => x"FF",
		324852 => x"FF",
		325876 => x"FF",
		326900 => x"FF",
		327924 => x"FF",
		328948 => x"FF",
		329972 => x"FF",
		330996 => x"FF",
		332020 => x"FF",
		333044 => x"FF",
		334068 => x"FF",
		335092 => x"FF",
		336116 => x"FF",
		337140 => x"FF",
		338164 => x"FF",
		339188 => x"FF",
		340212 => x"FF",
		341236 => x"FF",
		342260 => x"FF",
		343284 => x"FF",
		344308 => x"FF",
		345332 => x"FF",
		346356 => x"FF",
		347380 => x"FF",
		348404 => x"FF",
		349428 => x"FF",
		350452 => x"FF",
		351476 => x"FF",
		352500 => x"FF",
		353524 => x"FF",
		354548 => x"FF",
		355572 => x"FF",
		356596 => x"FF",
		357620 => x"FF",
		358644 => x"FF",
		359668 => x"FF",
		360692 => x"FF",
		361716 => x"FF",
		362740 => x"FF",
		363764 => x"FF",
		364788 => x"FF",
		365812 => x"FF",
		366836 => x"FF",
		367860 => x"FF",
		368884 => x"FF",
		369908 => x"FF",
		370932 => x"FF",
		371956 => x"FF",
		372980 => x"FF",
		374004 => x"FF",
		375028 => x"FF",
		376052 => x"FF",
		377076 => x"FF",
		378100 => x"FF",
		379124 => x"FF",
		380148 => x"FF",
		381172 => x"FF",
		382196 => x"FF",
		383220 => x"FF",
		384244 => x"FF",
		385268 => x"FF",
		386292 => x"FF",
		387316 => x"FF",
		388340 => x"FF",
		389364 => x"FF",
		390388 => x"FF",
		391412 => x"FF",
		392436 => x"FF",
		393460 => x"FF",
		394484 => x"FF",
		395508 => x"FF",
		396532 => x"FF",
		397556 => x"FF",
		398580 => x"FF",
		399604 => x"FF",
		400628 => x"FF",
		401652 => x"FF",
		402676 => x"FF",
		403700 => x"FF",
		404724 => x"FF",
		405748 => x"FF",
		406772 => x"FF",
		407796 => x"FF",
		408820 => x"FF",
		409844 => x"FF",
		410868 => x"FF",
		411892 => x"FF",
		412916 => x"FF",
		413940 => x"FF",
		414964 => x"FF",
		415988 => x"FF",
		417012 => x"FF",
		418036 => x"FF",
		419060 => x"FF",
		420084 => x"FF",
		421108 => x"FF",
		422132 => x"FF",
		423156 => x"FF",
		424180 => x"FF",
		425204 => x"FF",
		426228 => x"FF",
		427252 => x"FF",
		428276 => x"FF",
		429300 => x"FF",
		430324 => x"FF",
		431348 => x"FF",
		432372 => x"FF",
		433396 => x"FF",
		434420 => x"FF",
		435444 => x"FF",
		436468 => x"FF",
		437492 => x"FF",
		438516 => x"FF",
		439540 => x"FF",
		440564 => x"FF",
		441588 => x"FF",
		442612 => x"FF",
		443636 => x"FF",
		444660 => x"FF",
		445684 => x"FF",
		446708 => x"FF",
		447732 => x"FF",
		448756 => x"FF",
		449780 => x"FF",
		450804 => x"FF",
		451828 => x"FF",
		452852 => x"FF",
		453876 => x"FF",
		454900 => x"FF",
		455924 => x"FF",
		456948 => x"FF",
		457972 => x"FF",
		458996 => x"FF",
		460020 => x"FF",
		461044 => x"FF",
		462068 => x"FF",
		463092 => x"FF",
		464116 => x"FF",
		465140 => x"FF",
		466164 => x"FF",
		467188 => x"FF",
		468212 => x"FF",
		469236 => x"FF",
		19701 => x"FF",
		20725 => x"FF",
		21749 => x"FF",
		22773 => x"FF",
		23797 => x"FF",
		24821 => x"FF",
		25845 => x"FF",
		26869 => x"FF",
		27893 => x"FF",
		28917 => x"FF",
		29941 => x"FF",
		30965 => x"FF",
		31989 => x"FF",
		33013 => x"FF",
		34037 => x"FF",
		35061 => x"FF",
		36085 => x"FF",
		37109 => x"FF",
		38133 => x"FF",
		39157 => x"FF",
		40181 => x"FF",
		41205 => x"FF",
		42229 => x"FF",
		43253 => x"FF",
		44277 => x"FF",
		45301 => x"FF",
		46325 => x"FF",
		47349 => x"FF",
		48373 => x"FF",
		49397 => x"FF",
		50421 => x"FF",
		51445 => x"FF",
		52469 => x"FF",
		53493 => x"FF",
		54517 => x"FF",
		55541 => x"FF",
		56565 => x"FF",
		57589 => x"FF",
		58613 => x"FF",
		59637 => x"FF",
		60661 => x"FF",
		61685 => x"FF",
		62709 => x"FF",
		63733 => x"FF",
		64757 => x"FF",
		65781 => x"FF",
		66805 => x"FF",
		67829 => x"FF",
		68853 => x"FF",
		69877 => x"FF",
		70901 => x"FF",
		71925 => x"FF",
		72949 => x"FF",
		73973 => x"FF",
		74997 => x"FF",
		76021 => x"FF",
		77045 => x"FF",
		78069 => x"FF",
		79093 => x"FF",
		80117 => x"FF",
		81141 => x"FF",
		82165 => x"FF",
		83189 => x"FF",
		84213 => x"FF",
		85237 => x"FF",
		86261 => x"FF",
		87285 => x"FF",
		88309 => x"FF",
		89333 => x"FF",
		90357 => x"FF",
		91381 => x"FF",
		92405 => x"FF",
		93429 => x"FF",
		94453 => x"FF",
		95477 => x"FF",
		96501 => x"FF",
		97525 => x"FF",
		98549 => x"FF",
		99573 => x"FF",
		100597 => x"FF",
		101621 => x"FF",
		102645 => x"FF",
		103669 => x"FF",
		104693 => x"FF",
		105717 => x"FF",
		106741 => x"FF",
		107765 => x"FF",
		108789 => x"FF",
		109813 => x"FF",
		110837 => x"FF",
		111861 => x"FF",
		112885 => x"FF",
		113909 => x"FF",
		114933 => x"FF",
		115957 => x"FF",
		116981 => x"FF",
		118005 => x"FF",
		119029 => x"FF",
		120053 => x"FF",
		121077 => x"FF",
		122101 => x"FF",
		123125 => x"FF",
		124149 => x"FF",
		125173 => x"FF",
		126197 => x"FF",
		127221 => x"FF",
		128245 => x"FF",
		129269 => x"FF",
		130293 => x"FF",
		131317 => x"FF",
		132341 => x"FF",
		133365 => x"FF",
		134389 => x"FF",
		135413 => x"FF",
		136437 => x"FF",
		137461 => x"FF",
		138485 => x"FF",
		139509 => x"FF",
		140533 => x"FF",
		141557 => x"FF",
		142581 => x"FF",
		143605 => x"FF",
		144629 => x"FF",
		145653 => x"FF",
		146677 => x"FF",
		147701 => x"FF",
		148725 => x"FF",
		149749 => x"FF",
		150773 => x"FF",
		151797 => x"FF",
		152821 => x"FF",
		153845 => x"FF",
		154869 => x"FF",
		155893 => x"FF",
		156917 => x"FF",
		157941 => x"FF",
		158965 => x"FF",
		159989 => x"FF",
		161013 => x"FF",
		162037 => x"FF",
		163061 => x"FF",
		164085 => x"FF",
		165109 => x"FF",
		166133 => x"FF",
		167157 => x"FF",
		168181 => x"FF",
		169205 => x"FF",
		170229 => x"FF",
		171253 => x"FF",
		172277 => x"FF",
		173301 => x"FF",
		174325 => x"FF",
		175349 => x"FF",
		176373 => x"FF",
		177397 => x"FF",
		178421 => x"FF",
		179445 => x"FF",
		180469 => x"FF",
		181493 => x"FF",
		182517 => x"FF",
		183541 => x"FF",
		184565 => x"FF",
		185589 => x"FF",
		186613 => x"FF",
		187637 => x"FF",
		188661 => x"FF",
		189685 => x"FF",
		190709 => x"FF",
		191733 => x"FF",
		192757 => x"FF",
		193781 => x"FF",
		194805 => x"FF",
		195829 => x"FF",
		196853 => x"FF",
		197877 => x"FF",
		198901 => x"FF",
		199925 => x"FF",
		200949 => x"FF",
		201973 => x"FF",
		202997 => x"FF",
		204021 => x"FF",
		205045 => x"FF",
		206069 => x"FF",
		207093 => x"FF",
		208117 => x"FF",
		209141 => x"FF",
		210165 => x"FF",
		211189 => x"FF",
		212213 => x"FF",
		213237 => x"FF",
		214261 => x"FF",
		215285 => x"FF",
		216309 => x"FF",
		217333 => x"FF",
		218357 => x"FF",
		219381 => x"FF",
		220405 => x"FF",
		221429 => x"FF",
		222453 => x"FF",
		223477 => x"FF",
		224501 => x"FF",
		225525 => x"FF",
		226549 => x"FF",
		227573 => x"FF",
		228597 => x"FF",
		229621 => x"FF",
		230645 => x"FF",
		231669 => x"FF",
		232693 => x"FF",
		233717 => x"FF",
		234741 => x"FF",
		235765 => x"FF",
		236789 => x"FF",
		237813 => x"FF",
		238837 => x"FF",
		239861 => x"FF",
		240885 => x"FF",
		241909 => x"FF",
		242933 => x"FF",
		243957 => x"FF",
		244981 => x"FF",
		246005 => x"FF",
		247029 => x"FF",
		248053 => x"FF",
		249077 => x"FF",
		250101 => x"FF",
		251125 => x"FF",
		252149 => x"FF",
		253173 => x"FF",
		254197 => x"FF",
		255221 => x"FF",
		256245 => x"FF",
		257269 => x"FF",
		258293 => x"FF",
		259317 => x"FF",
		260341 => x"FF",
		261365 => x"FF",
		262389 => x"FF",
		263413 => x"FF",
		264437 => x"FF",
		265461 => x"FF",
		266485 => x"FF",
		267509 => x"FF",
		268533 => x"FF",
		269557 => x"FF",
		270581 => x"FF",
		271605 => x"FF",
		272629 => x"FF",
		273653 => x"FF",
		274677 => x"FF",
		275701 => x"FF",
		276725 => x"FF",
		277749 => x"FF",
		278773 => x"FF",
		279797 => x"FF",
		280821 => x"FF",
		281845 => x"FF",
		282869 => x"FF",
		283893 => x"FF",
		284917 => x"FF",
		285941 => x"FF",
		286965 => x"FF",
		287989 => x"FF",
		289013 => x"FF",
		290037 => x"FF",
		291061 => x"FF",
		292085 => x"FF",
		293109 => x"FF",
		294133 => x"FF",
		295157 => x"FF",
		296181 => x"FF",
		297205 => x"FF",
		298229 => x"FF",
		299253 => x"FF",
		300277 => x"FF",
		301301 => x"FF",
		302325 => x"FF",
		303349 => x"FF",
		304373 => x"FF",
		305397 => x"FF",
		306421 => x"FF",
		307445 => x"FF",
		308469 => x"FF",
		309493 => x"FF",
		310517 => x"FF",
		311541 => x"FF",
		312565 => x"FF",
		313589 => x"FF",
		314613 => x"FF",
		315637 => x"FF",
		316661 => x"FF",
		317685 => x"FF",
		318709 => x"FF",
		319733 => x"FF",
		320757 => x"FF",
		321781 => x"FF",
		322805 => x"FF",
		323829 => x"FF",
		324853 => x"FF",
		325877 => x"FF",
		326901 => x"FF",
		327925 => x"FF",
		328949 => x"FF",
		329973 => x"FF",
		330997 => x"FF",
		332021 => x"FF",
		333045 => x"FF",
		334069 => x"FF",
		335093 => x"FF",
		336117 => x"FF",
		337141 => x"FF",
		338165 => x"FF",
		339189 => x"FF",
		340213 => x"FF",
		341237 => x"FF",
		342261 => x"FF",
		343285 => x"FF",
		344309 => x"FF",
		345333 => x"FF",
		346357 => x"FF",
		347381 => x"FF",
		348405 => x"FF",
		349429 => x"FF",
		350453 => x"FF",
		351477 => x"FF",
		352501 => x"FF",
		353525 => x"FF",
		354549 => x"FF",
		355573 => x"FF",
		356597 => x"FF",
		357621 => x"FF",
		358645 => x"FF",
		359669 => x"FF",
		360693 => x"FF",
		361717 => x"FF",
		362741 => x"FF",
		363765 => x"FF",
		364789 => x"FF",
		365813 => x"FF",
		366837 => x"FF",
		367861 => x"FF",
		368885 => x"FF",
		369909 => x"FF",
		370933 => x"FF",
		371957 => x"FF",
		372981 => x"FF",
		374005 => x"FF",
		375029 => x"FF",
		376053 => x"FF",
		377077 => x"FF",
		378101 => x"FF",
		379125 => x"FF",
		380149 => x"FF",
		381173 => x"FF",
		382197 => x"FF",
		383221 => x"FF",
		384245 => x"FF",
		385269 => x"FF",
		386293 => x"FF",
		387317 => x"FF",
		388341 => x"FF",
		389365 => x"FF",
		390389 => x"FF",
		391413 => x"FF",
		392437 => x"FF",
		393461 => x"FF",
		394485 => x"FF",
		395509 => x"FF",
		396533 => x"FF",
		397557 => x"FF",
		398581 => x"FF",
		399605 => x"FF",
		400629 => x"FF",
		401653 => x"FF",
		402677 => x"FF",
		403701 => x"FF",
		404725 => x"FF",
		405749 => x"FF",
		406773 => x"FF",
		407797 => x"FF",
		408821 => x"FF",
		409845 => x"FF",
		410869 => x"FF",
		411893 => x"FF",
		412917 => x"FF",
		413941 => x"FF",
		414965 => x"FF",
		415989 => x"FF",
		417013 => x"FF",
		418037 => x"FF",
		419061 => x"FF",
		420085 => x"FF",
		421109 => x"FF",
		422133 => x"FF",
		423157 => x"FF",
		424181 => x"FF",
		425205 => x"FF",
		426229 => x"FF",
		427253 => x"FF",
		428277 => x"FF",
		429301 => x"FF",
		430325 => x"FF",
		431349 => x"FF",
		432373 => x"FF",
		433397 => x"FF",
		434421 => x"FF",
		435445 => x"FF",
		436469 => x"FF",
		437493 => x"FF",
		438517 => x"FF",
		439541 => x"FF",
		440565 => x"FF",
		441589 => x"FF",
		442613 => x"FF",
		443637 => x"FF",
		444661 => x"FF",
		445685 => x"FF",
		446709 => x"FF",
		447733 => x"FF",
		448757 => x"FF",
		449781 => x"FF",
		450805 => x"FF",
		451829 => x"FF",
		452853 => x"FF",
		453877 => x"FF",
		454901 => x"FF",
		455925 => x"FF",
		456949 => x"FF",
		457973 => x"FF",
		458997 => x"FF",
		460021 => x"FF",
		461045 => x"FF",
		462069 => x"FF",
		463093 => x"FF",
		464117 => x"FF",
		465141 => x"FF",
		466165 => x"FF",
		467189 => x"FF",
		468213 => x"FF",
		469237 => x"FF",
		19702 => x"FF",
		20726 => x"FF",
		21750 => x"FF",
		22774 => x"FF",
		23798 => x"FF",
		24822 => x"FF",
		25846 => x"FF",
		26870 => x"FF",
		27894 => x"FF",
		28918 => x"FF",
		29942 => x"FF",
		30966 => x"FF",
		31990 => x"FF",
		33014 => x"FF",
		34038 => x"FF",
		35062 => x"FF",
		36086 => x"FF",
		37110 => x"FF",
		38134 => x"FF",
		39158 => x"FF",
		40182 => x"FF",
		41206 => x"FF",
		42230 => x"FF",
		43254 => x"FF",
		44278 => x"FF",
		45302 => x"FF",
		46326 => x"FF",
		47350 => x"FF",
		48374 => x"FF",
		49398 => x"FF",
		50422 => x"FF",
		51446 => x"FF",
		52470 => x"FF",
		53494 => x"FF",
		54518 => x"FF",
		55542 => x"FF",
		56566 => x"FF",
		57590 => x"FF",
		58614 => x"FF",
		59638 => x"FF",
		60662 => x"FF",
		61686 => x"FF",
		62710 => x"FF",
		63734 => x"FF",
		64758 => x"FF",
		65782 => x"FF",
		66806 => x"FF",
		67830 => x"FF",
		68854 => x"FF",
		69878 => x"FF",
		70902 => x"FF",
		71926 => x"FF",
		72950 => x"FF",
		73974 => x"FF",
		74998 => x"FF",
		76022 => x"FF",
		77046 => x"FF",
		78070 => x"FF",
		79094 => x"FF",
		80118 => x"FF",
		81142 => x"FF",
		82166 => x"FF",
		83190 => x"FF",
		84214 => x"FF",
		85238 => x"FF",
		86262 => x"FF",
		87286 => x"FF",
		88310 => x"FF",
		89334 => x"FF",
		90358 => x"FF",
		91382 => x"FF",
		92406 => x"FF",
		93430 => x"FF",
		94454 => x"FF",
		95478 => x"FF",
		96502 => x"FF",
		97526 => x"FF",
		98550 => x"FF",
		99574 => x"FF",
		100598 => x"FF",
		101622 => x"FF",
		102646 => x"FF",
		103670 => x"FF",
		104694 => x"FF",
		105718 => x"FF",
		106742 => x"FF",
		107766 => x"FF",
		108790 => x"FF",
		109814 => x"FF",
		110838 => x"FF",
		111862 => x"FF",
		112886 => x"FF",
		113910 => x"FF",
		114934 => x"FF",
		115958 => x"FF",
		116982 => x"FF",
		118006 => x"FF",
		119030 => x"FF",
		120054 => x"FF",
		121078 => x"FF",
		122102 => x"FF",
		123126 => x"FF",
		124150 => x"FF",
		125174 => x"FF",
		126198 => x"FF",
		127222 => x"FF",
		128246 => x"FF",
		129270 => x"FF",
		130294 => x"FF",
		131318 => x"FF",
		132342 => x"FF",
		133366 => x"FF",
		134390 => x"FF",
		135414 => x"FF",
		136438 => x"FF",
		137462 => x"FF",
		138486 => x"FF",
		139510 => x"FF",
		140534 => x"FF",
		141558 => x"FF",
		142582 => x"FF",
		143606 => x"FF",
		144630 => x"FF",
		145654 => x"FF",
		146678 => x"FF",
		147702 => x"FF",
		148726 => x"FF",
		149750 => x"FF",
		150774 => x"FF",
		151798 => x"FF",
		152822 => x"FF",
		153846 => x"FF",
		154870 => x"FF",
		155894 => x"FF",
		156918 => x"FF",
		157942 => x"FF",
		158966 => x"FF",
		159990 => x"FF",
		161014 => x"FF",
		162038 => x"FF",
		163062 => x"FF",
		164086 => x"FF",
		165110 => x"FF",
		166134 => x"FF",
		167158 => x"FF",
		168182 => x"FF",
		169206 => x"FF",
		170230 => x"FF",
		171254 => x"FF",
		172278 => x"FF",
		173302 => x"FF",
		174326 => x"FF",
		175350 => x"FF",
		176374 => x"FF",
		177398 => x"FF",
		178422 => x"FF",
		179446 => x"FF",
		180470 => x"FF",
		181494 => x"FF",
		182518 => x"FF",
		183542 => x"FF",
		184566 => x"FF",
		185590 => x"FF",
		186614 => x"FF",
		187638 => x"FF",
		188662 => x"FF",
		189686 => x"FF",
		190710 => x"FF",
		191734 => x"FF",
		192758 => x"FF",
		193782 => x"FF",
		194806 => x"FF",
		195830 => x"FF",
		196854 => x"FF",
		197878 => x"FF",
		198902 => x"FF",
		199926 => x"FF",
		200950 => x"FF",
		201974 => x"FF",
		202998 => x"FF",
		204022 => x"FF",
		205046 => x"FF",
		206070 => x"FF",
		207094 => x"FF",
		208118 => x"FF",
		209142 => x"FF",
		210166 => x"FF",
		211190 => x"FF",
		212214 => x"FF",
		213238 => x"FF",
		214262 => x"FF",
		215286 => x"FF",
		216310 => x"FF",
		217334 => x"FF",
		218358 => x"FF",
		219382 => x"FF",
		220406 => x"FF",
		221430 => x"FF",
		222454 => x"FF",
		223478 => x"FF",
		224502 => x"FF",
		225526 => x"FF",
		226550 => x"FF",
		227574 => x"FF",
		228598 => x"FF",
		229622 => x"FF",
		230646 => x"FF",
		231670 => x"FF",
		232694 => x"FF",
		233718 => x"FF",
		234742 => x"FF",
		235766 => x"FF",
		236790 => x"FF",
		237814 => x"FF",
		238838 => x"FF",
		239862 => x"FF",
		240886 => x"FF",
		241910 => x"FF",
		242934 => x"FF",
		243958 => x"FF",
		244982 => x"FF",
		246006 => x"FF",
		247030 => x"FF",
		248054 => x"FF",
		249078 => x"FF",
		250102 => x"FF",
		251126 => x"FF",
		252150 => x"FF",
		253174 => x"FF",
		254198 => x"FF",
		255222 => x"FF",
		256246 => x"FF",
		257270 => x"FF",
		258294 => x"FF",
		259318 => x"FF",
		260342 => x"FF",
		261366 => x"FF",
		262390 => x"FF",
		263414 => x"FF",
		264438 => x"FF",
		265462 => x"FF",
		266486 => x"FF",
		267510 => x"FF",
		268534 => x"FF",
		269558 => x"FF",
		270582 => x"FF",
		271606 => x"FF",
		272630 => x"FF",
		273654 => x"FF",
		274678 => x"FF",
		275702 => x"FF",
		276726 => x"FF",
		277750 => x"FF",
		278774 => x"FF",
		279798 => x"FF",
		280822 => x"FF",
		281846 => x"FF",
		282870 => x"FF",
		283894 => x"FF",
		284918 => x"FF",
		285942 => x"FF",
		286966 => x"FF",
		287990 => x"FF",
		289014 => x"FF",
		290038 => x"FF",
		291062 => x"FF",
		292086 => x"FF",
		293110 => x"FF",
		294134 => x"FF",
		295158 => x"FF",
		296182 => x"FF",
		297206 => x"FF",
		298230 => x"FF",
		299254 => x"FF",
		300278 => x"FF",
		301302 => x"FF",
		302326 => x"FF",
		303350 => x"FF",
		304374 => x"FF",
		305398 => x"FF",
		306422 => x"FF",
		307446 => x"FF",
		308470 => x"FF",
		309494 => x"FF",
		310518 => x"FF",
		311542 => x"FF",
		312566 => x"FF",
		313590 => x"FF",
		314614 => x"FF",
		315638 => x"FF",
		316662 => x"FF",
		317686 => x"FF",
		318710 => x"FF",
		319734 => x"FF",
		320758 => x"FF",
		321782 => x"FF",
		322806 => x"FF",
		323830 => x"FF",
		324854 => x"FF",
		325878 => x"FF",
		326902 => x"FF",
		327926 => x"FF",
		328950 => x"FF",
		329974 => x"FF",
		330998 => x"FF",
		332022 => x"FF",
		333046 => x"FF",
		334070 => x"FF",
		335094 => x"FF",
		336118 => x"FF",
		337142 => x"FF",
		338166 => x"FF",
		339190 => x"FF",
		340214 => x"FF",
		341238 => x"FF",
		342262 => x"FF",
		343286 => x"FF",
		344310 => x"FF",
		345334 => x"FF",
		346358 => x"FF",
		347382 => x"FF",
		348406 => x"FF",
		349430 => x"FF",
		350454 => x"FF",
		351478 => x"FF",
		352502 => x"FF",
		353526 => x"FF",
		354550 => x"FF",
		355574 => x"FF",
		356598 => x"FF",
		357622 => x"FF",
		358646 => x"FF",
		359670 => x"FF",
		360694 => x"FF",
		361718 => x"FF",
		362742 => x"FF",
		363766 => x"FF",
		364790 => x"FF",
		365814 => x"FF",
		366838 => x"FF",
		367862 => x"FF",
		368886 => x"FF",
		369910 => x"FF",
		370934 => x"FF",
		371958 => x"FF",
		372982 => x"FF",
		374006 => x"FF",
		375030 => x"FF",
		376054 => x"FF",
		377078 => x"FF",
		378102 => x"FF",
		379126 => x"FF",
		380150 => x"FF",
		381174 => x"FF",
		382198 => x"FF",
		383222 => x"FF",
		384246 => x"FF",
		385270 => x"FF",
		386294 => x"FF",
		387318 => x"FF",
		388342 => x"FF",
		389366 => x"FF",
		390390 => x"FF",
		391414 => x"FF",
		392438 => x"FF",
		393462 => x"FF",
		394486 => x"FF",
		395510 => x"FF",
		396534 => x"FF",
		397558 => x"FF",
		398582 => x"FF",
		399606 => x"FF",
		400630 => x"FF",
		401654 => x"FF",
		402678 => x"FF",
		403702 => x"FF",
		404726 => x"FF",
		405750 => x"FF",
		406774 => x"FF",
		407798 => x"FF",
		408822 => x"FF",
		409846 => x"FF",
		410870 => x"FF",
		411894 => x"FF",
		412918 => x"FF",
		413942 => x"FF",
		414966 => x"FF",
		415990 => x"FF",
		417014 => x"FF",
		418038 => x"FF",
		419062 => x"FF",
		420086 => x"FF",
		421110 => x"FF",
		422134 => x"FF",
		423158 => x"FF",
		424182 => x"FF",
		425206 => x"FF",
		426230 => x"FF",
		427254 => x"FF",
		428278 => x"FF",
		429302 => x"FF",
		430326 => x"FF",
		431350 => x"FF",
		432374 => x"FF",
		433398 => x"FF",
		434422 => x"FF",
		435446 => x"FF",
		436470 => x"FF",
		437494 => x"FF",
		438518 => x"FF",
		439542 => x"FF",
		440566 => x"FF",
		441590 => x"FF",
		442614 => x"FF",
		443638 => x"FF",
		444662 => x"FF",
		445686 => x"FF",
		446710 => x"FF",
		447734 => x"FF",
		448758 => x"FF",
		449782 => x"FF",
		450806 => x"FF",
		451830 => x"FF",
		452854 => x"FF",
		453878 => x"FF",
		454902 => x"FF",
		455926 => x"FF",
		456950 => x"FF",
		457974 => x"FF",
		458998 => x"FF",
		460022 => x"FF",
		461046 => x"FF",
		462070 => x"FF",
		463094 => x"FF",
		464118 => x"FF",
		465142 => x"FF",
		466166 => x"FF",
		467190 => x"FF",
		468214 => x"FF",
		469238 => x"FF",
		19703 => x"FF",
		20727 => x"FF",
		21751 => x"FF",
		22775 => x"FF",
		23799 => x"FF",
		24823 => x"FF",
		25847 => x"FF",
		26871 => x"FF",
		27895 => x"FF",
		28919 => x"FF",
		29943 => x"FF",
		30967 => x"FF",
		31991 => x"FF",
		33015 => x"FF",
		34039 => x"FF",
		35063 => x"FF",
		36087 => x"FF",
		37111 => x"FF",
		38135 => x"FF",
		39159 => x"FF",
		40183 => x"FF",
		41207 => x"FF",
		42231 => x"FF",
		43255 => x"FF",
		44279 => x"FF",
		45303 => x"FF",
		46327 => x"FF",
		47351 => x"FF",
		48375 => x"FF",
		49399 => x"FF",
		50423 => x"FF",
		51447 => x"FF",
		52471 => x"FF",
		53495 => x"FF",
		54519 => x"FF",
		55543 => x"FF",
		56567 => x"FF",
		57591 => x"FF",
		58615 => x"FF",
		59639 => x"FF",
		60663 => x"FF",
		61687 => x"FF",
		62711 => x"FF",
		63735 => x"FF",
		64759 => x"FF",
		65783 => x"FF",
		66807 => x"FF",
		67831 => x"FF",
		68855 => x"FF",
		69879 => x"FF",
		70903 => x"FF",
		71927 => x"FF",
		72951 => x"FF",
		73975 => x"FF",
		74999 => x"FF",
		76023 => x"FF",
		77047 => x"FF",
		78071 => x"FF",
		79095 => x"FF",
		80119 => x"FF",
		81143 => x"FF",
		82167 => x"FF",
		83191 => x"FF",
		84215 => x"FF",
		85239 => x"FF",
		86263 => x"FF",
		87287 => x"FF",
		88311 => x"FF",
		89335 => x"FF",
		90359 => x"FF",
		91383 => x"FF",
		92407 => x"FF",
		93431 => x"FF",
		94455 => x"FF",
		95479 => x"FF",
		96503 => x"FF",
		97527 => x"FF",
		98551 => x"FF",
		99575 => x"FF",
		100599 => x"FF",
		101623 => x"FF",
		102647 => x"FF",
		103671 => x"FF",
		104695 => x"FF",
		105719 => x"FF",
		106743 => x"FF",
		107767 => x"FF",
		108791 => x"FF",
		109815 => x"FF",
		110839 => x"FF",
		111863 => x"FF",
		112887 => x"FF",
		113911 => x"FF",
		114935 => x"FF",
		115959 => x"FF",
		116983 => x"FF",
		118007 => x"FF",
		119031 => x"FF",
		120055 => x"FF",
		121079 => x"FF",
		122103 => x"FF",
		123127 => x"FF",
		124151 => x"FF",
		125175 => x"FF",
		126199 => x"FF",
		127223 => x"FF",
		128247 => x"FF",
		129271 => x"FF",
		130295 => x"FF",
		131319 => x"FF",
		132343 => x"FF",
		133367 => x"FF",
		134391 => x"FF",
		135415 => x"FF",
		136439 => x"FF",
		137463 => x"FF",
		138487 => x"FF",
		139511 => x"FF",
		140535 => x"FF",
		141559 => x"FF",
		142583 => x"FF",
		143607 => x"FF",
		144631 => x"FF",
		145655 => x"FF",
		146679 => x"FF",
		147703 => x"FF",
		148727 => x"FF",
		149751 => x"FF",
		150775 => x"FF",
		151799 => x"FF",
		152823 => x"FF",
		153847 => x"FF",
		154871 => x"FF",
		155895 => x"FF",
		156919 => x"FF",
		157943 => x"FF",
		158967 => x"FF",
		159991 => x"FF",
		161015 => x"FF",
		162039 => x"FF",
		163063 => x"FF",
		164087 => x"FF",
		165111 => x"FF",
		166135 => x"FF",
		167159 => x"FF",
		168183 => x"FF",
		169207 => x"FF",
		170231 => x"FF",
		171255 => x"FF",
		172279 => x"FF",
		173303 => x"FF",
		174327 => x"FF",
		175351 => x"FF",
		176375 => x"FF",
		177399 => x"FF",
		178423 => x"FF",
		179447 => x"FF",
		180471 => x"FF",
		181495 => x"FF",
		182519 => x"FF",
		183543 => x"FF",
		184567 => x"FF",
		185591 => x"FF",
		186615 => x"FF",
		187639 => x"FF",
		188663 => x"FF",
		189687 => x"FF",
		190711 => x"FF",
		191735 => x"FF",
		192759 => x"FF",
		193783 => x"FF",
		194807 => x"FF",
		195831 => x"FF",
		196855 => x"FF",
		197879 => x"FF",
		198903 => x"FF",
		199927 => x"FF",
		200951 => x"FF",
		201975 => x"FF",
		202999 => x"FF",
		204023 => x"FF",
		205047 => x"FF",
		206071 => x"FF",
		207095 => x"FF",
		208119 => x"FF",
		209143 => x"FF",
		210167 => x"FF",
		211191 => x"FF",
		212215 => x"FF",
		213239 => x"FF",
		214263 => x"FF",
		215287 => x"FF",
		216311 => x"FF",
		217335 => x"FF",
		218359 => x"FF",
		219383 => x"FF",
		220407 => x"FF",
		221431 => x"FF",
		222455 => x"FF",
		223479 => x"FF",
		224503 => x"FF",
		225527 => x"FF",
		226551 => x"FF",
		227575 => x"FF",
		228599 => x"FF",
		229623 => x"FF",
		230647 => x"FF",
		231671 => x"FF",
		232695 => x"FF",
		233719 => x"FF",
		234743 => x"FF",
		235767 => x"FF",
		236791 => x"FF",
		237815 => x"FF",
		238839 => x"FF",
		239863 => x"FF",
		240887 => x"FF",
		241911 => x"FF",
		242935 => x"FF",
		243959 => x"FF",
		244983 => x"FF",
		246007 => x"FF",
		247031 => x"FF",
		248055 => x"FF",
		249079 => x"FF",
		250103 => x"FF",
		251127 => x"FF",
		252151 => x"FF",
		253175 => x"FF",
		254199 => x"FF",
		255223 => x"FF",
		256247 => x"FF",
		257271 => x"FF",
		258295 => x"FF",
		259319 => x"FF",
		260343 => x"FF",
		261367 => x"FF",
		262391 => x"FF",
		263415 => x"FF",
		264439 => x"FF",
		265463 => x"FF",
		266487 => x"FF",
		267511 => x"FF",
		268535 => x"FF",
		269559 => x"FF",
		270583 => x"FF",
		271607 => x"FF",
		272631 => x"FF",
		273655 => x"FF",
		274679 => x"FF",
		275703 => x"FF",
		276727 => x"FF",
		277751 => x"FF",
		278775 => x"FF",
		279799 => x"FF",
		280823 => x"FF",
		281847 => x"FF",
		282871 => x"FF",
		283895 => x"FF",
		284919 => x"FF",
		285943 => x"FF",
		286967 => x"FF",
		287991 => x"FF",
		289015 => x"FF",
		290039 => x"FF",
		291063 => x"FF",
		292087 => x"FF",
		293111 => x"FF",
		294135 => x"FF",
		295159 => x"FF",
		296183 => x"FF",
		297207 => x"FF",
		298231 => x"FF",
		299255 => x"FF",
		300279 => x"FF",
		301303 => x"FF",
		302327 => x"FF",
		303351 => x"FF",
		304375 => x"FF",
		305399 => x"FF",
		306423 => x"FF",
		307447 => x"FF",
		308471 => x"FF",
		309495 => x"FF",
		310519 => x"FF",
		311543 => x"FF",
		312567 => x"FF",
		313591 => x"FF",
		314615 => x"FF",
		315639 => x"FF",
		316663 => x"FF",
		317687 => x"FF",
		318711 => x"FF",
		319735 => x"FF",
		320759 => x"FF",
		321783 => x"FF",
		322807 => x"FF",
		323831 => x"FF",
		324855 => x"FF",
		325879 => x"FF",
		326903 => x"FF",
		327927 => x"FF",
		328951 => x"FF",
		329975 => x"FF",
		330999 => x"FF",
		332023 => x"FF",
		333047 => x"FF",
		334071 => x"FF",
		335095 => x"FF",
		336119 => x"FF",
		337143 => x"FF",
		338167 => x"FF",
		339191 => x"FF",
		340215 => x"FF",
		341239 => x"FF",
		342263 => x"FF",
		343287 => x"FF",
		344311 => x"FF",
		345335 => x"FF",
		346359 => x"FF",
		347383 => x"FF",
		348407 => x"FF",
		349431 => x"FF",
		350455 => x"FF",
		351479 => x"FF",
		352503 => x"FF",
		353527 => x"FF",
		354551 => x"FF",
		355575 => x"FF",
		356599 => x"FF",
		357623 => x"FF",
		358647 => x"FF",
		359671 => x"FF",
		360695 => x"FF",
		361719 => x"FF",
		362743 => x"FF",
		363767 => x"FF",
		364791 => x"FF",
		365815 => x"FF",
		366839 => x"FF",
		367863 => x"FF",
		368887 => x"FF",
		369911 => x"FF",
		370935 => x"FF",
		371959 => x"FF",
		372983 => x"FF",
		374007 => x"FF",
		375031 => x"FF",
		376055 => x"FF",
		377079 => x"FF",
		378103 => x"FF",
		379127 => x"FF",
		380151 => x"FF",
		381175 => x"FF",
		382199 => x"FF",
		383223 => x"FF",
		384247 => x"FF",
		385271 => x"FF",
		386295 => x"FF",
		387319 => x"FF",
		388343 => x"FF",
		389367 => x"FF",
		390391 => x"FF",
		391415 => x"FF",
		392439 => x"FF",
		393463 => x"FF",
		394487 => x"FF",
		395511 => x"FF",
		396535 => x"FF",
		397559 => x"FF",
		398583 => x"FF",
		399607 => x"FF",
		400631 => x"FF",
		401655 => x"FF",
		402679 => x"FF",
		403703 => x"FF",
		404727 => x"FF",
		405751 => x"FF",
		406775 => x"FF",
		407799 => x"FF",
		408823 => x"FF",
		409847 => x"FF",
		410871 => x"FF",
		411895 => x"FF",
		412919 => x"FF",
		413943 => x"FF",
		414967 => x"FF",
		415991 => x"FF",
		417015 => x"FF",
		418039 => x"FF",
		419063 => x"FF",
		420087 => x"FF",
		421111 => x"FF",
		422135 => x"FF",
		423159 => x"FF",
		424183 => x"FF",
		425207 => x"FF",
		426231 => x"FF",
		427255 => x"FF",
		428279 => x"FF",
		429303 => x"FF",
		430327 => x"FF",
		431351 => x"FF",
		432375 => x"FF",
		433399 => x"FF",
		434423 => x"FF",
		435447 => x"FF",
		436471 => x"FF",
		437495 => x"FF",
		438519 => x"FF",
		439543 => x"FF",
		440567 => x"FF",
		441591 => x"FF",
		442615 => x"FF",
		443639 => x"FF",
		444663 => x"FF",
		445687 => x"FF",
		446711 => x"FF",
		447735 => x"FF",
		448759 => x"FF",
		449783 => x"FF",
		450807 => x"FF",
		451831 => x"FF",
		452855 => x"FF",
		453879 => x"FF",
		454903 => x"FF",
		455927 => x"FF",
		456951 => x"FF",
		457975 => x"FF",
		458999 => x"FF",
		460023 => x"FF",
		461047 => x"FF",
		462071 => x"FF",
		463095 => x"FF",
		464119 => x"FF",
		465143 => x"FF",
		466167 => x"FF",
		467191 => x"FF",
		468215 => x"FF",
		469239 => x"FF",
		19704 => x"FF",
		20728 => x"FF",
		21752 => x"FF",
		22776 => x"FF",
		23800 => x"FF",
		24824 => x"FF",
		25848 => x"FF",
		26872 => x"FF",
		27896 => x"FF",
		28920 => x"FF",
		29944 => x"FF",
		30968 => x"FF",
		31992 => x"FF",
		33016 => x"FF",
		34040 => x"FF",
		35064 => x"FF",
		36088 => x"FF",
		37112 => x"FF",
		38136 => x"FF",
		39160 => x"FF",
		40184 => x"FF",
		41208 => x"FF",
		42232 => x"FF",
		43256 => x"FF",
		44280 => x"FF",
		45304 => x"FF",
		46328 => x"FF",
		47352 => x"FF",
		48376 => x"FF",
		49400 => x"FF",
		50424 => x"FF",
		51448 => x"FF",
		52472 => x"FF",
		53496 => x"FF",
		54520 => x"FF",
		55544 => x"FF",
		56568 => x"FF",
		57592 => x"FF",
		58616 => x"FF",
		59640 => x"FF",
		60664 => x"FF",
		61688 => x"FF",
		62712 => x"FF",
		63736 => x"FF",
		64760 => x"FF",
		65784 => x"FF",
		66808 => x"FF",
		67832 => x"FF",
		68856 => x"FF",
		69880 => x"FF",
		70904 => x"FF",
		71928 => x"FF",
		72952 => x"FF",
		73976 => x"FF",
		75000 => x"FF",
		76024 => x"FF",
		77048 => x"FF",
		78072 => x"FF",
		79096 => x"FF",
		80120 => x"FF",
		81144 => x"FF",
		82168 => x"FF",
		83192 => x"FF",
		84216 => x"FF",
		85240 => x"FF",
		86264 => x"FF",
		87288 => x"FF",
		88312 => x"FF",
		89336 => x"FF",
		90360 => x"FF",
		91384 => x"FF",
		92408 => x"FF",
		93432 => x"FF",
		94456 => x"FF",
		95480 => x"FF",
		96504 => x"FF",
		97528 => x"FF",
		98552 => x"FF",
		99576 => x"FF",
		100600 => x"FF",
		101624 => x"FF",
		102648 => x"FF",
		103672 => x"FF",
		104696 => x"FF",
		105720 => x"FF",
		106744 => x"FF",
		107768 => x"FF",
		108792 => x"FF",
		109816 => x"FF",
		110840 => x"FF",
		111864 => x"FF",
		112888 => x"FF",
		113912 => x"FF",
		114936 => x"FF",
		115960 => x"FF",
		116984 => x"FF",
		118008 => x"FF",
		119032 => x"FF",
		120056 => x"FF",
		121080 => x"FF",
		122104 => x"FF",
		123128 => x"FF",
		124152 => x"FF",
		125176 => x"FF",
		126200 => x"FF",
		127224 => x"FF",
		128248 => x"FF",
		129272 => x"FF",
		130296 => x"FF",
		131320 => x"FF",
		132344 => x"FF",
		133368 => x"FF",
		134392 => x"FF",
		135416 => x"FF",
		136440 => x"FF",
		137464 => x"FF",
		138488 => x"FF",
		139512 => x"FF",
		140536 => x"FF",
		141560 => x"FF",
		142584 => x"FF",
		143608 => x"FF",
		144632 => x"FF",
		145656 => x"FF",
		146680 => x"FF",
		147704 => x"FF",
		148728 => x"FF",
		149752 => x"FF",
		150776 => x"FF",
		151800 => x"FF",
		152824 => x"FF",
		153848 => x"FF",
		154872 => x"FF",
		155896 => x"FF",
		156920 => x"FF",
		157944 => x"FF",
		158968 => x"FF",
		159992 => x"FF",
		161016 => x"FF",
		162040 => x"FF",
		163064 => x"FF",
		164088 => x"FF",
		165112 => x"FF",
		166136 => x"FF",
		167160 => x"FF",
		168184 => x"FF",
		169208 => x"FF",
		170232 => x"FF",
		171256 => x"FF",
		172280 => x"FF",
		173304 => x"FF",
		174328 => x"FF",
		175352 => x"FF",
		176376 => x"FF",
		177400 => x"FF",
		178424 => x"FF",
		179448 => x"FF",
		180472 => x"FF",
		181496 => x"FF",
		182520 => x"FF",
		183544 => x"FF",
		184568 => x"FF",
		185592 => x"FF",
		186616 => x"FF",
		187640 => x"FF",
		188664 => x"FF",
		189688 => x"FF",
		190712 => x"FF",
		191736 => x"FF",
		192760 => x"FF",
		193784 => x"FF",
		194808 => x"FF",
		195832 => x"FF",
		196856 => x"FF",
		197880 => x"FF",
		198904 => x"FF",
		199928 => x"FF",
		200952 => x"FF",
		201976 => x"FF",
		203000 => x"FF",
		204024 => x"FF",
		205048 => x"FF",
		206072 => x"FF",
		207096 => x"FF",
		208120 => x"FF",
		209144 => x"FF",
		210168 => x"FF",
		211192 => x"FF",
		212216 => x"FF",
		213240 => x"FF",
		214264 => x"FF",
		215288 => x"FF",
		216312 => x"FF",
		217336 => x"FF",
		218360 => x"FF",
		219384 => x"FF",
		220408 => x"FF",
		221432 => x"FF",
		222456 => x"FF",
		223480 => x"FF",
		224504 => x"FF",
		225528 => x"FF",
		226552 => x"FF",
		227576 => x"FF",
		228600 => x"FF",
		229624 => x"FF",
		230648 => x"FF",
		231672 => x"FF",
		232696 => x"FF",
		233720 => x"FF",
		234744 => x"FF",
		235768 => x"FF",
		236792 => x"FF",
		237816 => x"FF",
		238840 => x"FF",
		239864 => x"FF",
		240888 => x"FF",
		241912 => x"FF",
		242936 => x"FF",
		243960 => x"FF",
		244984 => x"FF",
		246008 => x"FF",
		247032 => x"FF",
		248056 => x"FF",
		249080 => x"FF",
		250104 => x"FF",
		251128 => x"FF",
		252152 => x"FF",
		253176 => x"FF",
		254200 => x"FF",
		255224 => x"FF",
		256248 => x"FF",
		257272 => x"FF",
		258296 => x"FF",
		259320 => x"FF",
		260344 => x"FF",
		261368 => x"FF",
		262392 => x"FF",
		263416 => x"FF",
		264440 => x"FF",
		265464 => x"FF",
		266488 => x"FF",
		267512 => x"FF",
		268536 => x"FF",
		269560 => x"FF",
		270584 => x"FF",
		271608 => x"FF",
		272632 => x"FF",
		273656 => x"FF",
		274680 => x"FF",
		275704 => x"FF",
		276728 => x"FF",
		277752 => x"FF",
		278776 => x"FF",
		279800 => x"FF",
		280824 => x"FF",
		281848 => x"FF",
		282872 => x"FF",
		283896 => x"FF",
		284920 => x"FF",
		285944 => x"FF",
		286968 => x"FF",
		287992 => x"FF",
		289016 => x"FF",
		290040 => x"FF",
		291064 => x"FF",
		292088 => x"FF",
		293112 => x"FF",
		294136 => x"FF",
		295160 => x"FF",
		296184 => x"FF",
		297208 => x"FF",
		298232 => x"FF",
		299256 => x"FF",
		300280 => x"FF",
		301304 => x"FF",
		302328 => x"FF",
		303352 => x"FF",
		304376 => x"FF",
		305400 => x"FF",
		306424 => x"FF",
		307448 => x"FF",
		308472 => x"FF",
		309496 => x"FF",
		310520 => x"FF",
		311544 => x"FF",
		312568 => x"FF",
		313592 => x"FF",
		314616 => x"FF",
		315640 => x"FF",
		316664 => x"FF",
		317688 => x"FF",
		318712 => x"FF",
		319736 => x"FF",
		320760 => x"FF",
		321784 => x"FF",
		322808 => x"FF",
		323832 => x"FF",
		324856 => x"FF",
		325880 => x"FF",
		326904 => x"FF",
		327928 => x"FF",
		328952 => x"FF",
		329976 => x"FF",
		331000 => x"FF",
		332024 => x"FF",
		333048 => x"FF",
		334072 => x"FF",
		335096 => x"FF",
		336120 => x"FF",
		337144 => x"FF",
		338168 => x"FF",
		339192 => x"FF",
		340216 => x"FF",
		341240 => x"FF",
		342264 => x"FF",
		343288 => x"FF",
		344312 => x"FF",
		345336 => x"FF",
		346360 => x"FF",
		347384 => x"FF",
		348408 => x"FF",
		349432 => x"FF",
		350456 => x"FF",
		351480 => x"FF",
		352504 => x"FF",
		353528 => x"FF",
		354552 => x"FF",
		355576 => x"FF",
		356600 => x"FF",
		357624 => x"FF",
		358648 => x"FF",
		359672 => x"FF",
		360696 => x"FF",
		361720 => x"FF",
		362744 => x"FF",
		363768 => x"FF",
		364792 => x"FF",
		365816 => x"FF",
		366840 => x"FF",
		367864 => x"FF",
		368888 => x"FF",
		369912 => x"FF",
		370936 => x"FF",
		371960 => x"FF",
		372984 => x"FF",
		374008 => x"FF",
		375032 => x"FF",
		376056 => x"FF",
		377080 => x"FF",
		378104 => x"FF",
		379128 => x"FF",
		380152 => x"FF",
		381176 => x"FF",
		382200 => x"FF",
		383224 => x"FF",
		384248 => x"FF",
		385272 => x"FF",
		386296 => x"FF",
		387320 => x"FF",
		388344 => x"FF",
		389368 => x"FF",
		390392 => x"FF",
		391416 => x"FF",
		392440 => x"FF",
		393464 => x"FF",
		394488 => x"FF",
		395512 => x"FF",
		396536 => x"FF",
		397560 => x"FF",
		398584 => x"FF",
		399608 => x"FF",
		400632 => x"FF",
		401656 => x"FF",
		402680 => x"FF",
		403704 => x"FF",
		404728 => x"FF",
		405752 => x"FF",
		406776 => x"FF",
		407800 => x"FF",
		408824 => x"FF",
		409848 => x"FF",
		410872 => x"FF",
		411896 => x"FF",
		412920 => x"FF",
		413944 => x"FF",
		414968 => x"FF",
		415992 => x"FF",
		417016 => x"FF",
		418040 => x"FF",
		419064 => x"FF",
		420088 => x"FF",
		421112 => x"FF",
		422136 => x"FF",
		423160 => x"FF",
		424184 => x"FF",
		425208 => x"FF",
		426232 => x"FF",
		427256 => x"FF",
		428280 => x"FF",
		429304 => x"FF",
		430328 => x"FF",
		431352 => x"FF",
		432376 => x"FF",
		433400 => x"FF",
		434424 => x"FF",
		435448 => x"FF",
		436472 => x"FF",
		437496 => x"FF",
		438520 => x"FF",
		439544 => x"FF",
		440568 => x"FF",
		441592 => x"FF",
		442616 => x"FF",
		443640 => x"FF",
		444664 => x"FF",
		445688 => x"FF",
		446712 => x"FF",
		447736 => x"FF",
		448760 => x"FF",
		449784 => x"FF",
		450808 => x"FF",
		451832 => x"FF",
		452856 => x"FF",
		453880 => x"FF",
		454904 => x"FF",
		455928 => x"FF",
		456952 => x"FF",
		457976 => x"FF",
		459000 => x"FF",
		460024 => x"FF",
		461048 => x"FF",
		462072 => x"FF",
		463096 => x"FF",
		464120 => x"FF",
		465144 => x"FF",
		466168 => x"FF",
		467192 => x"FF",
		468216 => x"FF",
		469240 => x"FF",
		19705 => x"FF",
		20729 => x"FF",
		21753 => x"FF",
		22777 => x"FF",
		23801 => x"FF",
		168185 => x"FF",
		169209 => x"FF",
		170233 => x"FF",
		171257 => x"FF",
		172281 => x"FF",
		316665 => x"FF",
		317689 => x"FF",
		318713 => x"FF",
		319737 => x"FF",
		320761 => x"FF",
		465145 => x"FF",
		466169 => x"FF",
		467193 => x"FF",
		468217 => x"FF",
		469241 => x"FF",
		19706 => x"FF",
		20730 => x"FF",
		21754 => x"FF",
		22778 => x"FF",
		23802 => x"FF",
		168186 => x"FF",
		169210 => x"FF",
		170234 => x"FF",
		171258 => x"FF",
		172282 => x"FF",
		316666 => x"FF",
		317690 => x"FF",
		318714 => x"FF",
		319738 => x"FF",
		320762 => x"FF",
		465146 => x"FF",
		466170 => x"FF",
		467194 => x"FF",
		468218 => x"FF",
		469242 => x"FF",
		19707 => x"FF",
		20731 => x"FF",
		21755 => x"FF",
		22779 => x"FF",
		23803 => x"FF",
		168187 => x"FF",
		169211 => x"FF",
		170235 => x"FF",
		171259 => x"FF",
		172283 => x"FF",
		316667 => x"FF",
		317691 => x"FF",
		318715 => x"FF",
		319739 => x"FF",
		320763 => x"FF",
		465147 => x"FF",
		466171 => x"FF",
		467195 => x"FF",
		468219 => x"FF",
		469243 => x"FF",
		19708 => x"FF",
		20732 => x"FF",
		21756 => x"FF",
		22780 => x"FF",
		23804 => x"FF",
		168188 => x"FF",
		169212 => x"FF",
		170236 => x"FF",
		171260 => x"FF",
		172284 => x"FF",
		316668 => x"FF",
		317692 => x"FF",
		318716 => x"FF",
		319740 => x"FF",
		320764 => x"FF",
		465148 => x"FF",
		466172 => x"FF",
		467196 => x"FF",
		468220 => x"FF",
		469244 => x"FF",
		19709 => x"FF",
		20733 => x"FF",
		21757 => x"FF",
		22781 => x"FF",
		23805 => x"FF",
		168189 => x"FF",
		169213 => x"FF",
		170237 => x"FF",
		171261 => x"FF",
		172285 => x"FF",
		316669 => x"FF",
		317693 => x"FF",
		318717 => x"FF",
		319741 => x"FF",
		320765 => x"FF",
		465149 => x"FF",
		466173 => x"FF",
		467197 => x"FF",
		468221 => x"FF",
		469245 => x"FF",
		19710 => x"FF",
		20734 => x"FF",
		21758 => x"FF",
		22782 => x"FF",
		23806 => x"FF",
		168190 => x"FF",
		169214 => x"FF",
		170238 => x"FF",
		171262 => x"FF",
		172286 => x"FF",
		316670 => x"FF",
		317694 => x"FF",
		318718 => x"FF",
		319742 => x"FF",
		320766 => x"FF",
		465150 => x"FF",
		466174 => x"FF",
		467198 => x"FF",
		468222 => x"FF",
		469246 => x"FF",
		19711 => x"FF",
		20735 => x"FF",
		21759 => x"FF",
		22783 => x"FF",
		23807 => x"FF",
		168191 => x"FF",
		169215 => x"FF",
		170239 => x"FF",
		171263 => x"FF",
		172287 => x"FF",
		316671 => x"FF",
		317695 => x"FF",
		318719 => x"FF",
		319743 => x"FF",
		320767 => x"FF",
		465151 => x"FF",
		466175 => x"FF",
		467199 => x"FF",
		468223 => x"FF",
		469247 => x"FF",
		19712 => x"FF",
		20736 => x"FF",
		21760 => x"FF",
		22784 => x"FF",
		23808 => x"FF",
		168192 => x"FF",
		169216 => x"FF",
		170240 => x"FF",
		171264 => x"FF",
		172288 => x"FF",
		316672 => x"FF",
		317696 => x"FF",
		318720 => x"FF",
		319744 => x"FF",
		320768 => x"FF",
		465152 => x"FF",
		466176 => x"FF",
		467200 => x"FF",
		468224 => x"FF",
		469248 => x"FF",
		19713 => x"FF",
		20737 => x"FF",
		21761 => x"FF",
		22785 => x"FF",
		23809 => x"FF",
		168193 => x"FF",
		169217 => x"FF",
		170241 => x"FF",
		171265 => x"FF",
		172289 => x"FF",
		316673 => x"FF",
		317697 => x"FF",
		318721 => x"FF",
		319745 => x"FF",
		320769 => x"FF",
		465153 => x"FF",
		466177 => x"FF",
		467201 => x"FF",
		468225 => x"FF",
		469249 => x"FF",
		19714 => x"FF",
		20738 => x"FF",
		21762 => x"FF",
		22786 => x"FF",
		23810 => x"FF",
		168194 => x"FF",
		169218 => x"FF",
		170242 => x"FF",
		171266 => x"FF",
		172290 => x"FF",
		316674 => x"FF",
		317698 => x"FF",
		318722 => x"FF",
		319746 => x"FF",
		320770 => x"FF",
		465154 => x"FF",
		466178 => x"FF",
		467202 => x"FF",
		468226 => x"FF",
		469250 => x"FF",
		19715 => x"FF",
		20739 => x"FF",
		21763 => x"FF",
		22787 => x"FF",
		23811 => x"FF",
		168195 => x"FF",
		169219 => x"FF",
		170243 => x"FF",
		171267 => x"FF",
		172291 => x"FF",
		316675 => x"FF",
		317699 => x"FF",
		318723 => x"FF",
		319747 => x"FF",
		320771 => x"FF",
		465155 => x"FF",
		466179 => x"FF",
		467203 => x"FF",
		468227 => x"FF",
		469251 => x"FF",
		19716 => x"FF",
		20740 => x"FF",
		21764 => x"FF",
		22788 => x"FF",
		23812 => x"FF",
		168196 => x"FF",
		169220 => x"FF",
		170244 => x"FF",
		171268 => x"FF",
		172292 => x"FF",
		316676 => x"FF",
		317700 => x"FF",
		318724 => x"FF",
		319748 => x"FF",
		320772 => x"FF",
		465156 => x"FF",
		466180 => x"FF",
		467204 => x"FF",
		468228 => x"FF",
		469252 => x"FF",
		19717 => x"FF",
		20741 => x"FF",
		21765 => x"FF",
		22789 => x"FF",
		23813 => x"FF",
		168197 => x"FF",
		169221 => x"FF",
		170245 => x"FF",
		171269 => x"FF",
		172293 => x"FF",
		316677 => x"FF",
		317701 => x"FF",
		318725 => x"FF",
		319749 => x"FF",
		320773 => x"FF",
		465157 => x"FF",
		466181 => x"FF",
		467205 => x"FF",
		468229 => x"FF",
		469253 => x"FF",
		19718 => x"FF",
		20742 => x"FF",
		21766 => x"FF",
		22790 => x"FF",
		23814 => x"FF",
		168198 => x"FF",
		169222 => x"FF",
		170246 => x"FF",
		171270 => x"FF",
		172294 => x"FF",
		316678 => x"FF",
		317702 => x"FF",
		318726 => x"FF",
		319750 => x"FF",
		320774 => x"FF",
		465158 => x"FF",
		466182 => x"FF",
		467206 => x"FF",
		468230 => x"FF",
		469254 => x"FF",
		19719 => x"FF",
		20743 => x"FF",
		21767 => x"FF",
		22791 => x"FF",
		23815 => x"FF",
		168199 => x"FF",
		169223 => x"FF",
		170247 => x"FF",
		171271 => x"FF",
		172295 => x"FF",
		316679 => x"FF",
		317703 => x"FF",
		318727 => x"FF",
		319751 => x"FF",
		320775 => x"FF",
		465159 => x"FF",
		466183 => x"FF",
		467207 => x"FF",
		468231 => x"FF",
		469255 => x"FF",
		19720 => x"FF",
		20744 => x"FF",
		21768 => x"FF",
		22792 => x"FF",
		23816 => x"FF",
		168200 => x"FF",
		169224 => x"FF",
		170248 => x"FF",
		171272 => x"FF",
		172296 => x"FF",
		316680 => x"FF",
		317704 => x"FF",
		318728 => x"FF",
		319752 => x"FF",
		320776 => x"FF",
		465160 => x"FF",
		466184 => x"FF",
		467208 => x"FF",
		468232 => x"FF",
		469256 => x"FF",
		19721 => x"FF",
		20745 => x"FF",
		21769 => x"FF",
		22793 => x"FF",
		23817 => x"FF",
		168201 => x"FF",
		169225 => x"FF",
		170249 => x"FF",
		171273 => x"FF",
		172297 => x"FF",
		316681 => x"FF",
		317705 => x"FF",
		318729 => x"FF",
		319753 => x"FF",
		320777 => x"FF",
		465161 => x"FF",
		466185 => x"FF",
		467209 => x"FF",
		468233 => x"FF",
		469257 => x"FF",
		19722 => x"FF",
		20746 => x"FF",
		21770 => x"FF",
		22794 => x"FF",
		23818 => x"FF",
		168202 => x"FF",
		169226 => x"FF",
		170250 => x"FF",
		171274 => x"FF",
		172298 => x"FF",
		316682 => x"FF",
		317706 => x"FF",
		318730 => x"FF",
		319754 => x"FF",
		320778 => x"FF",
		465162 => x"FF",
		466186 => x"FF",
		467210 => x"FF",
		468234 => x"FF",
		469258 => x"FF",
		19723 => x"FF",
		20747 => x"FF",
		21771 => x"FF",
		22795 => x"FF",
		23819 => x"FF",
		168203 => x"FF",
		169227 => x"FF",
		170251 => x"FF",
		171275 => x"FF",
		172299 => x"FF",
		316683 => x"FF",
		317707 => x"FF",
		318731 => x"FF",
		319755 => x"FF",
		320779 => x"FF",
		465163 => x"FF",
		466187 => x"FF",
		467211 => x"FF",
		468235 => x"FF",
		469259 => x"FF",
		19724 => x"FF",
		20748 => x"FF",
		21772 => x"FF",
		22796 => x"FF",
		23820 => x"FF",
		168204 => x"FF",
		169228 => x"FF",
		170252 => x"FF",
		171276 => x"FF",
		172300 => x"FF",
		316684 => x"FF",
		317708 => x"FF",
		318732 => x"FF",
		319756 => x"FF",
		320780 => x"FF",
		465164 => x"FF",
		466188 => x"FF",
		467212 => x"FF",
		468236 => x"FF",
		469260 => x"FF",
		19725 => x"FF",
		20749 => x"FF",
		21773 => x"FF",
		22797 => x"FF",
		23821 => x"FF",
		168205 => x"FF",
		169229 => x"FF",
		170253 => x"FF",
		171277 => x"FF",
		172301 => x"FF",
		316685 => x"FF",
		317709 => x"FF",
		318733 => x"FF",
		319757 => x"FF",
		320781 => x"FF",
		465165 => x"FF",
		466189 => x"FF",
		467213 => x"FF",
		468237 => x"FF",
		469261 => x"FF",
		19726 => x"FF",
		20750 => x"FF",
		21774 => x"FF",
		22798 => x"FF",
		23822 => x"FF",
		168206 => x"FF",
		169230 => x"FF",
		170254 => x"FF",
		171278 => x"FF",
		172302 => x"FF",
		316686 => x"FF",
		317710 => x"FF",
		318734 => x"FF",
		319758 => x"FF",
		320782 => x"FF",
		465166 => x"FF",
		466190 => x"FF",
		467214 => x"FF",
		468238 => x"FF",
		469262 => x"FF",
		19727 => x"FF",
		20751 => x"FF",
		21775 => x"FF",
		22799 => x"FF",
		23823 => x"FF",
		168207 => x"FF",
		169231 => x"FF",
		170255 => x"FF",
		171279 => x"FF",
		172303 => x"FF",
		316687 => x"FF",
		317711 => x"FF",
		318735 => x"FF",
		319759 => x"FF",
		320783 => x"FF",
		465167 => x"FF",
		466191 => x"FF",
		467215 => x"FF",
		468239 => x"FF",
		469263 => x"FF",
		19728 => x"FF",
		20752 => x"FF",
		21776 => x"FF",
		22800 => x"FF",
		23824 => x"FF",
		168208 => x"FF",
		169232 => x"FF",
		170256 => x"FF",
		171280 => x"FF",
		172304 => x"FF",
		316688 => x"FF",
		317712 => x"FF",
		318736 => x"FF",
		319760 => x"FF",
		320784 => x"FF",
		465168 => x"FF",
		466192 => x"FF",
		467216 => x"FF",
		468240 => x"FF",
		469264 => x"FF",
		19729 => x"FF",
		20753 => x"FF",
		21777 => x"FF",
		22801 => x"FF",
		23825 => x"FF",
		168209 => x"FF",
		169233 => x"FF",
		170257 => x"FF",
		171281 => x"FF",
		172305 => x"FF",
		316689 => x"FF",
		317713 => x"FF",
		318737 => x"FF",
		319761 => x"FF",
		320785 => x"FF",
		465169 => x"FF",
		466193 => x"FF",
		467217 => x"FF",
		468241 => x"FF",
		469265 => x"FF",
		19730 => x"FF",
		20754 => x"FF",
		21778 => x"FF",
		22802 => x"FF",
		23826 => x"FF",
		168210 => x"FF",
		169234 => x"FF",
		170258 => x"FF",
		171282 => x"FF",
		172306 => x"FF",
		316690 => x"FF",
		317714 => x"FF",
		318738 => x"FF",
		319762 => x"FF",
		320786 => x"FF",
		465170 => x"FF",
		466194 => x"FF",
		467218 => x"FF",
		468242 => x"FF",
		469266 => x"FF",
		19731 => x"FF",
		20755 => x"FF",
		21779 => x"FF",
		22803 => x"FF",
		23827 => x"FF",
		168211 => x"FF",
		169235 => x"FF",
		170259 => x"FF",
		171283 => x"FF",
		172307 => x"FF",
		316691 => x"FF",
		317715 => x"FF",
		318739 => x"FF",
		319763 => x"FF",
		320787 => x"FF",
		465171 => x"FF",
		466195 => x"FF",
		467219 => x"FF",
		468243 => x"FF",
		469267 => x"FF",
		19732 => x"FF",
		20756 => x"FF",
		21780 => x"FF",
		22804 => x"FF",
		23828 => x"FF",
		168212 => x"FF",
		169236 => x"FF",
		170260 => x"FF",
		171284 => x"FF",
		172308 => x"FF",
		316692 => x"FF",
		317716 => x"FF",
		318740 => x"FF",
		319764 => x"FF",
		320788 => x"FF",
		465172 => x"FF",
		466196 => x"FF",
		467220 => x"FF",
		468244 => x"FF",
		469268 => x"FF",
		19733 => x"FF",
		20757 => x"FF",
		21781 => x"FF",
		22805 => x"FF",
		23829 => x"FF",
		168213 => x"FF",
		169237 => x"FF",
		170261 => x"FF",
		171285 => x"FF",
		172309 => x"FF",
		316693 => x"FF",
		317717 => x"FF",
		318741 => x"FF",
		319765 => x"FF",
		320789 => x"FF",
		465173 => x"FF",
		466197 => x"FF",
		467221 => x"FF",
		468245 => x"FF",
		469269 => x"FF",
		19734 => x"FF",
		20758 => x"FF",
		21782 => x"FF",
		22806 => x"FF",
		23830 => x"FF",
		168214 => x"FF",
		169238 => x"FF",
		170262 => x"FF",
		171286 => x"FF",
		172310 => x"FF",
		316694 => x"FF",
		317718 => x"FF",
		318742 => x"FF",
		319766 => x"FF",
		320790 => x"FF",
		465174 => x"FF",
		466198 => x"FF",
		467222 => x"FF",
		468246 => x"FF",
		469270 => x"FF",
		19735 => x"FF",
		20759 => x"FF",
		21783 => x"FF",
		22807 => x"FF",
		23831 => x"FF",
		168215 => x"FF",
		169239 => x"FF",
		170263 => x"FF",
		171287 => x"FF",
		172311 => x"FF",
		316695 => x"FF",
		317719 => x"FF",
		318743 => x"FF",
		319767 => x"FF",
		320791 => x"FF",
		465175 => x"FF",
		466199 => x"FF",
		467223 => x"FF",
		468247 => x"FF",
		469271 => x"FF",
		19736 => x"FF",
		20760 => x"FF",
		21784 => x"FF",
		22808 => x"FF",
		23832 => x"FF",
		168216 => x"FF",
		169240 => x"FF",
		170264 => x"FF",
		171288 => x"FF",
		172312 => x"FF",
		316696 => x"FF",
		317720 => x"FF",
		318744 => x"FF",
		319768 => x"FF",
		320792 => x"FF",
		465176 => x"FF",
		466200 => x"FF",
		467224 => x"FF",
		468248 => x"FF",
		469272 => x"FF",
		19737 => x"FF",
		20761 => x"FF",
		21785 => x"FF",
		22809 => x"FF",
		23833 => x"FF",
		168217 => x"FF",
		169241 => x"FF",
		170265 => x"FF",
		171289 => x"FF",
		172313 => x"FF",
		316697 => x"FF",
		317721 => x"FF",
		318745 => x"FF",
		319769 => x"FF",
		320793 => x"FF",
		465177 => x"FF",
		466201 => x"FF",
		467225 => x"FF",
		468249 => x"FF",
		469273 => x"FF",
		19738 => x"FF",
		20762 => x"FF",
		21786 => x"FF",
		22810 => x"FF",
		23834 => x"FF",
		168218 => x"FF",
		169242 => x"FF",
		170266 => x"FF",
		171290 => x"FF",
		172314 => x"FF",
		316698 => x"FF",
		317722 => x"FF",
		318746 => x"FF",
		319770 => x"FF",
		320794 => x"FF",
		465178 => x"FF",
		466202 => x"FF",
		467226 => x"FF",
		468250 => x"FF",
		469274 => x"FF",
		19739 => x"FF",
		20763 => x"FF",
		21787 => x"FF",
		22811 => x"FF",
		23835 => x"FF",
		168219 => x"FF",
		169243 => x"FF",
		170267 => x"FF",
		171291 => x"FF",
		172315 => x"FF",
		316699 => x"FF",
		317723 => x"FF",
		318747 => x"FF",
		319771 => x"FF",
		320795 => x"FF",
		465179 => x"FF",
		466203 => x"FF",
		467227 => x"FF",
		468251 => x"FF",
		469275 => x"FF",
		19740 => x"FF",
		20764 => x"FF",
		21788 => x"FF",
		22812 => x"FF",
		23836 => x"FF",
		168220 => x"FF",
		169244 => x"FF",
		170268 => x"FF",
		171292 => x"FF",
		172316 => x"FF",
		316700 => x"FF",
		317724 => x"FF",
		318748 => x"FF",
		319772 => x"FF",
		320796 => x"FF",
		465180 => x"FF",
		466204 => x"FF",
		467228 => x"FF",
		468252 => x"FF",
		469276 => x"FF",
		19741 => x"FF",
		20765 => x"FF",
		21789 => x"FF",
		22813 => x"FF",
		23837 => x"FF",
		168221 => x"FF",
		169245 => x"FF",
		170269 => x"FF",
		171293 => x"FF",
		172317 => x"FF",
		316701 => x"FF",
		317725 => x"FF",
		318749 => x"FF",
		319773 => x"FF",
		320797 => x"FF",
		465181 => x"FF",
		466205 => x"FF",
		467229 => x"FF",
		468253 => x"FF",
		469277 => x"FF",
		19742 => x"FF",
		20766 => x"FF",
		21790 => x"FF",
		22814 => x"FF",
		23838 => x"FF",
		168222 => x"FF",
		169246 => x"FF",
		170270 => x"FF",
		171294 => x"FF",
		172318 => x"FF",
		316702 => x"FF",
		317726 => x"FF",
		318750 => x"FF",
		319774 => x"FF",
		320798 => x"FF",
		465182 => x"FF",
		466206 => x"FF",
		467230 => x"FF",
		468254 => x"FF",
		469278 => x"FF",
		19743 => x"FF",
		20767 => x"FF",
		21791 => x"FF",
		22815 => x"FF",
		23839 => x"FF",
		168223 => x"FF",
		169247 => x"FF",
		170271 => x"FF",
		171295 => x"FF",
		172319 => x"FF",
		316703 => x"FF",
		317727 => x"FF",
		318751 => x"FF",
		319775 => x"FF",
		320799 => x"FF",
		465183 => x"FF",
		466207 => x"FF",
		467231 => x"FF",
		468255 => x"FF",
		469279 => x"FF",
		19744 => x"FF",
		20768 => x"FF",
		21792 => x"FF",
		22816 => x"FF",
		23840 => x"FF",
		168224 => x"FF",
		169248 => x"FF",
		170272 => x"FF",
		171296 => x"FF",
		172320 => x"FF",
		316704 => x"FF",
		317728 => x"FF",
		318752 => x"FF",
		319776 => x"FF",
		320800 => x"FF",
		465184 => x"FF",
		466208 => x"FF",
		467232 => x"FF",
		468256 => x"FF",
		469280 => x"FF",
		19745 => x"FF",
		20769 => x"FF",
		21793 => x"FF",
		22817 => x"FF",
		23841 => x"FF",
		168225 => x"FF",
		169249 => x"FF",
		170273 => x"FF",
		171297 => x"FF",
		172321 => x"FF",
		316705 => x"FF",
		317729 => x"FF",
		318753 => x"FF",
		319777 => x"FF",
		320801 => x"FF",
		465185 => x"FF",
		466209 => x"FF",
		467233 => x"FF",
		468257 => x"FF",
		469281 => x"FF",
		19746 => x"FF",
		20770 => x"FF",
		21794 => x"FF",
		22818 => x"FF",
		23842 => x"FF",
		168226 => x"FF",
		169250 => x"FF",
		170274 => x"FF",
		171298 => x"FF",
		172322 => x"FF",
		316706 => x"FF",
		317730 => x"FF",
		318754 => x"FF",
		319778 => x"FF",
		320802 => x"FF",
		465186 => x"FF",
		466210 => x"FF",
		467234 => x"FF",
		468258 => x"FF",
		469282 => x"FF",
		19747 => x"FF",
		20771 => x"FF",
		21795 => x"FF",
		22819 => x"FF",
		23843 => x"FF",
		168227 => x"FF",
		169251 => x"FF",
		170275 => x"FF",
		171299 => x"FF",
		172323 => x"FF",
		316707 => x"FF",
		317731 => x"FF",
		318755 => x"FF",
		319779 => x"FF",
		320803 => x"FF",
		465187 => x"FF",
		466211 => x"FF",
		467235 => x"FF",
		468259 => x"FF",
		469283 => x"FF",
		19748 => x"FF",
		20772 => x"FF",
		21796 => x"FF",
		22820 => x"FF",
		23844 => x"FF",
		168228 => x"FF",
		169252 => x"FF",
		170276 => x"FF",
		171300 => x"FF",
		172324 => x"FF",
		316708 => x"FF",
		317732 => x"FF",
		318756 => x"FF",
		319780 => x"FF",
		320804 => x"FF",
		465188 => x"FF",
		466212 => x"FF",
		467236 => x"FF",
		468260 => x"FF",
		469284 => x"FF",
		19749 => x"FF",
		20773 => x"FF",
		21797 => x"FF",
		22821 => x"FF",
		23845 => x"FF",
		168229 => x"FF",
		169253 => x"FF",
		170277 => x"FF",
		171301 => x"FF",
		172325 => x"FF",
		316709 => x"FF",
		317733 => x"FF",
		318757 => x"FF",
		319781 => x"FF",
		320805 => x"FF",
		465189 => x"FF",
		466213 => x"FF",
		467237 => x"FF",
		468261 => x"FF",
		469285 => x"FF",
		19750 => x"FF",
		20774 => x"FF",
		21798 => x"FF",
		22822 => x"FF",
		23846 => x"FF",
		168230 => x"FF",
		169254 => x"FF",
		170278 => x"FF",
		171302 => x"FF",
		172326 => x"FF",
		316710 => x"FF",
		317734 => x"FF",
		318758 => x"FF",
		319782 => x"FF",
		320806 => x"FF",
		465190 => x"FF",
		466214 => x"FF",
		467238 => x"FF",
		468262 => x"FF",
		469286 => x"FF",
		19751 => x"FF",
		20775 => x"FF",
		21799 => x"FF",
		22823 => x"FF",
		23847 => x"FF",
		168231 => x"FF",
		169255 => x"FF",
		170279 => x"FF",
		171303 => x"FF",
		172327 => x"FF",
		316711 => x"FF",
		317735 => x"FF",
		318759 => x"FF",
		319783 => x"FF",
		320807 => x"FF",
		465191 => x"FF",
		466215 => x"FF",
		467239 => x"FF",
		468263 => x"FF",
		469287 => x"FF",
		19752 => x"FF",
		20776 => x"FF",
		21800 => x"FF",
		22824 => x"FF",
		23848 => x"FF",
		168232 => x"FF",
		169256 => x"FF",
		170280 => x"FF",
		171304 => x"FF",
		172328 => x"FF",
		316712 => x"FF",
		317736 => x"FF",
		318760 => x"FF",
		319784 => x"FF",
		320808 => x"FF",
		465192 => x"FF",
		466216 => x"FF",
		467240 => x"FF",
		468264 => x"FF",
		469288 => x"FF",
		19753 => x"FF",
		20777 => x"FF",
		21801 => x"FF",
		22825 => x"FF",
		23849 => x"FF",
		168233 => x"FF",
		169257 => x"FF",
		170281 => x"FF",
		171305 => x"FF",
		172329 => x"FF",
		316713 => x"FF",
		317737 => x"FF",
		318761 => x"FF",
		319785 => x"FF",
		320809 => x"FF",
		465193 => x"FF",
		466217 => x"FF",
		467241 => x"FF",
		468265 => x"FF",
		469289 => x"FF",
		19754 => x"FF",
		20778 => x"FF",
		21802 => x"FF",
		22826 => x"FF",
		23850 => x"FF",
		168234 => x"FF",
		169258 => x"FF",
		170282 => x"FF",
		171306 => x"FF",
		172330 => x"FF",
		316714 => x"FF",
		317738 => x"FF",
		318762 => x"FF",
		319786 => x"FF",
		320810 => x"FF",
		465194 => x"FF",
		466218 => x"FF",
		467242 => x"FF",
		468266 => x"FF",
		469290 => x"FF",
		19755 => x"FF",
		20779 => x"FF",
		21803 => x"FF",
		22827 => x"FF",
		23851 => x"FF",
		168235 => x"FF",
		169259 => x"FF",
		170283 => x"FF",
		171307 => x"FF",
		172331 => x"FF",
		316715 => x"FF",
		317739 => x"FF",
		318763 => x"FF",
		319787 => x"FF",
		320811 => x"FF",
		465195 => x"FF",
		466219 => x"FF",
		467243 => x"FF",
		468267 => x"FF",
		469291 => x"FF",
		19756 => x"FF",
		20780 => x"FF",
		21804 => x"FF",
		22828 => x"FF",
		23852 => x"FF",
		168236 => x"FF",
		169260 => x"FF",
		170284 => x"FF",
		171308 => x"FF",
		172332 => x"FF",
		316716 => x"FF",
		317740 => x"FF",
		318764 => x"FF",
		319788 => x"FF",
		320812 => x"FF",
		465196 => x"FF",
		466220 => x"FF",
		467244 => x"FF",
		468268 => x"FF",
		469292 => x"FF",
		19757 => x"FF",
		20781 => x"FF",
		21805 => x"FF",
		22829 => x"FF",
		23853 => x"FF",
		168237 => x"FF",
		169261 => x"FF",
		170285 => x"FF",
		171309 => x"FF",
		172333 => x"FF",
		316717 => x"FF",
		317741 => x"FF",
		318765 => x"FF",
		319789 => x"FF",
		320813 => x"FF",
		465197 => x"FF",
		466221 => x"FF",
		467245 => x"FF",
		468269 => x"FF",
		469293 => x"FF",
		19758 => x"FF",
		20782 => x"FF",
		21806 => x"FF",
		22830 => x"FF",
		23854 => x"FF",
		168238 => x"FF",
		169262 => x"FF",
		170286 => x"FF",
		171310 => x"FF",
		172334 => x"FF",
		316718 => x"FF",
		317742 => x"FF",
		318766 => x"FF",
		319790 => x"FF",
		320814 => x"FF",
		465198 => x"FF",
		466222 => x"FF",
		467246 => x"FF",
		468270 => x"FF",
		469294 => x"FF",
		19759 => x"FF",
		20783 => x"FF",
		21807 => x"FF",
		22831 => x"FF",
		23855 => x"FF",
		168239 => x"FF",
		169263 => x"FF",
		170287 => x"FF",
		171311 => x"FF",
		172335 => x"FF",
		316719 => x"FF",
		317743 => x"FF",
		318767 => x"FF",
		319791 => x"FF",
		320815 => x"FF",
		465199 => x"FF",
		466223 => x"FF",
		467247 => x"FF",
		468271 => x"FF",
		469295 => x"FF",
		19760 => x"FF",
		20784 => x"FF",
		21808 => x"FF",
		22832 => x"FF",
		23856 => x"FF",
		168240 => x"FF",
		169264 => x"FF",
		170288 => x"FF",
		171312 => x"FF",
		172336 => x"FF",
		316720 => x"FF",
		317744 => x"FF",
		318768 => x"FF",
		319792 => x"FF",
		320816 => x"FF",
		465200 => x"FF",
		466224 => x"FF",
		467248 => x"FF",
		468272 => x"FF",
		469296 => x"FF",
		19761 => x"FF",
		20785 => x"FF",
		21809 => x"FF",
		22833 => x"FF",
		23857 => x"FF",
		168241 => x"FF",
		169265 => x"FF",
		170289 => x"FF",
		171313 => x"FF",
		172337 => x"FF",
		316721 => x"FF",
		317745 => x"FF",
		318769 => x"FF",
		319793 => x"FF",
		320817 => x"FF",
		465201 => x"FF",
		466225 => x"FF",
		467249 => x"FF",
		468273 => x"FF",
		469297 => x"FF",
		19762 => x"FF",
		20786 => x"FF",
		21810 => x"FF",
		22834 => x"FF",
		23858 => x"FF",
		168242 => x"FF",
		169266 => x"FF",
		170290 => x"FF",
		171314 => x"FF",
		172338 => x"FF",
		316722 => x"FF",
		317746 => x"FF",
		318770 => x"FF",
		319794 => x"FF",
		320818 => x"FF",
		465202 => x"FF",
		466226 => x"FF",
		467250 => x"FF",
		468274 => x"FF",
		469298 => x"FF",
		19763 => x"FF",
		20787 => x"FF",
		21811 => x"FF",
		22835 => x"FF",
		23859 => x"FF",
		168243 => x"FF",
		169267 => x"FF",
		170291 => x"FF",
		171315 => x"FF",
		172339 => x"FF",
		316723 => x"FF",
		317747 => x"FF",
		318771 => x"FF",
		319795 => x"FF",
		320819 => x"FF",
		465203 => x"FF",
		466227 => x"FF",
		467251 => x"FF",
		468275 => x"FF",
		469299 => x"FF",
		19764 => x"FF",
		20788 => x"FF",
		21812 => x"FF",
		22836 => x"FF",
		23860 => x"FF",
		168244 => x"FF",
		169268 => x"FF",
		170292 => x"FF",
		171316 => x"FF",
		172340 => x"FF",
		316724 => x"FF",
		317748 => x"FF",
		318772 => x"FF",
		319796 => x"FF",
		320820 => x"FF",
		465204 => x"FF",
		466228 => x"FF",
		467252 => x"FF",
		468276 => x"FF",
		469300 => x"FF",
		19765 => x"FF",
		20789 => x"FF",
		21813 => x"FF",
		22837 => x"FF",
		23861 => x"FF",
		168245 => x"FF",
		169269 => x"FF",
		170293 => x"FF",
		171317 => x"FF",
		172341 => x"FF",
		316725 => x"FF",
		317749 => x"FF",
		318773 => x"FF",
		319797 => x"FF",
		320821 => x"FF",
		465205 => x"FF",
		466229 => x"FF",
		467253 => x"FF",
		468277 => x"FF",
		469301 => x"FF",
		19766 => x"FF",
		20790 => x"FF",
		21814 => x"FF",
		22838 => x"FF",
		23862 => x"FF",
		168246 => x"FF",
		169270 => x"FF",
		170294 => x"FF",
		171318 => x"FF",
		172342 => x"FF",
		316726 => x"FF",
		317750 => x"FF",
		318774 => x"FF",
		319798 => x"FF",
		320822 => x"FF",
		465206 => x"FF",
		466230 => x"FF",
		467254 => x"FF",
		468278 => x"FF",
		469302 => x"FF",
		19767 => x"FF",
		20791 => x"FF",
		21815 => x"FF",
		22839 => x"FF",
		23863 => x"FF",
		168247 => x"FF",
		169271 => x"FF",
		170295 => x"FF",
		171319 => x"FF",
		172343 => x"FF",
		316727 => x"FF",
		317751 => x"FF",
		318775 => x"FF",
		319799 => x"FF",
		320823 => x"FF",
		465207 => x"FF",
		466231 => x"FF",
		467255 => x"FF",
		468279 => x"FF",
		469303 => x"FF",
		19768 => x"FF",
		20792 => x"FF",
		21816 => x"FF",
		22840 => x"FF",
		23864 => x"FF",
		168248 => x"FF",
		169272 => x"FF",
		170296 => x"FF",
		171320 => x"FF",
		172344 => x"FF",
		316728 => x"FF",
		317752 => x"FF",
		318776 => x"FF",
		319800 => x"FF",
		320824 => x"FF",
		465208 => x"FF",
		466232 => x"FF",
		467256 => x"FF",
		468280 => x"FF",
		469304 => x"FF",
		19769 => x"FF",
		20793 => x"FF",
		21817 => x"FF",
		22841 => x"FF",
		23865 => x"FF",
		168249 => x"FF",
		169273 => x"FF",
		170297 => x"FF",
		171321 => x"FF",
		172345 => x"FF",
		316729 => x"FF",
		317753 => x"FF",
		318777 => x"FF",
		319801 => x"FF",
		320825 => x"FF",
		465209 => x"FF",
		466233 => x"FF",
		467257 => x"FF",
		468281 => x"FF",
		469305 => x"FF",
		19770 => x"FF",
		20794 => x"FF",
		21818 => x"FF",
		22842 => x"FF",
		23866 => x"FF",
		168250 => x"FF",
		169274 => x"FF",
		170298 => x"FF",
		171322 => x"FF",
		172346 => x"FF",
		316730 => x"FF",
		317754 => x"FF",
		318778 => x"FF",
		319802 => x"FF",
		320826 => x"FF",
		465210 => x"FF",
		466234 => x"FF",
		467258 => x"FF",
		468282 => x"FF",
		469306 => x"FF",
		19771 => x"FF",
		20795 => x"FF",
		21819 => x"FF",
		22843 => x"FF",
		23867 => x"FF",
		168251 => x"FF",
		169275 => x"FF",
		170299 => x"FF",
		171323 => x"FF",
		172347 => x"FF",
		316731 => x"FF",
		317755 => x"FF",
		318779 => x"FF",
		319803 => x"FF",
		320827 => x"FF",
		465211 => x"FF",
		466235 => x"FF",
		467259 => x"FF",
		468283 => x"FF",
		469307 => x"FF",
		19772 => x"FF",
		20796 => x"FF",
		21820 => x"FF",
		22844 => x"FF",
		23868 => x"FF",
		168252 => x"FF",
		169276 => x"FF",
		170300 => x"FF",
		171324 => x"FF",
		172348 => x"FF",
		316732 => x"FF",
		317756 => x"FF",
		318780 => x"FF",
		319804 => x"FF",
		320828 => x"FF",
		465212 => x"FF",
		466236 => x"FF",
		467260 => x"FF",
		468284 => x"FF",
		469308 => x"FF",
		19773 => x"FF",
		20797 => x"FF",
		21821 => x"FF",
		22845 => x"FF",
		23869 => x"FF",
		168253 => x"FF",
		169277 => x"FF",
		170301 => x"FF",
		171325 => x"FF",
		172349 => x"FF",
		316733 => x"FF",
		317757 => x"FF",
		318781 => x"FF",
		319805 => x"FF",
		320829 => x"FF",
		465213 => x"FF",
		466237 => x"FF",
		467261 => x"FF",
		468285 => x"FF",
		469309 => x"FF",
		19774 => x"FF",
		20798 => x"FF",
		21822 => x"FF",
		22846 => x"FF",
		23870 => x"FF",
		168254 => x"FF",
		169278 => x"FF",
		170302 => x"FF",
		171326 => x"FF",
		172350 => x"FF",
		316734 => x"FF",
		317758 => x"FF",
		318782 => x"FF",
		319806 => x"FF",
		320830 => x"FF",
		465214 => x"FF",
		466238 => x"FF",
		467262 => x"FF",
		468286 => x"FF",
		469310 => x"FF",
		19775 => x"FF",
		20799 => x"FF",
		21823 => x"FF",
		22847 => x"FF",
		23871 => x"FF",
		168255 => x"FF",
		169279 => x"FF",
		170303 => x"FF",
		171327 => x"FF",
		172351 => x"FF",
		316735 => x"FF",
		317759 => x"FF",
		318783 => x"FF",
		319807 => x"FF",
		320831 => x"FF",
		465215 => x"FF",
		466239 => x"FF",
		467263 => x"FF",
		468287 => x"FF",
		469311 => x"FF",
		19776 => x"FF",
		20800 => x"FF",
		21824 => x"FF",
		22848 => x"FF",
		23872 => x"FF",
		168256 => x"FF",
		169280 => x"FF",
		170304 => x"FF",
		171328 => x"FF",
		172352 => x"FF",
		316736 => x"FF",
		317760 => x"FF",
		318784 => x"FF",
		319808 => x"FF",
		320832 => x"FF",
		465216 => x"FF",
		466240 => x"FF",
		467264 => x"FF",
		468288 => x"FF",
		469312 => x"FF",
		19777 => x"FF",
		20801 => x"FF",
		21825 => x"FF",
		22849 => x"FF",
		23873 => x"FF",
		168257 => x"FF",
		169281 => x"FF",
		170305 => x"FF",
		171329 => x"FF",
		172353 => x"FF",
		316737 => x"FF",
		317761 => x"FF",
		318785 => x"FF",
		319809 => x"FF",
		320833 => x"FF",
		465217 => x"FF",
		466241 => x"FF",
		467265 => x"FF",
		468289 => x"FF",
		469313 => x"FF",
		19778 => x"FF",
		20802 => x"FF",
		21826 => x"FF",
		22850 => x"FF",
		23874 => x"FF",
		168258 => x"FF",
		169282 => x"FF",
		170306 => x"FF",
		171330 => x"FF",
		172354 => x"FF",
		316738 => x"FF",
		317762 => x"FF",
		318786 => x"FF",
		319810 => x"FF",
		320834 => x"FF",
		465218 => x"FF",
		466242 => x"FF",
		467266 => x"FF",
		468290 => x"FF",
		469314 => x"FF",
		19779 => x"FF",
		20803 => x"FF",
		21827 => x"FF",
		22851 => x"FF",
		23875 => x"FF",
		168259 => x"FF",
		169283 => x"FF",
		170307 => x"FF",
		171331 => x"FF",
		172355 => x"FF",
		316739 => x"FF",
		317763 => x"FF",
		318787 => x"FF",
		319811 => x"FF",
		320835 => x"FF",
		465219 => x"FF",
		466243 => x"FF",
		467267 => x"FF",
		468291 => x"FF",
		469315 => x"FF",
		19780 => x"FF",
		20804 => x"FF",
		21828 => x"FF",
		22852 => x"FF",
		23876 => x"FF",
		168260 => x"FF",
		169284 => x"FF",
		170308 => x"FF",
		171332 => x"FF",
		172356 => x"FF",
		316740 => x"FF",
		317764 => x"FF",
		318788 => x"FF",
		319812 => x"FF",
		320836 => x"FF",
		465220 => x"FF",
		466244 => x"FF",
		467268 => x"FF",
		468292 => x"FF",
		469316 => x"FF",
		19781 => x"FF",
		20805 => x"FF",
		21829 => x"FF",
		22853 => x"FF",
		23877 => x"FF",
		168261 => x"FF",
		169285 => x"FF",
		170309 => x"FF",
		171333 => x"FF",
		172357 => x"FF",
		316741 => x"FF",
		317765 => x"FF",
		318789 => x"FF",
		319813 => x"FF",
		320837 => x"FF",
		465221 => x"FF",
		466245 => x"FF",
		467269 => x"FF",
		468293 => x"FF",
		469317 => x"FF",
		19782 => x"FF",
		20806 => x"FF",
		21830 => x"FF",
		22854 => x"FF",
		23878 => x"FF",
		168262 => x"FF",
		169286 => x"FF",
		170310 => x"FF",
		171334 => x"FF",
		172358 => x"FF",
		316742 => x"FF",
		317766 => x"FF",
		318790 => x"FF",
		319814 => x"FF",
		320838 => x"FF",
		465222 => x"FF",
		466246 => x"FF",
		467270 => x"FF",
		468294 => x"FF",
		469318 => x"FF",
		19783 => x"FF",
		20807 => x"FF",
		21831 => x"FF",
		22855 => x"FF",
		23879 => x"FF",
		168263 => x"FF",
		169287 => x"FF",
		170311 => x"FF",
		171335 => x"FF",
		172359 => x"FF",
		316743 => x"FF",
		317767 => x"FF",
		318791 => x"FF",
		319815 => x"FF",
		320839 => x"FF",
		465223 => x"FF",
		466247 => x"FF",
		467271 => x"FF",
		468295 => x"FF",
		469319 => x"FF",
		19784 => x"FF",
		20808 => x"FF",
		21832 => x"FF",
		22856 => x"FF",
		23880 => x"FF",
		168264 => x"FF",
		169288 => x"FF",
		170312 => x"FF",
		171336 => x"FF",
		172360 => x"FF",
		316744 => x"FF",
		317768 => x"FF",
		318792 => x"FF",
		319816 => x"FF",
		320840 => x"FF",
		465224 => x"FF",
		466248 => x"FF",
		467272 => x"FF",
		468296 => x"FF",
		469320 => x"FF",
		19785 => x"FF",
		20809 => x"FF",
		21833 => x"FF",
		22857 => x"FF",
		23881 => x"FF",
		168265 => x"FF",
		169289 => x"FF",
		170313 => x"FF",
		171337 => x"FF",
		172361 => x"FF",
		316745 => x"FF",
		317769 => x"FF",
		318793 => x"FF",
		319817 => x"FF",
		320841 => x"FF",
		465225 => x"FF",
		466249 => x"FF",
		467273 => x"FF",
		468297 => x"FF",
		469321 => x"FF",
		19786 => x"FF",
		20810 => x"FF",
		21834 => x"FF",
		22858 => x"FF",
		23882 => x"FF",
		168266 => x"FF",
		169290 => x"FF",
		170314 => x"FF",
		171338 => x"FF",
		172362 => x"FF",
		316746 => x"FF",
		317770 => x"FF",
		318794 => x"FF",
		319818 => x"FF",
		320842 => x"FF",
		465226 => x"FF",
		466250 => x"FF",
		467274 => x"FF",
		468298 => x"FF",
		469322 => x"FF",
		19787 => x"FF",
		20811 => x"FF",
		21835 => x"FF",
		22859 => x"FF",
		23883 => x"FF",
		168267 => x"FF",
		169291 => x"FF",
		170315 => x"FF",
		171339 => x"FF",
		172363 => x"FF",
		316747 => x"FF",
		317771 => x"FF",
		318795 => x"FF",
		319819 => x"FF",
		320843 => x"FF",
		465227 => x"FF",
		466251 => x"FF",
		467275 => x"FF",
		468299 => x"FF",
		469323 => x"FF",
		19788 => x"FF",
		20812 => x"FF",
		21836 => x"FF",
		22860 => x"FF",
		23884 => x"FF",
		168268 => x"FF",
		169292 => x"FF",
		170316 => x"FF",
		171340 => x"FF",
		172364 => x"FF",
		316748 => x"FF",
		317772 => x"FF",
		318796 => x"FF",
		319820 => x"FF",
		320844 => x"FF",
		465228 => x"FF",
		466252 => x"FF",
		467276 => x"FF",
		468300 => x"FF",
		469324 => x"FF",
		19789 => x"FF",
		20813 => x"FF",
		21837 => x"FF",
		22861 => x"FF",
		23885 => x"FF",
		168269 => x"FF",
		169293 => x"FF",
		170317 => x"FF",
		171341 => x"FF",
		172365 => x"FF",
		316749 => x"FF",
		317773 => x"FF",
		318797 => x"FF",
		319821 => x"FF",
		320845 => x"FF",
		465229 => x"FF",
		466253 => x"FF",
		467277 => x"FF",
		468301 => x"FF",
		469325 => x"FF",
		19790 => x"FF",
		20814 => x"FF",
		21838 => x"FF",
		22862 => x"FF",
		23886 => x"FF",
		168270 => x"FF",
		169294 => x"FF",
		170318 => x"FF",
		171342 => x"FF",
		172366 => x"FF",
		316750 => x"FF",
		317774 => x"FF",
		318798 => x"FF",
		319822 => x"FF",
		320846 => x"FF",
		465230 => x"FF",
		466254 => x"FF",
		467278 => x"FF",
		468302 => x"FF",
		469326 => x"FF",
		19791 => x"FF",
		20815 => x"FF",
		21839 => x"FF",
		22863 => x"FF",
		23887 => x"FF",
		168271 => x"FF",
		169295 => x"FF",
		170319 => x"FF",
		171343 => x"FF",
		172367 => x"FF",
		316751 => x"FF",
		317775 => x"FF",
		318799 => x"FF",
		319823 => x"FF",
		320847 => x"FF",
		465231 => x"FF",
		466255 => x"FF",
		467279 => x"FF",
		468303 => x"FF",
		469327 => x"FF",
		19792 => x"FF",
		20816 => x"FF",
		21840 => x"FF",
		22864 => x"FF",
		23888 => x"FF",
		168272 => x"FF",
		169296 => x"FF",
		170320 => x"FF",
		171344 => x"FF",
		172368 => x"FF",
		316752 => x"FF",
		317776 => x"FF",
		318800 => x"FF",
		319824 => x"FF",
		320848 => x"FF",
		465232 => x"FF",
		466256 => x"FF",
		467280 => x"FF",
		468304 => x"FF",
		469328 => x"FF",
		19793 => x"FF",
		20817 => x"FF",
		21841 => x"FF",
		22865 => x"FF",
		23889 => x"FF",
		168273 => x"FF",
		169297 => x"FF",
		170321 => x"FF",
		171345 => x"FF",
		172369 => x"FF",
		316753 => x"FF",
		317777 => x"FF",
		318801 => x"FF",
		319825 => x"FF",
		320849 => x"FF",
		465233 => x"FF",
		466257 => x"FF",
		467281 => x"FF",
		468305 => x"FF",
		469329 => x"FF",
		19794 => x"FF",
		20818 => x"FF",
		21842 => x"FF",
		22866 => x"FF",
		23890 => x"FF",
		168274 => x"FF",
		169298 => x"FF",
		170322 => x"FF",
		171346 => x"FF",
		172370 => x"FF",
		316754 => x"FF",
		317778 => x"FF",
		318802 => x"FF",
		319826 => x"FF",
		320850 => x"FF",
		465234 => x"FF",
		466258 => x"FF",
		467282 => x"FF",
		468306 => x"FF",
		469330 => x"FF",
		19795 => x"FF",
		20819 => x"FF",
		21843 => x"FF",
		22867 => x"FF",
		23891 => x"FF",
		168275 => x"FF",
		169299 => x"FF",
		170323 => x"FF",
		171347 => x"FF",
		172371 => x"FF",
		316755 => x"FF",
		317779 => x"FF",
		318803 => x"FF",
		319827 => x"FF",
		320851 => x"FF",
		465235 => x"FF",
		466259 => x"FF",
		467283 => x"FF",
		468307 => x"FF",
		469331 => x"FF",
		19796 => x"FF",
		20820 => x"FF",
		21844 => x"FF",
		22868 => x"FF",
		23892 => x"FF",
		168276 => x"FF",
		169300 => x"FF",
		170324 => x"FF",
		171348 => x"FF",
		172372 => x"FF",
		316756 => x"FF",
		317780 => x"FF",
		318804 => x"FF",
		319828 => x"FF",
		320852 => x"FF",
		465236 => x"FF",
		466260 => x"FF",
		467284 => x"FF",
		468308 => x"FF",
		469332 => x"FF",
		19797 => x"FF",
		20821 => x"FF",
		21845 => x"FF",
		22869 => x"FF",
		23893 => x"FF",
		168277 => x"FF",
		169301 => x"FF",
		170325 => x"FF",
		171349 => x"FF",
		172373 => x"FF",
		316757 => x"FF",
		317781 => x"FF",
		318805 => x"FF",
		319829 => x"FF",
		320853 => x"FF",
		465237 => x"FF",
		466261 => x"FF",
		467285 => x"FF",
		468309 => x"FF",
		469333 => x"FF",
		19798 => x"FF",
		20822 => x"FF",
		21846 => x"FF",
		22870 => x"FF",
		23894 => x"FF",
		168278 => x"FF",
		169302 => x"FF",
		170326 => x"FF",
		171350 => x"FF",
		172374 => x"FF",
		316758 => x"FF",
		317782 => x"FF",
		318806 => x"FF",
		319830 => x"FF",
		320854 => x"FF",
		465238 => x"FF",
		466262 => x"FF",
		467286 => x"FF",
		468310 => x"FF",
		469334 => x"FF",
		19799 => x"FF",
		20823 => x"FF",
		21847 => x"FF",
		22871 => x"FF",
		23895 => x"FF",
		168279 => x"FF",
		169303 => x"FF",
		170327 => x"FF",
		171351 => x"FF",
		172375 => x"FF",
		316759 => x"FF",
		317783 => x"FF",
		318807 => x"FF",
		319831 => x"FF",
		320855 => x"FF",
		465239 => x"FF",
		466263 => x"FF",
		467287 => x"FF",
		468311 => x"FF",
		469335 => x"FF",
		19800 => x"FF",
		20824 => x"FF",
		21848 => x"FF",
		22872 => x"FF",
		23896 => x"FF",
		168280 => x"FF",
		169304 => x"FF",
		170328 => x"FF",
		171352 => x"FF",
		172376 => x"FF",
		316760 => x"FF",
		317784 => x"FF",
		318808 => x"FF",
		319832 => x"FF",
		320856 => x"FF",
		465240 => x"FF",
		466264 => x"FF",
		467288 => x"FF",
		468312 => x"FF",
		469336 => x"FF",
		19801 => x"FF",
		20825 => x"FF",
		21849 => x"FF",
		22873 => x"FF",
		23897 => x"FF",
		168281 => x"FF",
		169305 => x"FF",
		170329 => x"FF",
		171353 => x"FF",
		172377 => x"FF",
		316761 => x"FF",
		317785 => x"FF",
		318809 => x"FF",
		319833 => x"FF",
		320857 => x"FF",
		465241 => x"FF",
		466265 => x"FF",
		467289 => x"FF",
		468313 => x"FF",
		469337 => x"FF",
		19802 => x"FF",
		20826 => x"FF",
		21850 => x"FF",
		22874 => x"FF",
		23898 => x"FF",
		168282 => x"FF",
		169306 => x"FF",
		170330 => x"FF",
		171354 => x"FF",
		172378 => x"FF",
		316762 => x"FF",
		317786 => x"FF",
		318810 => x"FF",
		319834 => x"FF",
		320858 => x"FF",
		465242 => x"FF",
		466266 => x"FF",
		467290 => x"FF",
		468314 => x"FF",
		469338 => x"FF",
		19803 => x"FF",
		20827 => x"FF",
		21851 => x"FF",
		22875 => x"FF",
		23899 => x"FF",
		168283 => x"FF",
		169307 => x"FF",
		170331 => x"FF",
		171355 => x"FF",
		172379 => x"FF",
		316763 => x"FF",
		317787 => x"FF",
		318811 => x"FF",
		319835 => x"FF",
		320859 => x"FF",
		465243 => x"FF",
		466267 => x"FF",
		467291 => x"FF",
		468315 => x"FF",
		469339 => x"FF",
		19804 => x"FF",
		20828 => x"FF",
		21852 => x"FF",
		22876 => x"FF",
		23900 => x"FF",
		168284 => x"FF",
		169308 => x"FF",
		170332 => x"FF",
		171356 => x"FF",
		172380 => x"FF",
		316764 => x"FF",
		317788 => x"FF",
		318812 => x"FF",
		319836 => x"FF",
		320860 => x"FF",
		465244 => x"FF",
		466268 => x"FF",
		467292 => x"FF",
		468316 => x"FF",
		469340 => x"FF",
		19805 => x"FF",
		20829 => x"FF",
		21853 => x"FF",
		22877 => x"FF",
		23901 => x"FF",
		168285 => x"FF",
		169309 => x"FF",
		170333 => x"FF",
		171357 => x"FF",
		172381 => x"FF",
		316765 => x"FF",
		317789 => x"FF",
		318813 => x"FF",
		319837 => x"FF",
		320861 => x"FF",
		465245 => x"FF",
		466269 => x"FF",
		467293 => x"FF",
		468317 => x"FF",
		469341 => x"FF",
		19806 => x"FF",
		20830 => x"FF",
		21854 => x"FF",
		22878 => x"FF",
		23902 => x"FF",
		168286 => x"FF",
		169310 => x"FF",
		170334 => x"FF",
		171358 => x"FF",
		172382 => x"FF",
		316766 => x"FF",
		317790 => x"FF",
		318814 => x"FF",
		319838 => x"FF",
		320862 => x"FF",
		465246 => x"FF",
		466270 => x"FF",
		467294 => x"FF",
		468318 => x"FF",
		469342 => x"FF",
		19807 => x"FF",
		20831 => x"FF",
		21855 => x"FF",
		22879 => x"FF",
		23903 => x"FF",
		168287 => x"FF",
		169311 => x"FF",
		170335 => x"FF",
		171359 => x"FF",
		172383 => x"FF",
		316767 => x"FF",
		317791 => x"FF",
		318815 => x"FF",
		319839 => x"FF",
		320863 => x"FF",
		465247 => x"FF",
		466271 => x"FF",
		467295 => x"FF",
		468319 => x"FF",
		469343 => x"FF",
		19808 => x"FF",
		20832 => x"FF",
		21856 => x"FF",
		22880 => x"FF",
		23904 => x"FF",
		168288 => x"FF",
		169312 => x"FF",
		170336 => x"FF",
		171360 => x"FF",
		172384 => x"FF",
		316768 => x"FF",
		317792 => x"FF",
		318816 => x"FF",
		319840 => x"FF",
		320864 => x"FF",
		465248 => x"FF",
		466272 => x"FF",
		467296 => x"FF",
		468320 => x"FF",
		469344 => x"FF",
		19809 => x"FF",
		20833 => x"FF",
		21857 => x"FF",
		22881 => x"FF",
		23905 => x"FF",
		168289 => x"FF",
		169313 => x"FF",
		170337 => x"FF",
		171361 => x"FF",
		172385 => x"FF",
		316769 => x"FF",
		317793 => x"FF",
		318817 => x"FF",
		319841 => x"FF",
		320865 => x"FF",
		465249 => x"FF",
		466273 => x"FF",
		467297 => x"FF",
		468321 => x"FF",
		469345 => x"FF",
		19810 => x"FF",
		20834 => x"FF",
		21858 => x"FF",
		22882 => x"FF",
		23906 => x"FF",
		168290 => x"FF",
		169314 => x"FF",
		170338 => x"FF",
		171362 => x"FF",
		172386 => x"FF",
		316770 => x"FF",
		317794 => x"FF",
		318818 => x"FF",
		319842 => x"FF",
		320866 => x"FF",
		465250 => x"FF",
		466274 => x"FF",
		467298 => x"FF",
		468322 => x"FF",
		469346 => x"FF",
		19811 => x"FF",
		20835 => x"FF",
		21859 => x"FF",
		22883 => x"FF",
		23907 => x"FF",
		168291 => x"FF",
		169315 => x"FF",
		170339 => x"FF",
		171363 => x"FF",
		172387 => x"FF",
		316771 => x"FF",
		317795 => x"FF",
		318819 => x"FF",
		319843 => x"FF",
		320867 => x"FF",
		465251 => x"FF",
		466275 => x"FF",
		467299 => x"FF",
		468323 => x"FF",
		469347 => x"FF",
		19812 => x"FF",
		20836 => x"FF",
		21860 => x"FF",
		22884 => x"FF",
		23908 => x"FF",
		168292 => x"FF",
		169316 => x"FF",
		170340 => x"FF",
		171364 => x"FF",
		172388 => x"FF",
		316772 => x"FF",
		317796 => x"FF",
		318820 => x"FF",
		319844 => x"FF",
		320868 => x"FF",
		465252 => x"FF",
		466276 => x"FF",
		467300 => x"FF",
		468324 => x"FF",
		469348 => x"FF",
		19813 => x"FF",
		20837 => x"FF",
		21861 => x"FF",
		22885 => x"FF",
		23909 => x"FF",
		168293 => x"FF",
		169317 => x"FF",
		170341 => x"FF",
		171365 => x"FF",
		172389 => x"FF",
		316773 => x"FF",
		317797 => x"FF",
		318821 => x"FF",
		319845 => x"FF",
		320869 => x"FF",
		465253 => x"FF",
		466277 => x"FF",
		467301 => x"FF",
		468325 => x"FF",
		469349 => x"FF",
		19814 => x"FF",
		20838 => x"FF",
		21862 => x"FF",
		22886 => x"FF",
		23910 => x"FF",
		168294 => x"FF",
		169318 => x"FF",
		170342 => x"FF",
		171366 => x"FF",
		172390 => x"FF",
		316774 => x"FF",
		317798 => x"FF",
		318822 => x"FF",
		319846 => x"FF",
		320870 => x"FF",
		465254 => x"FF",
		466278 => x"FF",
		467302 => x"FF",
		468326 => x"FF",
		469350 => x"FF",
		19815 => x"FF",
		20839 => x"FF",
		21863 => x"FF",
		22887 => x"FF",
		23911 => x"FF",
		168295 => x"FF",
		169319 => x"FF",
		170343 => x"FF",
		171367 => x"FF",
		172391 => x"FF",
		316775 => x"FF",
		317799 => x"FF",
		318823 => x"FF",
		319847 => x"FF",
		320871 => x"FF",
		465255 => x"FF",
		466279 => x"FF",
		467303 => x"FF",
		468327 => x"FF",
		469351 => x"FF",
		19816 => x"FF",
		20840 => x"FF",
		21864 => x"FF",
		22888 => x"FF",
		23912 => x"FF",
		168296 => x"FF",
		169320 => x"FF",
		170344 => x"FF",
		171368 => x"FF",
		172392 => x"FF",
		316776 => x"FF",
		317800 => x"FF",
		318824 => x"FF",
		319848 => x"FF",
		320872 => x"FF",
		465256 => x"FF",
		466280 => x"FF",
		467304 => x"FF",
		468328 => x"FF",
		469352 => x"FF",
		19817 => x"FF",
		20841 => x"FF",
		21865 => x"FF",
		22889 => x"FF",
		23913 => x"FF",
		168297 => x"FF",
		169321 => x"FF",
		170345 => x"FF",
		171369 => x"FF",
		172393 => x"FF",
		316777 => x"FF",
		317801 => x"FF",
		318825 => x"FF",
		319849 => x"FF",
		320873 => x"FF",
		465257 => x"FF",
		466281 => x"FF",
		467305 => x"FF",
		468329 => x"FF",
		469353 => x"FF",
		19818 => x"FF",
		20842 => x"FF",
		21866 => x"FF",
		22890 => x"FF",
		23914 => x"FF",
		168298 => x"FF",
		169322 => x"FF",
		170346 => x"FF",
		171370 => x"FF",
		172394 => x"FF",
		316778 => x"FF",
		317802 => x"FF",
		318826 => x"FF",
		319850 => x"FF",
		320874 => x"FF",
		465258 => x"FF",
		466282 => x"FF",
		467306 => x"FF",
		468330 => x"FF",
		469354 => x"FF",
		19819 => x"FF",
		20843 => x"FF",
		21867 => x"FF",
		22891 => x"FF",
		23915 => x"FF",
		168299 => x"FF",
		169323 => x"FF",
		170347 => x"FF",
		171371 => x"FF",
		172395 => x"FF",
		316779 => x"FF",
		317803 => x"FF",
		318827 => x"FF",
		319851 => x"FF",
		320875 => x"FF",
		465259 => x"FF",
		466283 => x"FF",
		467307 => x"FF",
		468331 => x"FF",
		469355 => x"FF",
		19820 => x"FF",
		20844 => x"FF",
		21868 => x"FF",
		22892 => x"FF",
		23916 => x"FF",
		168300 => x"FF",
		169324 => x"FF",
		170348 => x"FF",
		171372 => x"FF",
		172396 => x"FF",
		316780 => x"FF",
		317804 => x"FF",
		318828 => x"FF",
		319852 => x"FF",
		320876 => x"FF",
		465260 => x"FF",
		466284 => x"FF",
		467308 => x"FF",
		468332 => x"FF",
		469356 => x"FF",
		19821 => x"FF",
		20845 => x"FF",
		21869 => x"FF",
		22893 => x"FF",
		23917 => x"FF",
		168301 => x"FF",
		169325 => x"FF",
		170349 => x"FF",
		171373 => x"FF",
		172397 => x"FF",
		316781 => x"FF",
		317805 => x"FF",
		318829 => x"FF",
		319853 => x"FF",
		320877 => x"FF",
		465261 => x"FF",
		466285 => x"FF",
		467309 => x"FF",
		468333 => x"FF",
		469357 => x"FF",
		19822 => x"FF",
		20846 => x"FF",
		21870 => x"FF",
		22894 => x"FF",
		23918 => x"FF",
		168302 => x"FF",
		169326 => x"FF",
		170350 => x"FF",
		171374 => x"FF",
		172398 => x"FF",
		316782 => x"FF",
		317806 => x"FF",
		318830 => x"FF",
		319854 => x"FF",
		320878 => x"FF",
		465262 => x"FF",
		466286 => x"FF",
		467310 => x"FF",
		468334 => x"FF",
		469358 => x"FF",
		19823 => x"FF",
		20847 => x"FF",
		21871 => x"FF",
		22895 => x"FF",
		23919 => x"FF",
		168303 => x"FF",
		169327 => x"FF",
		170351 => x"FF",
		171375 => x"FF",
		172399 => x"FF",
		316783 => x"FF",
		317807 => x"FF",
		318831 => x"FF",
		319855 => x"FF",
		320879 => x"FF",
		465263 => x"FF",
		466287 => x"FF",
		467311 => x"FF",
		468335 => x"FF",
		469359 => x"FF",
		19824 => x"FF",
		20848 => x"FF",
		21872 => x"FF",
		22896 => x"FF",
		23920 => x"FF",
		168304 => x"FF",
		169328 => x"FF",
		170352 => x"FF",
		171376 => x"FF",
		172400 => x"FF",
		316784 => x"FF",
		317808 => x"FF",
		318832 => x"FF",
		319856 => x"FF",
		320880 => x"FF",
		465264 => x"FF",
		466288 => x"FF",
		467312 => x"FF",
		468336 => x"FF",
		469360 => x"FF",
		19825 => x"FF",
		20849 => x"FF",
		21873 => x"FF",
		22897 => x"FF",
		23921 => x"FF",
		168305 => x"FF",
		169329 => x"FF",
		170353 => x"FF",
		171377 => x"FF",
		172401 => x"FF",
		316785 => x"FF",
		317809 => x"FF",
		318833 => x"FF",
		319857 => x"FF",
		320881 => x"FF",
		465265 => x"FF",
		466289 => x"FF",
		467313 => x"FF",
		468337 => x"FF",
		469361 => x"FF",
		19826 => x"FF",
		20850 => x"FF",
		21874 => x"FF",
		22898 => x"FF",
		23922 => x"FF",
		168306 => x"FF",
		169330 => x"FF",
		170354 => x"FF",
		171378 => x"FF",
		172402 => x"FF",
		316786 => x"FF",
		317810 => x"FF",
		318834 => x"FF",
		319858 => x"FF",
		320882 => x"FF",
		465266 => x"FF",
		466290 => x"FF",
		467314 => x"FF",
		468338 => x"FF",
		469362 => x"FF",
		19827 => x"FF",
		20851 => x"FF",
		21875 => x"FF",
		22899 => x"FF",
		23923 => x"FF",
		168307 => x"FF",
		169331 => x"FF",
		170355 => x"FF",
		171379 => x"FF",
		172403 => x"FF",
		316787 => x"FF",
		317811 => x"FF",
		318835 => x"FF",
		319859 => x"FF",
		320883 => x"FF",
		465267 => x"FF",
		466291 => x"FF",
		467315 => x"FF",
		468339 => x"FF",
		469363 => x"FF",
		19828 => x"FF",
		20852 => x"FF",
		21876 => x"FF",
		22900 => x"FF",
		23924 => x"FF",
		168308 => x"FF",
		169332 => x"FF",
		170356 => x"FF",
		171380 => x"FF",
		172404 => x"FF",
		316788 => x"FF",
		317812 => x"FF",
		318836 => x"FF",
		319860 => x"FF",
		320884 => x"FF",
		465268 => x"FF",
		466292 => x"FF",
		467316 => x"FF",
		468340 => x"FF",
		469364 => x"FF",
		19829 => x"FF",
		20853 => x"FF",
		21877 => x"FF",
		22901 => x"FF",
		23925 => x"FF",
		168309 => x"FF",
		169333 => x"FF",
		170357 => x"FF",
		171381 => x"FF",
		172405 => x"FF",
		316789 => x"FF",
		317813 => x"FF",
		318837 => x"FF",
		319861 => x"FF",
		320885 => x"FF",
		465269 => x"FF",
		466293 => x"FF",
		467317 => x"FF",
		468341 => x"FF",
		469365 => x"FF",
		19830 => x"FF",
		20854 => x"FF",
		21878 => x"FF",
		22902 => x"FF",
		23926 => x"FF",
		168310 => x"FF",
		169334 => x"FF",
		170358 => x"FF",
		171382 => x"FF",
		172406 => x"FF",
		316790 => x"FF",
		317814 => x"FF",
		318838 => x"FF",
		319862 => x"FF",
		320886 => x"FF",
		465270 => x"FF",
		466294 => x"FF",
		467318 => x"FF",
		468342 => x"FF",
		469366 => x"FF",
		19831 => x"FF",
		20855 => x"FF",
		21879 => x"FF",
		22903 => x"FF",
		23927 => x"FF",
		168311 => x"FF",
		169335 => x"FF",
		170359 => x"FF",
		171383 => x"FF",
		172407 => x"FF",
		316791 => x"FF",
		317815 => x"FF",
		318839 => x"FF",
		319863 => x"FF",
		320887 => x"FF",
		465271 => x"FF",
		466295 => x"FF",
		467319 => x"FF",
		468343 => x"FF",
		469367 => x"FF",
		19832 => x"FF",
		20856 => x"FF",
		21880 => x"FF",
		22904 => x"FF",
		23928 => x"FF",
		168312 => x"FF",
		169336 => x"FF",
		170360 => x"FF",
		171384 => x"FF",
		172408 => x"FF",
		316792 => x"FF",
		317816 => x"FF",
		318840 => x"FF",
		319864 => x"FF",
		320888 => x"FF",
		465272 => x"FF",
		466296 => x"FF",
		467320 => x"FF",
		468344 => x"FF",
		469368 => x"FF",
		19833 => x"FF",
		20857 => x"FF",
		21881 => x"FF",
		22905 => x"FF",
		23929 => x"FF",
		168313 => x"FF",
		169337 => x"FF",
		170361 => x"FF",
		171385 => x"FF",
		172409 => x"FF",
		316793 => x"FF",
		317817 => x"FF",
		318841 => x"FF",
		319865 => x"FF",
		320889 => x"FF",
		465273 => x"FF",
		466297 => x"FF",
		467321 => x"FF",
		468345 => x"FF",
		469369 => x"FF",
		19834 => x"FF",
		20858 => x"FF",
		21882 => x"FF",
		22906 => x"FF",
		23930 => x"FF",
		168314 => x"FF",
		169338 => x"FF",
		170362 => x"FF",
		171386 => x"FF",
		172410 => x"FF",
		316794 => x"FF",
		317818 => x"FF",
		318842 => x"FF",
		319866 => x"FF",
		320890 => x"FF",
		465274 => x"FF",
		466298 => x"FF",
		467322 => x"FF",
		468346 => x"FF",
		469370 => x"FF",
		19835 => x"FF",
		20859 => x"FF",
		21883 => x"FF",
		22907 => x"FF",
		23931 => x"FF",
		168315 => x"FF",
		169339 => x"FF",
		170363 => x"FF",
		171387 => x"FF",
		172411 => x"FF",
		316795 => x"FF",
		317819 => x"FF",
		318843 => x"FF",
		319867 => x"FF",
		320891 => x"FF",
		465275 => x"FF",
		466299 => x"FF",
		467323 => x"FF",
		468347 => x"FF",
		469371 => x"FF",
		19836 => x"FF",
		20860 => x"FF",
		21884 => x"FF",
		22908 => x"FF",
		23932 => x"FF",
		168316 => x"FF",
		169340 => x"FF",
		170364 => x"FF",
		171388 => x"FF",
		172412 => x"FF",
		316796 => x"FF",
		317820 => x"FF",
		318844 => x"FF",
		319868 => x"FF",
		320892 => x"FF",
		465276 => x"FF",
		466300 => x"FF",
		467324 => x"FF",
		468348 => x"FF",
		469372 => x"FF",
		19837 => x"FF",
		20861 => x"FF",
		21885 => x"FF",
		22909 => x"FF",
		23933 => x"FF",
		168317 => x"FF",
		169341 => x"FF",
		170365 => x"FF",
		171389 => x"FF",
		172413 => x"FF",
		316797 => x"FF",
		317821 => x"FF",
		318845 => x"FF",
		319869 => x"FF",
		320893 => x"FF",
		465277 => x"FF",
		466301 => x"FF",
		467325 => x"FF",
		468349 => x"FF",
		469373 => x"FF",
		19838 => x"FF",
		20862 => x"FF",
		21886 => x"FF",
		22910 => x"FF",
		23934 => x"FF",
		168318 => x"FF",
		169342 => x"FF",
		170366 => x"FF",
		171390 => x"FF",
		172414 => x"FF",
		316798 => x"FF",
		317822 => x"FF",
		318846 => x"FF",
		319870 => x"FF",
		320894 => x"FF",
		465278 => x"FF",
		466302 => x"FF",
		467326 => x"FF",
		468350 => x"FF",
		469374 => x"FF",
		19839 => x"FF",
		20863 => x"FF",
		21887 => x"FF",
		22911 => x"FF",
		23935 => x"FF",
		168319 => x"FF",
		169343 => x"FF",
		170367 => x"FF",
		171391 => x"FF",
		172415 => x"FF",
		316799 => x"FF",
		317823 => x"FF",
		318847 => x"FF",
		319871 => x"FF",
		320895 => x"FF",
		465279 => x"FF",
		466303 => x"FF",
		467327 => x"FF",
		468351 => x"FF",
		469375 => x"FF",
		19840 => x"FF",
		20864 => x"FF",
		21888 => x"FF",
		22912 => x"FF",
		23936 => x"FF",
		168320 => x"FF",
		169344 => x"FF",
		170368 => x"FF",
		171392 => x"FF",
		172416 => x"FF",
		316800 => x"FF",
		317824 => x"FF",
		318848 => x"FF",
		319872 => x"FF",
		320896 => x"FF",
		465280 => x"FF",
		466304 => x"FF",
		467328 => x"FF",
		468352 => x"FF",
		469376 => x"FF",
		19841 => x"FF",
		20865 => x"FF",
		21889 => x"FF",
		22913 => x"FF",
		23937 => x"FF",
		168321 => x"FF",
		169345 => x"FF",
		170369 => x"FF",
		171393 => x"FF",
		172417 => x"FF",
		316801 => x"FF",
		317825 => x"FF",
		318849 => x"FF",
		319873 => x"FF",
		320897 => x"FF",
		465281 => x"FF",
		466305 => x"FF",
		467329 => x"FF",
		468353 => x"FF",
		469377 => x"FF",
		19842 => x"FF",
		20866 => x"FF",
		21890 => x"FF",
		22914 => x"FF",
		23938 => x"FF",
		168322 => x"FF",
		169346 => x"FF",
		170370 => x"FF",
		171394 => x"FF",
		172418 => x"FF",
		316802 => x"FF",
		317826 => x"FF",
		318850 => x"FF",
		319874 => x"FF",
		320898 => x"FF",
		465282 => x"FF",
		466306 => x"FF",
		467330 => x"FF",
		468354 => x"FF",
		469378 => x"FF",
		19843 => x"FF",
		20867 => x"FF",
		21891 => x"FF",
		22915 => x"FF",
		23939 => x"FF",
		168323 => x"FF",
		169347 => x"FF",
		170371 => x"FF",
		171395 => x"FF",
		172419 => x"FF",
		316803 => x"FF",
		317827 => x"FF",
		318851 => x"FF",
		319875 => x"FF",
		320899 => x"FF",
		465283 => x"FF",
		466307 => x"FF",
		467331 => x"FF",
		468355 => x"FF",
		469379 => x"FF",
		19844 => x"FF",
		20868 => x"FF",
		21892 => x"FF",
		22916 => x"FF",
		23940 => x"FF",
		168324 => x"FF",
		169348 => x"FF",
		170372 => x"FF",
		171396 => x"FF",
		172420 => x"FF",
		316804 => x"FF",
		317828 => x"FF",
		318852 => x"FF",
		319876 => x"FF",
		320900 => x"FF",
		465284 => x"FF",
		466308 => x"FF",
		467332 => x"FF",
		468356 => x"FF",
		469380 => x"FF",
		19845 => x"FF",
		20869 => x"FF",
		21893 => x"FF",
		22917 => x"FF",
		23941 => x"FF",
		24965 => x"FF",
		25989 => x"FF",
		27013 => x"FF",
		28037 => x"FF",
		29061 => x"FF",
		30085 => x"FF",
		31109 => x"FF",
		32133 => x"FF",
		33157 => x"FF",
		34181 => x"FF",
		35205 => x"FF",
		36229 => x"FF",
		37253 => x"FF",
		38277 => x"FF",
		39301 => x"FF",
		40325 => x"FF",
		41349 => x"FF",
		42373 => x"FF",
		43397 => x"FF",
		44421 => x"FF",
		45445 => x"FF",
		46469 => x"FF",
		47493 => x"FF",
		48517 => x"FF",
		49541 => x"FF",
		50565 => x"FF",
		51589 => x"FF",
		52613 => x"FF",
		53637 => x"FF",
		54661 => x"FF",
		55685 => x"FF",
		56709 => x"FF",
		57733 => x"FF",
		58757 => x"FF",
		59781 => x"FF",
		60805 => x"FF",
		61829 => x"FF",
		62853 => x"FF",
		63877 => x"FF",
		64901 => x"FF",
		65925 => x"FF",
		66949 => x"FF",
		67973 => x"FF",
		68997 => x"FF",
		70021 => x"FF",
		71045 => x"FF",
		72069 => x"FF",
		73093 => x"FF",
		74117 => x"FF",
		75141 => x"FF",
		76165 => x"FF",
		77189 => x"FF",
		78213 => x"FF",
		79237 => x"FF",
		80261 => x"FF",
		81285 => x"FF",
		82309 => x"FF",
		83333 => x"FF",
		84357 => x"FF",
		85381 => x"FF",
		86405 => x"FF",
		87429 => x"FF",
		88453 => x"FF",
		89477 => x"FF",
		90501 => x"FF",
		91525 => x"FF",
		92549 => x"FF",
		93573 => x"FF",
		94597 => x"FF",
		95621 => x"FF",
		96645 => x"FF",
		97669 => x"FF",
		98693 => x"FF",
		99717 => x"FF",
		100741 => x"FF",
		101765 => x"FF",
		102789 => x"FF",
		103813 => x"FF",
		104837 => x"FF",
		105861 => x"FF",
		106885 => x"FF",
		107909 => x"FF",
		108933 => x"FF",
		109957 => x"FF",
		110981 => x"FF",
		112005 => x"FF",
		113029 => x"FF",
		114053 => x"FF",
		115077 => x"FF",
		116101 => x"FF",
		117125 => x"FF",
		118149 => x"FF",
		119173 => x"FF",
		120197 => x"FF",
		121221 => x"FF",
		122245 => x"FF",
		123269 => x"FF",
		124293 => x"FF",
		125317 => x"FF",
		126341 => x"FF",
		127365 => x"FF",
		128389 => x"FF",
		129413 => x"FF",
		130437 => x"FF",
		131461 => x"FF",
		132485 => x"FF",
		133509 => x"FF",
		134533 => x"FF",
		135557 => x"FF",
		136581 => x"FF",
		137605 => x"FF",
		138629 => x"FF",
		139653 => x"FF",
		140677 => x"FF",
		141701 => x"FF",
		142725 => x"FF",
		143749 => x"FF",
		144773 => x"FF",
		145797 => x"FF",
		146821 => x"FF",
		147845 => x"FF",
		148869 => x"FF",
		149893 => x"FF",
		150917 => x"FF",
		151941 => x"FF",
		152965 => x"FF",
		153989 => x"FF",
		155013 => x"FF",
		156037 => x"FF",
		157061 => x"FF",
		158085 => x"FF",
		159109 => x"FF",
		160133 => x"FF",
		161157 => x"FF",
		162181 => x"FF",
		163205 => x"FF",
		164229 => x"FF",
		165253 => x"FF",
		166277 => x"FF",
		167301 => x"FF",
		168325 => x"FF",
		169349 => x"FF",
		170373 => x"FF",
		171397 => x"FF",
		172421 => x"FF",
		173445 => x"FF",
		174469 => x"FF",
		175493 => x"FF",
		176517 => x"FF",
		177541 => x"FF",
		178565 => x"FF",
		179589 => x"FF",
		180613 => x"FF",
		181637 => x"FF",
		182661 => x"FF",
		183685 => x"FF",
		184709 => x"FF",
		185733 => x"FF",
		186757 => x"FF",
		187781 => x"FF",
		188805 => x"FF",
		189829 => x"FF",
		190853 => x"FF",
		191877 => x"FF",
		192901 => x"FF",
		193925 => x"FF",
		194949 => x"FF",
		195973 => x"FF",
		196997 => x"FF",
		198021 => x"FF",
		199045 => x"FF",
		200069 => x"FF",
		201093 => x"FF",
		202117 => x"FF",
		203141 => x"FF",
		204165 => x"FF",
		205189 => x"FF",
		206213 => x"FF",
		207237 => x"FF",
		208261 => x"FF",
		209285 => x"FF",
		210309 => x"FF",
		211333 => x"FF",
		212357 => x"FF",
		213381 => x"FF",
		214405 => x"FF",
		215429 => x"FF",
		216453 => x"FF",
		217477 => x"FF",
		218501 => x"FF",
		219525 => x"FF",
		220549 => x"FF",
		221573 => x"FF",
		222597 => x"FF",
		223621 => x"FF",
		224645 => x"FF",
		225669 => x"FF",
		226693 => x"FF",
		227717 => x"FF",
		228741 => x"FF",
		229765 => x"FF",
		230789 => x"FF",
		231813 => x"FF",
		232837 => x"FF",
		233861 => x"FF",
		234885 => x"FF",
		235909 => x"FF",
		236933 => x"FF",
		237957 => x"FF",
		238981 => x"FF",
		240005 => x"FF",
		241029 => x"FF",
		242053 => x"FF",
		243077 => x"FF",
		244101 => x"FF",
		245125 => x"FF",
		246149 => x"FF",
		247173 => x"FF",
		248197 => x"FF",
		249221 => x"FF",
		250245 => x"FF",
		251269 => x"FF",
		252293 => x"FF",
		253317 => x"FF",
		254341 => x"FF",
		255365 => x"FF",
		256389 => x"FF",
		257413 => x"FF",
		258437 => x"FF",
		259461 => x"FF",
		260485 => x"FF",
		261509 => x"FF",
		262533 => x"FF",
		263557 => x"FF",
		264581 => x"FF",
		265605 => x"FF",
		266629 => x"FF",
		267653 => x"FF",
		268677 => x"FF",
		269701 => x"FF",
		270725 => x"FF",
		271749 => x"FF",
		272773 => x"FF",
		273797 => x"FF",
		274821 => x"FF",
		275845 => x"FF",
		276869 => x"FF",
		277893 => x"FF",
		278917 => x"FF",
		279941 => x"FF",
		280965 => x"FF",
		281989 => x"FF",
		283013 => x"FF",
		284037 => x"FF",
		285061 => x"FF",
		286085 => x"FF",
		287109 => x"FF",
		288133 => x"FF",
		289157 => x"FF",
		290181 => x"FF",
		291205 => x"FF",
		292229 => x"FF",
		293253 => x"FF",
		294277 => x"FF",
		295301 => x"FF",
		296325 => x"FF",
		297349 => x"FF",
		298373 => x"FF",
		299397 => x"FF",
		300421 => x"FF",
		301445 => x"FF",
		302469 => x"FF",
		303493 => x"FF",
		304517 => x"FF",
		305541 => x"FF",
		306565 => x"FF",
		307589 => x"FF",
		308613 => x"FF",
		309637 => x"FF",
		310661 => x"FF",
		311685 => x"FF",
		312709 => x"FF",
		313733 => x"FF",
		314757 => x"FF",
		315781 => x"FF",
		316805 => x"FF",
		317829 => x"FF",
		318853 => x"FF",
		319877 => x"FF",
		320901 => x"FF",
		321925 => x"FF",
		322949 => x"FF",
		323973 => x"FF",
		324997 => x"FF",
		326021 => x"FF",
		327045 => x"FF",
		328069 => x"FF",
		329093 => x"FF",
		330117 => x"FF",
		331141 => x"FF",
		332165 => x"FF",
		333189 => x"FF",
		334213 => x"FF",
		335237 => x"FF",
		336261 => x"FF",
		337285 => x"FF",
		338309 => x"FF",
		339333 => x"FF",
		340357 => x"FF",
		341381 => x"FF",
		342405 => x"FF",
		343429 => x"FF",
		344453 => x"FF",
		345477 => x"FF",
		346501 => x"FF",
		347525 => x"FF",
		348549 => x"FF",
		349573 => x"FF",
		350597 => x"FF",
		351621 => x"FF",
		352645 => x"FF",
		353669 => x"FF",
		354693 => x"FF",
		355717 => x"FF",
		356741 => x"FF",
		357765 => x"FF",
		358789 => x"FF",
		359813 => x"FF",
		360837 => x"FF",
		361861 => x"FF",
		362885 => x"FF",
		363909 => x"FF",
		364933 => x"FF",
		365957 => x"FF",
		366981 => x"FF",
		368005 => x"FF",
		369029 => x"FF",
		370053 => x"FF",
		371077 => x"FF",
		372101 => x"FF",
		373125 => x"FF",
		374149 => x"FF",
		375173 => x"FF",
		376197 => x"FF",
		377221 => x"FF",
		378245 => x"FF",
		379269 => x"FF",
		380293 => x"FF",
		381317 => x"FF",
		382341 => x"FF",
		383365 => x"FF",
		384389 => x"FF",
		385413 => x"FF",
		386437 => x"FF",
		387461 => x"FF",
		388485 => x"FF",
		389509 => x"FF",
		390533 => x"FF",
		391557 => x"FF",
		392581 => x"FF",
		393605 => x"FF",
		394629 => x"FF",
		395653 => x"FF",
		396677 => x"FF",
		397701 => x"FF",
		398725 => x"FF",
		399749 => x"FF",
		400773 => x"FF",
		401797 => x"FF",
		402821 => x"FF",
		403845 => x"FF",
		404869 => x"FF",
		405893 => x"FF",
		406917 => x"FF",
		407941 => x"FF",
		408965 => x"FF",
		409989 => x"FF",
		411013 => x"FF",
		412037 => x"FF",
		413061 => x"FF",
		414085 => x"FF",
		415109 => x"FF",
		416133 => x"FF",
		417157 => x"FF",
		418181 => x"FF",
		419205 => x"FF",
		420229 => x"FF",
		421253 => x"FF",
		422277 => x"FF",
		423301 => x"FF",
		424325 => x"FF",
		425349 => x"FF",
		426373 => x"FF",
		427397 => x"FF",
		428421 => x"FF",
		429445 => x"FF",
		430469 => x"FF",
		431493 => x"FF",
		432517 => x"FF",
		433541 => x"FF",
		434565 => x"FF",
		435589 => x"FF",
		436613 => x"FF",
		437637 => x"FF",
		438661 => x"FF",
		439685 => x"FF",
		440709 => x"FF",
		441733 => x"FF",
		442757 => x"FF",
		443781 => x"FF",
		444805 => x"FF",
		445829 => x"FF",
		446853 => x"FF",
		447877 => x"FF",
		448901 => x"FF",
		449925 => x"FF",
		450949 => x"FF",
		451973 => x"FF",
		452997 => x"FF",
		454021 => x"FF",
		455045 => x"FF",
		456069 => x"FF",
		457093 => x"FF",
		458117 => x"FF",
		459141 => x"FF",
		460165 => x"FF",
		461189 => x"FF",
		462213 => x"FF",
		463237 => x"FF",
		464261 => x"FF",
		465285 => x"FF",
		466309 => x"FF",
		467333 => x"FF",
		468357 => x"FF",
		469381 => x"FF",
		19846 => x"FF",
		20870 => x"FF",
		21894 => x"FF",
		22918 => x"FF",
		23942 => x"FF",
		24966 => x"FF",
		25990 => x"FF",
		27014 => x"FF",
		28038 => x"FF",
		29062 => x"FF",
		30086 => x"FF",
		31110 => x"FF",
		32134 => x"FF",
		33158 => x"FF",
		34182 => x"FF",
		35206 => x"FF",
		36230 => x"FF",
		37254 => x"FF",
		38278 => x"FF",
		39302 => x"FF",
		40326 => x"FF",
		41350 => x"FF",
		42374 => x"FF",
		43398 => x"FF",
		44422 => x"FF",
		45446 => x"FF",
		46470 => x"FF",
		47494 => x"FF",
		48518 => x"FF",
		49542 => x"FF",
		50566 => x"FF",
		51590 => x"FF",
		52614 => x"FF",
		53638 => x"FF",
		54662 => x"FF",
		55686 => x"FF",
		56710 => x"FF",
		57734 => x"FF",
		58758 => x"FF",
		59782 => x"FF",
		60806 => x"FF",
		61830 => x"FF",
		62854 => x"FF",
		63878 => x"FF",
		64902 => x"FF",
		65926 => x"FF",
		66950 => x"FF",
		67974 => x"FF",
		68998 => x"FF",
		70022 => x"FF",
		71046 => x"FF",
		72070 => x"FF",
		73094 => x"FF",
		74118 => x"FF",
		75142 => x"FF",
		76166 => x"FF",
		77190 => x"FF",
		78214 => x"FF",
		79238 => x"FF",
		80262 => x"FF",
		81286 => x"FF",
		82310 => x"FF",
		83334 => x"FF",
		84358 => x"FF",
		85382 => x"FF",
		86406 => x"FF",
		87430 => x"FF",
		88454 => x"FF",
		89478 => x"FF",
		90502 => x"FF",
		91526 => x"FF",
		92550 => x"FF",
		93574 => x"FF",
		94598 => x"FF",
		95622 => x"FF",
		96646 => x"FF",
		97670 => x"FF",
		98694 => x"FF",
		99718 => x"FF",
		100742 => x"FF",
		101766 => x"FF",
		102790 => x"FF",
		103814 => x"FF",
		104838 => x"FF",
		105862 => x"FF",
		106886 => x"FF",
		107910 => x"FF",
		108934 => x"FF",
		109958 => x"FF",
		110982 => x"FF",
		112006 => x"FF",
		113030 => x"FF",
		114054 => x"FF",
		115078 => x"FF",
		116102 => x"FF",
		117126 => x"FF",
		118150 => x"FF",
		119174 => x"FF",
		120198 => x"FF",
		121222 => x"FF",
		122246 => x"FF",
		123270 => x"FF",
		124294 => x"FF",
		125318 => x"FF",
		126342 => x"FF",
		127366 => x"FF",
		128390 => x"FF",
		129414 => x"FF",
		130438 => x"FF",
		131462 => x"FF",
		132486 => x"FF",
		133510 => x"FF",
		134534 => x"FF",
		135558 => x"FF",
		136582 => x"FF",
		137606 => x"FF",
		138630 => x"FF",
		139654 => x"FF",
		140678 => x"FF",
		141702 => x"FF",
		142726 => x"FF",
		143750 => x"FF",
		144774 => x"FF",
		145798 => x"FF",
		146822 => x"FF",
		147846 => x"FF",
		148870 => x"FF",
		149894 => x"FF",
		150918 => x"FF",
		151942 => x"FF",
		152966 => x"FF",
		153990 => x"FF",
		155014 => x"FF",
		156038 => x"FF",
		157062 => x"FF",
		158086 => x"FF",
		159110 => x"FF",
		160134 => x"FF",
		161158 => x"FF",
		162182 => x"FF",
		163206 => x"FF",
		164230 => x"FF",
		165254 => x"FF",
		166278 => x"FF",
		167302 => x"FF",
		168326 => x"FF",
		169350 => x"FF",
		170374 => x"FF",
		171398 => x"FF",
		172422 => x"FF",
		173446 => x"FF",
		174470 => x"FF",
		175494 => x"FF",
		176518 => x"FF",
		177542 => x"FF",
		178566 => x"FF",
		179590 => x"FF",
		180614 => x"FF",
		181638 => x"FF",
		182662 => x"FF",
		183686 => x"FF",
		184710 => x"FF",
		185734 => x"FF",
		186758 => x"FF",
		187782 => x"FF",
		188806 => x"FF",
		189830 => x"FF",
		190854 => x"FF",
		191878 => x"FF",
		192902 => x"FF",
		193926 => x"FF",
		194950 => x"FF",
		195974 => x"FF",
		196998 => x"FF",
		198022 => x"FF",
		199046 => x"FF",
		200070 => x"FF",
		201094 => x"FF",
		202118 => x"FF",
		203142 => x"FF",
		204166 => x"FF",
		205190 => x"FF",
		206214 => x"FF",
		207238 => x"FF",
		208262 => x"FF",
		209286 => x"FF",
		210310 => x"FF",
		211334 => x"FF",
		212358 => x"FF",
		213382 => x"FF",
		214406 => x"FF",
		215430 => x"FF",
		216454 => x"FF",
		217478 => x"FF",
		218502 => x"FF",
		219526 => x"FF",
		220550 => x"FF",
		221574 => x"FF",
		222598 => x"FF",
		223622 => x"FF",
		224646 => x"FF",
		225670 => x"FF",
		226694 => x"FF",
		227718 => x"FF",
		228742 => x"FF",
		229766 => x"FF",
		230790 => x"FF",
		231814 => x"FF",
		232838 => x"FF",
		233862 => x"FF",
		234886 => x"FF",
		235910 => x"FF",
		236934 => x"FF",
		237958 => x"FF",
		238982 => x"FF",
		240006 => x"FF",
		241030 => x"FF",
		242054 => x"FF",
		243078 => x"FF",
		244102 => x"FF",
		245126 => x"FF",
		246150 => x"FF",
		247174 => x"FF",
		248198 => x"FF",
		249222 => x"FF",
		250246 => x"FF",
		251270 => x"FF",
		252294 => x"FF",
		253318 => x"FF",
		254342 => x"FF",
		255366 => x"FF",
		256390 => x"FF",
		257414 => x"FF",
		258438 => x"FF",
		259462 => x"FF",
		260486 => x"FF",
		261510 => x"FF",
		262534 => x"FF",
		263558 => x"FF",
		264582 => x"FF",
		265606 => x"FF",
		266630 => x"FF",
		267654 => x"FF",
		268678 => x"FF",
		269702 => x"FF",
		270726 => x"FF",
		271750 => x"FF",
		272774 => x"FF",
		273798 => x"FF",
		274822 => x"FF",
		275846 => x"FF",
		276870 => x"FF",
		277894 => x"FF",
		278918 => x"FF",
		279942 => x"FF",
		280966 => x"FF",
		281990 => x"FF",
		283014 => x"FF",
		284038 => x"FF",
		285062 => x"FF",
		286086 => x"FF",
		287110 => x"FF",
		288134 => x"FF",
		289158 => x"FF",
		290182 => x"FF",
		291206 => x"FF",
		292230 => x"FF",
		293254 => x"FF",
		294278 => x"FF",
		295302 => x"FF",
		296326 => x"FF",
		297350 => x"FF",
		298374 => x"FF",
		299398 => x"FF",
		300422 => x"FF",
		301446 => x"FF",
		302470 => x"FF",
		303494 => x"FF",
		304518 => x"FF",
		305542 => x"FF",
		306566 => x"FF",
		307590 => x"FF",
		308614 => x"FF",
		309638 => x"FF",
		310662 => x"FF",
		311686 => x"FF",
		312710 => x"FF",
		313734 => x"FF",
		314758 => x"FF",
		315782 => x"FF",
		316806 => x"FF",
		317830 => x"FF",
		318854 => x"FF",
		319878 => x"FF",
		320902 => x"FF",
		321926 => x"FF",
		322950 => x"FF",
		323974 => x"FF",
		324998 => x"FF",
		326022 => x"FF",
		327046 => x"FF",
		328070 => x"FF",
		329094 => x"FF",
		330118 => x"FF",
		331142 => x"FF",
		332166 => x"FF",
		333190 => x"FF",
		334214 => x"FF",
		335238 => x"FF",
		336262 => x"FF",
		337286 => x"FF",
		338310 => x"FF",
		339334 => x"FF",
		340358 => x"FF",
		341382 => x"FF",
		342406 => x"FF",
		343430 => x"FF",
		344454 => x"FF",
		345478 => x"FF",
		346502 => x"FF",
		347526 => x"FF",
		348550 => x"FF",
		349574 => x"FF",
		350598 => x"FF",
		351622 => x"FF",
		352646 => x"FF",
		353670 => x"FF",
		354694 => x"FF",
		355718 => x"FF",
		356742 => x"FF",
		357766 => x"FF",
		358790 => x"FF",
		359814 => x"FF",
		360838 => x"FF",
		361862 => x"FF",
		362886 => x"FF",
		363910 => x"FF",
		364934 => x"FF",
		365958 => x"FF",
		366982 => x"FF",
		368006 => x"FF",
		369030 => x"FF",
		370054 => x"FF",
		371078 => x"FF",
		372102 => x"FF",
		373126 => x"FF",
		374150 => x"FF",
		375174 => x"FF",
		376198 => x"FF",
		377222 => x"FF",
		378246 => x"FF",
		379270 => x"FF",
		380294 => x"FF",
		381318 => x"FF",
		382342 => x"FF",
		383366 => x"FF",
		384390 => x"FF",
		385414 => x"FF",
		386438 => x"FF",
		387462 => x"FF",
		388486 => x"FF",
		389510 => x"FF",
		390534 => x"FF",
		391558 => x"FF",
		392582 => x"FF",
		393606 => x"FF",
		394630 => x"FF",
		395654 => x"FF",
		396678 => x"FF",
		397702 => x"FF",
		398726 => x"FF",
		399750 => x"FF",
		400774 => x"FF",
		401798 => x"FF",
		402822 => x"FF",
		403846 => x"FF",
		404870 => x"FF",
		405894 => x"FF",
		406918 => x"FF",
		407942 => x"FF",
		408966 => x"FF",
		409990 => x"FF",
		411014 => x"FF",
		412038 => x"FF",
		413062 => x"FF",
		414086 => x"FF",
		415110 => x"FF",
		416134 => x"FF",
		417158 => x"FF",
		418182 => x"FF",
		419206 => x"FF",
		420230 => x"FF",
		421254 => x"FF",
		422278 => x"FF",
		423302 => x"FF",
		424326 => x"FF",
		425350 => x"FF",
		426374 => x"FF",
		427398 => x"FF",
		428422 => x"FF",
		429446 => x"FF",
		430470 => x"FF",
		431494 => x"FF",
		432518 => x"FF",
		433542 => x"FF",
		434566 => x"FF",
		435590 => x"FF",
		436614 => x"FF",
		437638 => x"FF",
		438662 => x"FF",
		439686 => x"FF",
		440710 => x"FF",
		441734 => x"FF",
		442758 => x"FF",
		443782 => x"FF",
		444806 => x"FF",
		445830 => x"FF",
		446854 => x"FF",
		447878 => x"FF",
		448902 => x"FF",
		449926 => x"FF",
		450950 => x"FF",
		451974 => x"FF",
		452998 => x"FF",
		454022 => x"FF",
		455046 => x"FF",
		456070 => x"FF",
		457094 => x"FF",
		458118 => x"FF",
		459142 => x"FF",
		460166 => x"FF",
		461190 => x"FF",
		462214 => x"FF",
		463238 => x"FF",
		464262 => x"FF",
		465286 => x"FF",
		466310 => x"FF",
		467334 => x"FF",
		468358 => x"FF",
		469382 => x"FF",
		19847 => x"FF",
		20871 => x"FF",
		21895 => x"FF",
		22919 => x"FF",
		23943 => x"FF",
		24967 => x"FF",
		25991 => x"FF",
		27015 => x"FF",
		28039 => x"FF",
		29063 => x"FF",
		30087 => x"FF",
		31111 => x"FF",
		32135 => x"FF",
		33159 => x"FF",
		34183 => x"FF",
		35207 => x"FF",
		36231 => x"FF",
		37255 => x"FF",
		38279 => x"FF",
		39303 => x"FF",
		40327 => x"FF",
		41351 => x"FF",
		42375 => x"FF",
		43399 => x"FF",
		44423 => x"FF",
		45447 => x"FF",
		46471 => x"FF",
		47495 => x"FF",
		48519 => x"FF",
		49543 => x"FF",
		50567 => x"FF",
		51591 => x"FF",
		52615 => x"FF",
		53639 => x"FF",
		54663 => x"FF",
		55687 => x"FF",
		56711 => x"FF",
		57735 => x"FF",
		58759 => x"FF",
		59783 => x"FF",
		60807 => x"FF",
		61831 => x"FF",
		62855 => x"FF",
		63879 => x"FF",
		64903 => x"FF",
		65927 => x"FF",
		66951 => x"FF",
		67975 => x"FF",
		68999 => x"FF",
		70023 => x"FF",
		71047 => x"FF",
		72071 => x"FF",
		73095 => x"FF",
		74119 => x"FF",
		75143 => x"FF",
		76167 => x"FF",
		77191 => x"FF",
		78215 => x"FF",
		79239 => x"FF",
		80263 => x"FF",
		81287 => x"FF",
		82311 => x"FF",
		83335 => x"FF",
		84359 => x"FF",
		85383 => x"FF",
		86407 => x"FF",
		87431 => x"FF",
		88455 => x"FF",
		89479 => x"FF",
		90503 => x"FF",
		91527 => x"FF",
		92551 => x"FF",
		93575 => x"FF",
		94599 => x"FF",
		95623 => x"FF",
		96647 => x"FF",
		97671 => x"FF",
		98695 => x"FF",
		99719 => x"FF",
		100743 => x"FF",
		101767 => x"FF",
		102791 => x"FF",
		103815 => x"FF",
		104839 => x"FF",
		105863 => x"FF",
		106887 => x"FF",
		107911 => x"FF",
		108935 => x"FF",
		109959 => x"FF",
		110983 => x"FF",
		112007 => x"FF",
		113031 => x"FF",
		114055 => x"FF",
		115079 => x"FF",
		116103 => x"FF",
		117127 => x"FF",
		118151 => x"FF",
		119175 => x"FF",
		120199 => x"FF",
		121223 => x"FF",
		122247 => x"FF",
		123271 => x"FF",
		124295 => x"FF",
		125319 => x"FF",
		126343 => x"FF",
		127367 => x"FF",
		128391 => x"FF",
		129415 => x"FF",
		130439 => x"FF",
		131463 => x"FF",
		132487 => x"FF",
		133511 => x"FF",
		134535 => x"FF",
		135559 => x"FF",
		136583 => x"FF",
		137607 => x"FF",
		138631 => x"FF",
		139655 => x"FF",
		140679 => x"FF",
		141703 => x"FF",
		142727 => x"FF",
		143751 => x"FF",
		144775 => x"FF",
		145799 => x"FF",
		146823 => x"FF",
		147847 => x"FF",
		148871 => x"FF",
		149895 => x"FF",
		150919 => x"FF",
		151943 => x"FF",
		152967 => x"FF",
		153991 => x"FF",
		155015 => x"FF",
		156039 => x"FF",
		157063 => x"FF",
		158087 => x"FF",
		159111 => x"FF",
		160135 => x"FF",
		161159 => x"FF",
		162183 => x"FF",
		163207 => x"FF",
		164231 => x"FF",
		165255 => x"FF",
		166279 => x"FF",
		167303 => x"FF",
		168327 => x"FF",
		169351 => x"FF",
		170375 => x"FF",
		171399 => x"FF",
		172423 => x"FF",
		173447 => x"FF",
		174471 => x"FF",
		175495 => x"FF",
		176519 => x"FF",
		177543 => x"FF",
		178567 => x"FF",
		179591 => x"FF",
		180615 => x"FF",
		181639 => x"FF",
		182663 => x"FF",
		183687 => x"FF",
		184711 => x"FF",
		185735 => x"FF",
		186759 => x"FF",
		187783 => x"FF",
		188807 => x"FF",
		189831 => x"FF",
		190855 => x"FF",
		191879 => x"FF",
		192903 => x"FF",
		193927 => x"FF",
		194951 => x"FF",
		195975 => x"FF",
		196999 => x"FF",
		198023 => x"FF",
		199047 => x"FF",
		200071 => x"FF",
		201095 => x"FF",
		202119 => x"FF",
		203143 => x"FF",
		204167 => x"FF",
		205191 => x"FF",
		206215 => x"FF",
		207239 => x"FF",
		208263 => x"FF",
		209287 => x"FF",
		210311 => x"FF",
		211335 => x"FF",
		212359 => x"FF",
		213383 => x"FF",
		214407 => x"FF",
		215431 => x"FF",
		216455 => x"FF",
		217479 => x"FF",
		218503 => x"FF",
		219527 => x"FF",
		220551 => x"FF",
		221575 => x"FF",
		222599 => x"FF",
		223623 => x"FF",
		224647 => x"FF",
		225671 => x"FF",
		226695 => x"FF",
		227719 => x"FF",
		228743 => x"FF",
		229767 => x"FF",
		230791 => x"FF",
		231815 => x"FF",
		232839 => x"FF",
		233863 => x"FF",
		234887 => x"FF",
		235911 => x"FF",
		236935 => x"FF",
		237959 => x"FF",
		238983 => x"FF",
		240007 => x"FF",
		241031 => x"FF",
		242055 => x"FF",
		243079 => x"FF",
		244103 => x"FF",
		245127 => x"FF",
		246151 => x"FF",
		247175 => x"FF",
		248199 => x"FF",
		249223 => x"FF",
		250247 => x"FF",
		251271 => x"FF",
		252295 => x"FF",
		253319 => x"FF",
		254343 => x"FF",
		255367 => x"FF",
		256391 => x"FF",
		257415 => x"FF",
		258439 => x"FF",
		259463 => x"FF",
		260487 => x"FF",
		261511 => x"FF",
		262535 => x"FF",
		263559 => x"FF",
		264583 => x"FF",
		265607 => x"FF",
		266631 => x"FF",
		267655 => x"FF",
		268679 => x"FF",
		269703 => x"FF",
		270727 => x"FF",
		271751 => x"FF",
		272775 => x"FF",
		273799 => x"FF",
		274823 => x"FF",
		275847 => x"FF",
		276871 => x"FF",
		277895 => x"FF",
		278919 => x"FF",
		279943 => x"FF",
		280967 => x"FF",
		281991 => x"FF",
		283015 => x"FF",
		284039 => x"FF",
		285063 => x"FF",
		286087 => x"FF",
		287111 => x"FF",
		288135 => x"FF",
		289159 => x"FF",
		290183 => x"FF",
		291207 => x"FF",
		292231 => x"FF",
		293255 => x"FF",
		294279 => x"FF",
		295303 => x"FF",
		296327 => x"FF",
		297351 => x"FF",
		298375 => x"FF",
		299399 => x"FF",
		300423 => x"FF",
		301447 => x"FF",
		302471 => x"FF",
		303495 => x"FF",
		304519 => x"FF",
		305543 => x"FF",
		306567 => x"FF",
		307591 => x"FF",
		308615 => x"FF",
		309639 => x"FF",
		310663 => x"FF",
		311687 => x"FF",
		312711 => x"FF",
		313735 => x"FF",
		314759 => x"FF",
		315783 => x"FF",
		316807 => x"FF",
		317831 => x"FF",
		318855 => x"FF",
		319879 => x"FF",
		320903 => x"FF",
		321927 => x"FF",
		322951 => x"FF",
		323975 => x"FF",
		324999 => x"FF",
		326023 => x"FF",
		327047 => x"FF",
		328071 => x"FF",
		329095 => x"FF",
		330119 => x"FF",
		331143 => x"FF",
		332167 => x"FF",
		333191 => x"FF",
		334215 => x"FF",
		335239 => x"FF",
		336263 => x"FF",
		337287 => x"FF",
		338311 => x"FF",
		339335 => x"FF",
		340359 => x"FF",
		341383 => x"FF",
		342407 => x"FF",
		343431 => x"FF",
		344455 => x"FF",
		345479 => x"FF",
		346503 => x"FF",
		347527 => x"FF",
		348551 => x"FF",
		349575 => x"FF",
		350599 => x"FF",
		351623 => x"FF",
		352647 => x"FF",
		353671 => x"FF",
		354695 => x"FF",
		355719 => x"FF",
		356743 => x"FF",
		357767 => x"FF",
		358791 => x"FF",
		359815 => x"FF",
		360839 => x"FF",
		361863 => x"FF",
		362887 => x"FF",
		363911 => x"FF",
		364935 => x"FF",
		365959 => x"FF",
		366983 => x"FF",
		368007 => x"FF",
		369031 => x"FF",
		370055 => x"FF",
		371079 => x"FF",
		372103 => x"FF",
		373127 => x"FF",
		374151 => x"FF",
		375175 => x"FF",
		376199 => x"FF",
		377223 => x"FF",
		378247 => x"FF",
		379271 => x"FF",
		380295 => x"FF",
		381319 => x"FF",
		382343 => x"FF",
		383367 => x"FF",
		384391 => x"FF",
		385415 => x"FF",
		386439 => x"FF",
		387463 => x"FF",
		388487 => x"FF",
		389511 => x"FF",
		390535 => x"FF",
		391559 => x"FF",
		392583 => x"FF",
		393607 => x"FF",
		394631 => x"FF",
		395655 => x"FF",
		396679 => x"FF",
		397703 => x"FF",
		398727 => x"FF",
		399751 => x"FF",
		400775 => x"FF",
		401799 => x"FF",
		402823 => x"FF",
		403847 => x"FF",
		404871 => x"FF",
		405895 => x"FF",
		406919 => x"FF",
		407943 => x"FF",
		408967 => x"FF",
		409991 => x"FF",
		411015 => x"FF",
		412039 => x"FF",
		413063 => x"FF",
		414087 => x"FF",
		415111 => x"FF",
		416135 => x"FF",
		417159 => x"FF",
		418183 => x"FF",
		419207 => x"FF",
		420231 => x"FF",
		421255 => x"FF",
		422279 => x"FF",
		423303 => x"FF",
		424327 => x"FF",
		425351 => x"FF",
		426375 => x"FF",
		427399 => x"FF",
		428423 => x"FF",
		429447 => x"FF",
		430471 => x"FF",
		431495 => x"FF",
		432519 => x"FF",
		433543 => x"FF",
		434567 => x"FF",
		435591 => x"FF",
		436615 => x"FF",
		437639 => x"FF",
		438663 => x"FF",
		439687 => x"FF",
		440711 => x"FF",
		441735 => x"FF",
		442759 => x"FF",
		443783 => x"FF",
		444807 => x"FF",
		445831 => x"FF",
		446855 => x"FF",
		447879 => x"FF",
		448903 => x"FF",
		449927 => x"FF",
		450951 => x"FF",
		451975 => x"FF",
		452999 => x"FF",
		454023 => x"FF",
		455047 => x"FF",
		456071 => x"FF",
		457095 => x"FF",
		458119 => x"FF",
		459143 => x"FF",
		460167 => x"FF",
		461191 => x"FF",
		462215 => x"FF",
		463239 => x"FF",
		464263 => x"FF",
		465287 => x"FF",
		466311 => x"FF",
		467335 => x"FF",
		468359 => x"FF",
		469383 => x"FF",
		19848 => x"FF",
		20872 => x"FF",
		21896 => x"FF",
		22920 => x"FF",
		23944 => x"FF",
		24968 => x"FF",
		25992 => x"FF",
		27016 => x"FF",
		28040 => x"FF",
		29064 => x"FF",
		30088 => x"FF",
		31112 => x"FF",
		32136 => x"FF",
		33160 => x"FF",
		34184 => x"FF",
		35208 => x"FF",
		36232 => x"FF",
		37256 => x"FF",
		38280 => x"FF",
		39304 => x"FF",
		40328 => x"FF",
		41352 => x"FF",
		42376 => x"FF",
		43400 => x"FF",
		44424 => x"FF",
		45448 => x"FF",
		46472 => x"FF",
		47496 => x"FF",
		48520 => x"FF",
		49544 => x"FF",
		50568 => x"FF",
		51592 => x"FF",
		52616 => x"FF",
		53640 => x"FF",
		54664 => x"FF",
		55688 => x"FF",
		56712 => x"FF",
		57736 => x"FF",
		58760 => x"FF",
		59784 => x"FF",
		60808 => x"FF",
		61832 => x"FF",
		62856 => x"FF",
		63880 => x"FF",
		64904 => x"FF",
		65928 => x"FF",
		66952 => x"FF",
		67976 => x"FF",
		69000 => x"FF",
		70024 => x"FF",
		71048 => x"FF",
		72072 => x"FF",
		73096 => x"FF",
		74120 => x"FF",
		75144 => x"FF",
		76168 => x"FF",
		77192 => x"FF",
		78216 => x"FF",
		79240 => x"FF",
		80264 => x"FF",
		81288 => x"FF",
		82312 => x"FF",
		83336 => x"FF",
		84360 => x"FF",
		85384 => x"FF",
		86408 => x"FF",
		87432 => x"FF",
		88456 => x"FF",
		89480 => x"FF",
		90504 => x"FF",
		91528 => x"FF",
		92552 => x"FF",
		93576 => x"FF",
		94600 => x"FF",
		95624 => x"FF",
		96648 => x"FF",
		97672 => x"FF",
		98696 => x"FF",
		99720 => x"FF",
		100744 => x"FF",
		101768 => x"FF",
		102792 => x"FF",
		103816 => x"FF",
		104840 => x"FF",
		105864 => x"FF",
		106888 => x"FF",
		107912 => x"FF",
		108936 => x"FF",
		109960 => x"FF",
		110984 => x"FF",
		112008 => x"FF",
		113032 => x"FF",
		114056 => x"FF",
		115080 => x"FF",
		116104 => x"FF",
		117128 => x"FF",
		118152 => x"FF",
		119176 => x"FF",
		120200 => x"FF",
		121224 => x"FF",
		122248 => x"FF",
		123272 => x"FF",
		124296 => x"FF",
		125320 => x"FF",
		126344 => x"FF",
		127368 => x"FF",
		128392 => x"FF",
		129416 => x"FF",
		130440 => x"FF",
		131464 => x"FF",
		132488 => x"FF",
		133512 => x"FF",
		134536 => x"FF",
		135560 => x"FF",
		136584 => x"FF",
		137608 => x"FF",
		138632 => x"FF",
		139656 => x"FF",
		140680 => x"FF",
		141704 => x"FF",
		142728 => x"FF",
		143752 => x"FF",
		144776 => x"FF",
		145800 => x"FF",
		146824 => x"FF",
		147848 => x"FF",
		148872 => x"FF",
		149896 => x"FF",
		150920 => x"FF",
		151944 => x"FF",
		152968 => x"FF",
		153992 => x"FF",
		155016 => x"FF",
		156040 => x"FF",
		157064 => x"FF",
		158088 => x"FF",
		159112 => x"FF",
		160136 => x"FF",
		161160 => x"FF",
		162184 => x"FF",
		163208 => x"FF",
		164232 => x"FF",
		165256 => x"FF",
		166280 => x"FF",
		167304 => x"FF",
		168328 => x"FF",
		169352 => x"FF",
		170376 => x"FF",
		171400 => x"FF",
		172424 => x"FF",
		173448 => x"FF",
		174472 => x"FF",
		175496 => x"FF",
		176520 => x"FF",
		177544 => x"FF",
		178568 => x"FF",
		179592 => x"FF",
		180616 => x"FF",
		181640 => x"FF",
		182664 => x"FF",
		183688 => x"FF",
		184712 => x"FF",
		185736 => x"FF",
		186760 => x"FF",
		187784 => x"FF",
		188808 => x"FF",
		189832 => x"FF",
		190856 => x"FF",
		191880 => x"FF",
		192904 => x"FF",
		193928 => x"FF",
		194952 => x"FF",
		195976 => x"FF",
		197000 => x"FF",
		198024 => x"FF",
		199048 => x"FF",
		200072 => x"FF",
		201096 => x"FF",
		202120 => x"FF",
		203144 => x"FF",
		204168 => x"FF",
		205192 => x"FF",
		206216 => x"FF",
		207240 => x"FF",
		208264 => x"FF",
		209288 => x"FF",
		210312 => x"FF",
		211336 => x"FF",
		212360 => x"FF",
		213384 => x"FF",
		214408 => x"FF",
		215432 => x"FF",
		216456 => x"FF",
		217480 => x"FF",
		218504 => x"FF",
		219528 => x"FF",
		220552 => x"FF",
		221576 => x"FF",
		222600 => x"FF",
		223624 => x"FF",
		224648 => x"FF",
		225672 => x"FF",
		226696 => x"FF",
		227720 => x"FF",
		228744 => x"FF",
		229768 => x"FF",
		230792 => x"FF",
		231816 => x"FF",
		232840 => x"FF",
		233864 => x"FF",
		234888 => x"FF",
		235912 => x"FF",
		236936 => x"FF",
		237960 => x"FF",
		238984 => x"FF",
		240008 => x"FF",
		241032 => x"FF",
		242056 => x"FF",
		243080 => x"FF",
		244104 => x"FF",
		245128 => x"FF",
		246152 => x"FF",
		247176 => x"FF",
		248200 => x"FF",
		249224 => x"FF",
		250248 => x"FF",
		251272 => x"FF",
		252296 => x"FF",
		253320 => x"FF",
		254344 => x"FF",
		255368 => x"FF",
		256392 => x"FF",
		257416 => x"FF",
		258440 => x"FF",
		259464 => x"FF",
		260488 => x"FF",
		261512 => x"FF",
		262536 => x"FF",
		263560 => x"FF",
		264584 => x"FF",
		265608 => x"FF",
		266632 => x"FF",
		267656 => x"FF",
		268680 => x"FF",
		269704 => x"FF",
		270728 => x"FF",
		271752 => x"FF",
		272776 => x"FF",
		273800 => x"FF",
		274824 => x"FF",
		275848 => x"FF",
		276872 => x"FF",
		277896 => x"FF",
		278920 => x"FF",
		279944 => x"FF",
		280968 => x"FF",
		281992 => x"FF",
		283016 => x"FF",
		284040 => x"FF",
		285064 => x"FF",
		286088 => x"FF",
		287112 => x"FF",
		288136 => x"FF",
		289160 => x"FF",
		290184 => x"FF",
		291208 => x"FF",
		292232 => x"FF",
		293256 => x"FF",
		294280 => x"FF",
		295304 => x"FF",
		296328 => x"FF",
		297352 => x"FF",
		298376 => x"FF",
		299400 => x"FF",
		300424 => x"FF",
		301448 => x"FF",
		302472 => x"FF",
		303496 => x"FF",
		304520 => x"FF",
		305544 => x"FF",
		306568 => x"FF",
		307592 => x"FF",
		308616 => x"FF",
		309640 => x"FF",
		310664 => x"FF",
		311688 => x"FF",
		312712 => x"FF",
		313736 => x"FF",
		314760 => x"FF",
		315784 => x"FF",
		316808 => x"FF",
		317832 => x"FF",
		318856 => x"FF",
		319880 => x"FF",
		320904 => x"FF",
		321928 => x"FF",
		322952 => x"FF",
		323976 => x"FF",
		325000 => x"FF",
		326024 => x"FF",
		327048 => x"FF",
		328072 => x"FF",
		329096 => x"FF",
		330120 => x"FF",
		331144 => x"FF",
		332168 => x"FF",
		333192 => x"FF",
		334216 => x"FF",
		335240 => x"FF",
		336264 => x"FF",
		337288 => x"FF",
		338312 => x"FF",
		339336 => x"FF",
		340360 => x"FF",
		341384 => x"FF",
		342408 => x"FF",
		343432 => x"FF",
		344456 => x"FF",
		345480 => x"FF",
		346504 => x"FF",
		347528 => x"FF",
		348552 => x"FF",
		349576 => x"FF",
		350600 => x"FF",
		351624 => x"FF",
		352648 => x"FF",
		353672 => x"FF",
		354696 => x"FF",
		355720 => x"FF",
		356744 => x"FF",
		357768 => x"FF",
		358792 => x"FF",
		359816 => x"FF",
		360840 => x"FF",
		361864 => x"FF",
		362888 => x"FF",
		363912 => x"FF",
		364936 => x"FF",
		365960 => x"FF",
		366984 => x"FF",
		368008 => x"FF",
		369032 => x"FF",
		370056 => x"FF",
		371080 => x"FF",
		372104 => x"FF",
		373128 => x"FF",
		374152 => x"FF",
		375176 => x"FF",
		376200 => x"FF",
		377224 => x"FF",
		378248 => x"FF",
		379272 => x"FF",
		380296 => x"FF",
		381320 => x"FF",
		382344 => x"FF",
		383368 => x"FF",
		384392 => x"FF",
		385416 => x"FF",
		386440 => x"FF",
		387464 => x"FF",
		388488 => x"FF",
		389512 => x"FF",
		390536 => x"FF",
		391560 => x"FF",
		392584 => x"FF",
		393608 => x"FF",
		394632 => x"FF",
		395656 => x"FF",
		396680 => x"FF",
		397704 => x"FF",
		398728 => x"FF",
		399752 => x"FF",
		400776 => x"FF",
		401800 => x"FF",
		402824 => x"FF",
		403848 => x"FF",
		404872 => x"FF",
		405896 => x"FF",
		406920 => x"FF",
		407944 => x"FF",
		408968 => x"FF",
		409992 => x"FF",
		411016 => x"FF",
		412040 => x"FF",
		413064 => x"FF",
		414088 => x"FF",
		415112 => x"FF",
		416136 => x"FF",
		417160 => x"FF",
		418184 => x"FF",
		419208 => x"FF",
		420232 => x"FF",
		421256 => x"FF",
		422280 => x"FF",
		423304 => x"FF",
		424328 => x"FF",
		425352 => x"FF",
		426376 => x"FF",
		427400 => x"FF",
		428424 => x"FF",
		429448 => x"FF",
		430472 => x"FF",
		431496 => x"FF",
		432520 => x"FF",
		433544 => x"FF",
		434568 => x"FF",
		435592 => x"FF",
		436616 => x"FF",
		437640 => x"FF",
		438664 => x"FF",
		439688 => x"FF",
		440712 => x"FF",
		441736 => x"FF",
		442760 => x"FF",
		443784 => x"FF",
		444808 => x"FF",
		445832 => x"FF",
		446856 => x"FF",
		447880 => x"FF",
		448904 => x"FF",
		449928 => x"FF",
		450952 => x"FF",
		451976 => x"FF",
		453000 => x"FF",
		454024 => x"FF",
		455048 => x"FF",
		456072 => x"FF",
		457096 => x"FF",
		458120 => x"FF",
		459144 => x"FF",
		460168 => x"FF",
		461192 => x"FF",
		462216 => x"FF",
		463240 => x"FF",
		464264 => x"FF",
		465288 => x"FF",
		466312 => x"FF",
		467336 => x"FF",
		468360 => x"FF",
		469384 => x"FF",
		19849 => x"FF",
		20873 => x"FF",
		21897 => x"FF",
		22921 => x"FF",
		23945 => x"FF",
		24969 => x"FF",
		25993 => x"FF",
		27017 => x"FF",
		28041 => x"FF",
		29065 => x"FF",
		30089 => x"FF",
		31113 => x"FF",
		32137 => x"FF",
		33161 => x"FF",
		34185 => x"FF",
		35209 => x"FF",
		36233 => x"FF",
		37257 => x"FF",
		38281 => x"FF",
		39305 => x"FF",
		40329 => x"FF",
		41353 => x"FF",
		42377 => x"FF",
		43401 => x"FF",
		44425 => x"FF",
		45449 => x"FF",
		46473 => x"FF",
		47497 => x"FF",
		48521 => x"FF",
		49545 => x"FF",
		50569 => x"FF",
		51593 => x"FF",
		52617 => x"FF",
		53641 => x"FF",
		54665 => x"FF",
		55689 => x"FF",
		56713 => x"FF",
		57737 => x"FF",
		58761 => x"FF",
		59785 => x"FF",
		60809 => x"FF",
		61833 => x"FF",
		62857 => x"FF",
		63881 => x"FF",
		64905 => x"FF",
		65929 => x"FF",
		66953 => x"FF",
		67977 => x"FF",
		69001 => x"FF",
		70025 => x"FF",
		71049 => x"FF",
		72073 => x"FF",
		73097 => x"FF",
		74121 => x"FF",
		75145 => x"FF",
		76169 => x"FF",
		77193 => x"FF",
		78217 => x"FF",
		79241 => x"FF",
		80265 => x"FF",
		81289 => x"FF",
		82313 => x"FF",
		83337 => x"FF",
		84361 => x"FF",
		85385 => x"FF",
		86409 => x"FF",
		87433 => x"FF",
		88457 => x"FF",
		89481 => x"FF",
		90505 => x"FF",
		91529 => x"FF",
		92553 => x"FF",
		93577 => x"FF",
		94601 => x"FF",
		95625 => x"FF",
		96649 => x"FF",
		97673 => x"FF",
		98697 => x"FF",
		99721 => x"FF",
		100745 => x"FF",
		101769 => x"FF",
		102793 => x"FF",
		103817 => x"FF",
		104841 => x"FF",
		105865 => x"FF",
		106889 => x"FF",
		107913 => x"FF",
		108937 => x"FF",
		109961 => x"FF",
		110985 => x"FF",
		112009 => x"FF",
		113033 => x"FF",
		114057 => x"FF",
		115081 => x"FF",
		116105 => x"FF",
		117129 => x"FF",
		118153 => x"FF",
		119177 => x"FF",
		120201 => x"FF",
		121225 => x"FF",
		122249 => x"FF",
		123273 => x"FF",
		124297 => x"FF",
		125321 => x"FF",
		126345 => x"FF",
		127369 => x"FF",
		128393 => x"FF",
		129417 => x"FF",
		130441 => x"FF",
		131465 => x"FF",
		132489 => x"FF",
		133513 => x"FF",
		134537 => x"FF",
		135561 => x"FF",
		136585 => x"FF",
		137609 => x"FF",
		138633 => x"FF",
		139657 => x"FF",
		140681 => x"FF",
		141705 => x"FF",
		142729 => x"FF",
		143753 => x"FF",
		144777 => x"FF",
		145801 => x"FF",
		146825 => x"FF",
		147849 => x"FF",
		148873 => x"FF",
		149897 => x"FF",
		150921 => x"FF",
		151945 => x"FF",
		152969 => x"FF",
		153993 => x"FF",
		155017 => x"FF",
		156041 => x"FF",
		157065 => x"FF",
		158089 => x"FF",
		159113 => x"FF",
		160137 => x"FF",
		161161 => x"FF",
		162185 => x"FF",
		163209 => x"FF",
		164233 => x"FF",
		165257 => x"FF",
		166281 => x"FF",
		167305 => x"FF",
		168329 => x"FF",
		169353 => x"FF",
		170377 => x"FF",
		171401 => x"FF",
		172425 => x"FF",
		173449 => x"FF",
		174473 => x"FF",
		175497 => x"FF",
		176521 => x"FF",
		177545 => x"FF",
		178569 => x"FF",
		179593 => x"FF",
		180617 => x"FF",
		181641 => x"FF",
		182665 => x"FF",
		183689 => x"FF",
		184713 => x"FF",
		185737 => x"FF",
		186761 => x"FF",
		187785 => x"FF",
		188809 => x"FF",
		189833 => x"FF",
		190857 => x"FF",
		191881 => x"FF",
		192905 => x"FF",
		193929 => x"FF",
		194953 => x"FF",
		195977 => x"FF",
		197001 => x"FF",
		198025 => x"FF",
		199049 => x"FF",
		200073 => x"FF",
		201097 => x"FF",
		202121 => x"FF",
		203145 => x"FF",
		204169 => x"FF",
		205193 => x"FF",
		206217 => x"FF",
		207241 => x"FF",
		208265 => x"FF",
		209289 => x"FF",
		210313 => x"FF",
		211337 => x"FF",
		212361 => x"FF",
		213385 => x"FF",
		214409 => x"FF",
		215433 => x"FF",
		216457 => x"FF",
		217481 => x"FF",
		218505 => x"FF",
		219529 => x"FF",
		220553 => x"FF",
		221577 => x"FF",
		222601 => x"FF",
		223625 => x"FF",
		224649 => x"FF",
		225673 => x"FF",
		226697 => x"FF",
		227721 => x"FF",
		228745 => x"FF",
		229769 => x"FF",
		230793 => x"FF",
		231817 => x"FF",
		232841 => x"FF",
		233865 => x"FF",
		234889 => x"FF",
		235913 => x"FF",
		236937 => x"FF",
		237961 => x"FF",
		238985 => x"FF",
		240009 => x"FF",
		241033 => x"FF",
		242057 => x"FF",
		243081 => x"FF",
		244105 => x"FF",
		245129 => x"FF",
		246153 => x"FF",
		247177 => x"FF",
		248201 => x"FF",
		249225 => x"FF",
		250249 => x"FF",
		251273 => x"FF",
		252297 => x"FF",
		253321 => x"FF",
		254345 => x"FF",
		255369 => x"FF",
		256393 => x"FF",
		257417 => x"FF",
		258441 => x"FF",
		259465 => x"FF",
		260489 => x"FF",
		261513 => x"FF",
		262537 => x"FF",
		263561 => x"FF",
		264585 => x"FF",
		265609 => x"FF",
		266633 => x"FF",
		267657 => x"FF",
		268681 => x"FF",
		269705 => x"FF",
		270729 => x"FF",
		271753 => x"FF",
		272777 => x"FF",
		273801 => x"FF",
		274825 => x"FF",
		275849 => x"FF",
		276873 => x"FF",
		277897 => x"FF",
		278921 => x"FF",
		279945 => x"FF",
		280969 => x"FF",
		281993 => x"FF",
		283017 => x"FF",
		284041 => x"FF",
		285065 => x"FF",
		286089 => x"FF",
		287113 => x"FF",
		288137 => x"FF",
		289161 => x"FF",
		290185 => x"FF",
		291209 => x"FF",
		292233 => x"FF",
		293257 => x"FF",
		294281 => x"FF",
		295305 => x"FF",
		296329 => x"FF",
		297353 => x"FF",
		298377 => x"FF",
		299401 => x"FF",
		300425 => x"FF",
		301449 => x"FF",
		302473 => x"FF",
		303497 => x"FF",
		304521 => x"FF",
		305545 => x"FF",
		306569 => x"FF",
		307593 => x"FF",
		308617 => x"FF",
		309641 => x"FF",
		310665 => x"FF",
		311689 => x"FF",
		312713 => x"FF",
		313737 => x"FF",
		314761 => x"FF",
		315785 => x"FF",
		316809 => x"FF",
		317833 => x"FF",
		318857 => x"FF",
		319881 => x"FF",
		320905 => x"FF",
		321929 => x"FF",
		322953 => x"FF",
		323977 => x"FF",
		325001 => x"FF",
		326025 => x"FF",
		327049 => x"FF",
		328073 => x"FF",
		329097 => x"FF",
		330121 => x"FF",
		331145 => x"FF",
		332169 => x"FF",
		333193 => x"FF",
		334217 => x"FF",
		335241 => x"FF",
		336265 => x"FF",
		337289 => x"FF",
		338313 => x"FF",
		339337 => x"FF",
		340361 => x"FF",
		341385 => x"FF",
		342409 => x"FF",
		343433 => x"FF",
		344457 => x"FF",
		345481 => x"FF",
		346505 => x"FF",
		347529 => x"FF",
		348553 => x"FF",
		349577 => x"FF",
		350601 => x"FF",
		351625 => x"FF",
		352649 => x"FF",
		353673 => x"FF",
		354697 => x"FF",
		355721 => x"FF",
		356745 => x"FF",
		357769 => x"FF",
		358793 => x"FF",
		359817 => x"FF",
		360841 => x"FF",
		361865 => x"FF",
		362889 => x"FF",
		363913 => x"FF",
		364937 => x"FF",
		365961 => x"FF",
		366985 => x"FF",
		368009 => x"FF",
		369033 => x"FF",
		370057 => x"FF",
		371081 => x"FF",
		372105 => x"FF",
		373129 => x"FF",
		374153 => x"FF",
		375177 => x"FF",
		376201 => x"FF",
		377225 => x"FF",
		378249 => x"FF",
		379273 => x"FF",
		380297 => x"FF",
		381321 => x"FF",
		382345 => x"FF",
		383369 => x"FF",
		384393 => x"FF",
		385417 => x"FF",
		386441 => x"FF",
		387465 => x"FF",
		388489 => x"FF",
		389513 => x"FF",
		390537 => x"FF",
		391561 => x"FF",
		392585 => x"FF",
		393609 => x"FF",
		394633 => x"FF",
		395657 => x"FF",
		396681 => x"FF",
		397705 => x"FF",
		398729 => x"FF",
		399753 => x"FF",
		400777 => x"FF",
		401801 => x"FF",
		402825 => x"FF",
		403849 => x"FF",
		404873 => x"FF",
		405897 => x"FF",
		406921 => x"FF",
		407945 => x"FF",
		408969 => x"FF",
		409993 => x"FF",
		411017 => x"FF",
		412041 => x"FF",
		413065 => x"FF",
		414089 => x"FF",
		415113 => x"FF",
		416137 => x"FF",
		417161 => x"FF",
		418185 => x"FF",
		419209 => x"FF",
		420233 => x"FF",
		421257 => x"FF",
		422281 => x"FF",
		423305 => x"FF",
		424329 => x"FF",
		425353 => x"FF",
		426377 => x"FF",
		427401 => x"FF",
		428425 => x"FF",
		429449 => x"FF",
		430473 => x"FF",
		431497 => x"FF",
		432521 => x"FF",
		433545 => x"FF",
		434569 => x"FF",
		435593 => x"FF",
		436617 => x"FF",
		437641 => x"FF",
		438665 => x"FF",
		439689 => x"FF",
		440713 => x"FF",
		441737 => x"FF",
		442761 => x"FF",
		443785 => x"FF",
		444809 => x"FF",
		445833 => x"FF",
		446857 => x"FF",
		447881 => x"FF",
		448905 => x"FF",
		449929 => x"FF",
		450953 => x"FF",
		451977 => x"FF",
		453001 => x"FF",
		454025 => x"FF",
		455049 => x"FF",
		456073 => x"FF",
		457097 => x"FF",
		458121 => x"FF",
		459145 => x"FF",
		460169 => x"FF",
		461193 => x"FF",
		462217 => x"FF",
		463241 => x"FF",
		464265 => x"FF",
		465289 => x"FF",
		466313 => x"FF",
		467337 => x"FF",
		468361 => x"FF",
		469385 => x"FF",
		19850 => x"FF",
		20874 => x"FF",
		21898 => x"FF",
		22922 => x"FF",
		23946 => x"FF",
		168330 => x"FF",
		169354 => x"FF",
		170378 => x"FF",
		171402 => x"FF",
		172426 => x"FF",
		316810 => x"FF",
		317834 => x"FF",
		318858 => x"FF",
		319882 => x"FF",
		320906 => x"FF",
		465290 => x"FF",
		466314 => x"FF",
		467338 => x"FF",
		468362 => x"FF",
		469386 => x"FF",
		19851 => x"FF",
		20875 => x"FF",
		21899 => x"FF",
		22923 => x"FF",
		23947 => x"FF",
		168331 => x"FF",
		169355 => x"FF",
		170379 => x"FF",
		171403 => x"FF",
		172427 => x"FF",
		316811 => x"FF",
		317835 => x"FF",
		318859 => x"FF",
		319883 => x"FF",
		320907 => x"FF",
		465291 => x"FF",
		466315 => x"FF",
		467339 => x"FF",
		468363 => x"FF",
		469387 => x"FF",
		19852 => x"FF",
		20876 => x"FF",
		21900 => x"FF",
		22924 => x"FF",
		23948 => x"FF",
		168332 => x"FF",
		169356 => x"FF",
		170380 => x"FF",
		171404 => x"FF",
		172428 => x"FF",
		316812 => x"FF",
		317836 => x"FF",
		318860 => x"FF",
		319884 => x"FF",
		320908 => x"FF",
		465292 => x"FF",
		466316 => x"FF",
		467340 => x"FF",
		468364 => x"FF",
		469388 => x"FF",
		19853 => x"FF",
		20877 => x"FF",
		21901 => x"FF",
		22925 => x"FF",
		23949 => x"FF",
		168333 => x"FF",
		169357 => x"FF",
		170381 => x"FF",
		171405 => x"FF",
		172429 => x"FF",
		316813 => x"FF",
		317837 => x"FF",
		318861 => x"FF",
		319885 => x"FF",
		320909 => x"FF",
		465293 => x"FF",
		466317 => x"FF",
		467341 => x"FF",
		468365 => x"FF",
		469389 => x"FF",
		19854 => x"FF",
		20878 => x"FF",
		21902 => x"FF",
		22926 => x"FF",
		23950 => x"FF",
		168334 => x"FF",
		169358 => x"FF",
		170382 => x"FF",
		171406 => x"FF",
		172430 => x"FF",
		316814 => x"FF",
		317838 => x"FF",
		318862 => x"FF",
		319886 => x"FF",
		320910 => x"FF",
		465294 => x"FF",
		466318 => x"FF",
		467342 => x"FF",
		468366 => x"FF",
		469390 => x"FF",
		19855 => x"FF",
		20879 => x"FF",
		21903 => x"FF",
		22927 => x"FF",
		23951 => x"FF",
		168335 => x"FF",
		169359 => x"FF",
		170383 => x"FF",
		171407 => x"FF",
		172431 => x"FF",
		316815 => x"FF",
		317839 => x"FF",
		318863 => x"FF",
		319887 => x"FF",
		320911 => x"FF",
		465295 => x"FF",
		466319 => x"FF",
		467343 => x"FF",
		468367 => x"FF",
		469391 => x"FF",
		19856 => x"FF",
		20880 => x"FF",
		21904 => x"FF",
		22928 => x"FF",
		23952 => x"FF",
		168336 => x"FF",
		169360 => x"FF",
		170384 => x"FF",
		171408 => x"FF",
		172432 => x"FF",
		316816 => x"FF",
		317840 => x"FF",
		318864 => x"FF",
		319888 => x"FF",
		320912 => x"FF",
		465296 => x"FF",
		466320 => x"FF",
		467344 => x"FF",
		468368 => x"FF",
		469392 => x"FF",
		19857 => x"FF",
		20881 => x"FF",
		21905 => x"FF",
		22929 => x"FF",
		23953 => x"FF",
		168337 => x"FF",
		169361 => x"FF",
		170385 => x"FF",
		171409 => x"FF",
		172433 => x"FF",
		316817 => x"FF",
		317841 => x"FF",
		318865 => x"FF",
		319889 => x"FF",
		320913 => x"FF",
		465297 => x"FF",
		466321 => x"FF",
		467345 => x"FF",
		468369 => x"FF",
		469393 => x"FF",
		19858 => x"FF",
		20882 => x"FF",
		21906 => x"FF",
		22930 => x"FF",
		23954 => x"FF",
		168338 => x"FF",
		169362 => x"FF",
		170386 => x"FF",
		171410 => x"FF",
		172434 => x"FF",
		316818 => x"FF",
		317842 => x"FF",
		318866 => x"FF",
		319890 => x"FF",
		320914 => x"FF",
		465298 => x"FF",
		466322 => x"FF",
		467346 => x"FF",
		468370 => x"FF",
		469394 => x"FF",
		19859 => x"FF",
		20883 => x"FF",
		21907 => x"FF",
		22931 => x"FF",
		23955 => x"FF",
		168339 => x"FF",
		169363 => x"FF",
		170387 => x"FF",
		171411 => x"FF",
		172435 => x"FF",
		316819 => x"FF",
		317843 => x"FF",
		318867 => x"FF",
		319891 => x"FF",
		320915 => x"FF",
		465299 => x"FF",
		466323 => x"FF",
		467347 => x"FF",
		468371 => x"FF",
		469395 => x"FF",
		19860 => x"FF",
		20884 => x"FF",
		21908 => x"FF",
		22932 => x"FF",
		23956 => x"FF",
		168340 => x"FF",
		169364 => x"FF",
		170388 => x"FF",
		171412 => x"FF",
		172436 => x"FF",
		316820 => x"FF",
		317844 => x"FF",
		318868 => x"FF",
		319892 => x"FF",
		320916 => x"FF",
		465300 => x"FF",
		466324 => x"FF",
		467348 => x"FF",
		468372 => x"FF",
		469396 => x"FF",
		19861 => x"FF",
		20885 => x"FF",
		21909 => x"FF",
		22933 => x"FF",
		23957 => x"FF",
		168341 => x"FF",
		169365 => x"FF",
		170389 => x"FF",
		171413 => x"FF",
		172437 => x"FF",
		316821 => x"FF",
		317845 => x"FF",
		318869 => x"FF",
		319893 => x"FF",
		320917 => x"FF",
		465301 => x"FF",
		466325 => x"FF",
		467349 => x"FF",
		468373 => x"FF",
		469397 => x"FF",
		19862 => x"FF",
		20886 => x"FF",
		21910 => x"FF",
		22934 => x"FF",
		23958 => x"FF",
		168342 => x"FF",
		169366 => x"FF",
		170390 => x"FF",
		171414 => x"FF",
		172438 => x"FF",
		316822 => x"FF",
		317846 => x"FF",
		318870 => x"FF",
		319894 => x"FF",
		320918 => x"FF",
		465302 => x"FF",
		466326 => x"FF",
		467350 => x"FF",
		468374 => x"FF",
		469398 => x"FF",
		19863 => x"FF",
		20887 => x"FF",
		21911 => x"FF",
		22935 => x"FF",
		23959 => x"FF",
		168343 => x"FF",
		169367 => x"FF",
		170391 => x"FF",
		171415 => x"FF",
		172439 => x"FF",
		316823 => x"FF",
		317847 => x"FF",
		318871 => x"FF",
		319895 => x"FF",
		320919 => x"FF",
		465303 => x"FF",
		466327 => x"FF",
		467351 => x"FF",
		468375 => x"FF",
		469399 => x"FF",
		19864 => x"FF",
		20888 => x"FF",
		21912 => x"FF",
		22936 => x"FF",
		23960 => x"FF",
		168344 => x"FF",
		169368 => x"FF",
		170392 => x"FF",
		171416 => x"FF",
		172440 => x"FF",
		316824 => x"FF",
		317848 => x"FF",
		318872 => x"FF",
		319896 => x"FF",
		320920 => x"FF",
		465304 => x"FF",
		466328 => x"FF",
		467352 => x"FF",
		468376 => x"FF",
		469400 => x"FF",
		19865 => x"FF",
		20889 => x"FF",
		21913 => x"FF",
		22937 => x"FF",
		23961 => x"FF",
		168345 => x"FF",
		169369 => x"FF",
		170393 => x"FF",
		171417 => x"FF",
		172441 => x"FF",
		316825 => x"FF",
		317849 => x"FF",
		318873 => x"FF",
		319897 => x"FF",
		320921 => x"FF",
		465305 => x"FF",
		466329 => x"FF",
		467353 => x"FF",
		468377 => x"FF",
		469401 => x"FF",
		19866 => x"FF",
		20890 => x"FF",
		21914 => x"FF",
		22938 => x"FF",
		23962 => x"FF",
		168346 => x"FF",
		169370 => x"FF",
		170394 => x"FF",
		171418 => x"FF",
		172442 => x"FF",
		316826 => x"FF",
		317850 => x"FF",
		318874 => x"FF",
		319898 => x"FF",
		320922 => x"FF",
		465306 => x"FF",
		466330 => x"FF",
		467354 => x"FF",
		468378 => x"FF",
		469402 => x"FF",
		19867 => x"FF",
		20891 => x"FF",
		21915 => x"FF",
		22939 => x"FF",
		23963 => x"FF",
		168347 => x"FF",
		169371 => x"FF",
		170395 => x"FF",
		171419 => x"FF",
		172443 => x"FF",
		316827 => x"FF",
		317851 => x"FF",
		318875 => x"FF",
		319899 => x"FF",
		320923 => x"FF",
		465307 => x"FF",
		466331 => x"FF",
		467355 => x"FF",
		468379 => x"FF",
		469403 => x"FF",
		19868 => x"FF",
		20892 => x"FF",
		21916 => x"FF",
		22940 => x"FF",
		23964 => x"FF",
		168348 => x"FF",
		169372 => x"FF",
		170396 => x"FF",
		171420 => x"FF",
		172444 => x"FF",
		316828 => x"FF",
		317852 => x"FF",
		318876 => x"FF",
		319900 => x"FF",
		320924 => x"FF",
		465308 => x"FF",
		466332 => x"FF",
		467356 => x"FF",
		468380 => x"FF",
		469404 => x"FF",
		19869 => x"FF",
		20893 => x"FF",
		21917 => x"FF",
		22941 => x"FF",
		23965 => x"FF",
		168349 => x"FF",
		169373 => x"FF",
		170397 => x"FF",
		171421 => x"FF",
		172445 => x"FF",
		316829 => x"FF",
		317853 => x"FF",
		318877 => x"FF",
		319901 => x"FF",
		320925 => x"FF",
		465309 => x"FF",
		466333 => x"FF",
		467357 => x"FF",
		468381 => x"FF",
		469405 => x"FF",
		19870 => x"FF",
		20894 => x"FF",
		21918 => x"FF",
		22942 => x"FF",
		23966 => x"FF",
		168350 => x"FF",
		169374 => x"FF",
		170398 => x"FF",
		171422 => x"FF",
		172446 => x"FF",
		316830 => x"FF",
		317854 => x"FF",
		318878 => x"FF",
		319902 => x"FF",
		320926 => x"FF",
		465310 => x"FF",
		466334 => x"FF",
		467358 => x"FF",
		468382 => x"FF",
		469406 => x"FF",
		19871 => x"FF",
		20895 => x"FF",
		21919 => x"FF",
		22943 => x"FF",
		23967 => x"FF",
		168351 => x"FF",
		169375 => x"FF",
		170399 => x"FF",
		171423 => x"FF",
		172447 => x"FF",
		316831 => x"FF",
		317855 => x"FF",
		318879 => x"FF",
		319903 => x"FF",
		320927 => x"FF",
		465311 => x"FF",
		466335 => x"FF",
		467359 => x"FF",
		468383 => x"FF",
		469407 => x"FF",
		19872 => x"FF",
		20896 => x"FF",
		21920 => x"FF",
		22944 => x"FF",
		23968 => x"FF",
		168352 => x"FF",
		169376 => x"FF",
		170400 => x"FF",
		171424 => x"FF",
		172448 => x"FF",
		316832 => x"FF",
		317856 => x"FF",
		318880 => x"FF",
		319904 => x"FF",
		320928 => x"FF",
		465312 => x"FF",
		466336 => x"FF",
		467360 => x"FF",
		468384 => x"FF",
		469408 => x"FF",
		19873 => x"FF",
		20897 => x"FF",
		21921 => x"FF",
		22945 => x"FF",
		23969 => x"FF",
		168353 => x"FF",
		169377 => x"FF",
		170401 => x"FF",
		171425 => x"FF",
		172449 => x"FF",
		316833 => x"FF",
		317857 => x"FF",
		318881 => x"FF",
		319905 => x"FF",
		320929 => x"FF",
		465313 => x"FF",
		466337 => x"FF",
		467361 => x"FF",
		468385 => x"FF",
		469409 => x"FF",
		19874 => x"FF",
		20898 => x"FF",
		21922 => x"FF",
		22946 => x"FF",
		23970 => x"FF",
		168354 => x"FF",
		169378 => x"FF",
		170402 => x"FF",
		171426 => x"FF",
		172450 => x"FF",
		316834 => x"FF",
		317858 => x"FF",
		318882 => x"FF",
		319906 => x"FF",
		320930 => x"FF",
		465314 => x"FF",
		466338 => x"FF",
		467362 => x"FF",
		468386 => x"FF",
		469410 => x"FF",
		19875 => x"FF",
		20899 => x"FF",
		21923 => x"FF",
		22947 => x"FF",
		23971 => x"FF",
		168355 => x"FF",
		169379 => x"FF",
		170403 => x"FF",
		171427 => x"FF",
		172451 => x"FF",
		316835 => x"FF",
		317859 => x"FF",
		318883 => x"FF",
		319907 => x"FF",
		320931 => x"FF",
		465315 => x"FF",
		466339 => x"FF",
		467363 => x"FF",
		468387 => x"FF",
		469411 => x"FF",
		19876 => x"FF",
		20900 => x"FF",
		21924 => x"FF",
		22948 => x"FF",
		23972 => x"FF",
		168356 => x"FF",
		169380 => x"FF",
		170404 => x"FF",
		171428 => x"FF",
		172452 => x"FF",
		316836 => x"FF",
		317860 => x"FF",
		318884 => x"FF",
		319908 => x"FF",
		320932 => x"FF",
		465316 => x"FF",
		466340 => x"FF",
		467364 => x"FF",
		468388 => x"FF",
		469412 => x"FF",
		19877 => x"FF",
		20901 => x"FF",
		21925 => x"FF",
		22949 => x"FF",
		23973 => x"FF",
		168357 => x"FF",
		169381 => x"FF",
		170405 => x"FF",
		171429 => x"FF",
		172453 => x"FF",
		316837 => x"FF",
		317861 => x"FF",
		318885 => x"FF",
		319909 => x"FF",
		320933 => x"FF",
		465317 => x"FF",
		466341 => x"FF",
		467365 => x"FF",
		468389 => x"FF",
		469413 => x"FF",
		19878 => x"FF",
		20902 => x"FF",
		21926 => x"FF",
		22950 => x"FF",
		23974 => x"FF",
		168358 => x"FF",
		169382 => x"FF",
		170406 => x"FF",
		171430 => x"FF",
		172454 => x"FF",
		316838 => x"FF",
		317862 => x"FF",
		318886 => x"FF",
		319910 => x"FF",
		320934 => x"FF",
		465318 => x"FF",
		466342 => x"FF",
		467366 => x"FF",
		468390 => x"FF",
		469414 => x"FF",
		19879 => x"FF",
		20903 => x"FF",
		21927 => x"FF",
		22951 => x"FF",
		23975 => x"FF",
		168359 => x"FF",
		169383 => x"FF",
		170407 => x"FF",
		171431 => x"FF",
		172455 => x"FF",
		316839 => x"FF",
		317863 => x"FF",
		318887 => x"FF",
		319911 => x"FF",
		320935 => x"FF",
		465319 => x"FF",
		466343 => x"FF",
		467367 => x"FF",
		468391 => x"FF",
		469415 => x"FF",
		19880 => x"FF",
		20904 => x"FF",
		21928 => x"FF",
		22952 => x"FF",
		23976 => x"FF",
		168360 => x"FF",
		169384 => x"FF",
		170408 => x"FF",
		171432 => x"FF",
		172456 => x"FF",
		316840 => x"FF",
		317864 => x"FF",
		318888 => x"FF",
		319912 => x"FF",
		320936 => x"FF",
		465320 => x"FF",
		466344 => x"FF",
		467368 => x"FF",
		468392 => x"FF",
		469416 => x"FF",
		19881 => x"FF",
		20905 => x"FF",
		21929 => x"FF",
		22953 => x"FF",
		23977 => x"FF",
		168361 => x"FF",
		169385 => x"FF",
		170409 => x"FF",
		171433 => x"FF",
		172457 => x"FF",
		316841 => x"FF",
		317865 => x"FF",
		318889 => x"FF",
		319913 => x"FF",
		320937 => x"FF",
		465321 => x"FF",
		466345 => x"FF",
		467369 => x"FF",
		468393 => x"FF",
		469417 => x"FF",
		19882 => x"FF",
		20906 => x"FF",
		21930 => x"FF",
		22954 => x"FF",
		23978 => x"FF",
		168362 => x"FF",
		169386 => x"FF",
		170410 => x"FF",
		171434 => x"FF",
		172458 => x"FF",
		316842 => x"FF",
		317866 => x"FF",
		318890 => x"FF",
		319914 => x"FF",
		320938 => x"FF",
		465322 => x"FF",
		466346 => x"FF",
		467370 => x"FF",
		468394 => x"FF",
		469418 => x"FF",
		19883 => x"FF",
		20907 => x"FF",
		21931 => x"FF",
		22955 => x"FF",
		23979 => x"FF",
		168363 => x"FF",
		169387 => x"FF",
		170411 => x"FF",
		171435 => x"FF",
		172459 => x"FF",
		316843 => x"FF",
		317867 => x"FF",
		318891 => x"FF",
		319915 => x"FF",
		320939 => x"FF",
		465323 => x"FF",
		466347 => x"FF",
		467371 => x"FF",
		468395 => x"FF",
		469419 => x"FF",
		19884 => x"FF",
		20908 => x"FF",
		21932 => x"FF",
		22956 => x"FF",
		23980 => x"FF",
		168364 => x"FF",
		169388 => x"FF",
		170412 => x"FF",
		171436 => x"FF",
		172460 => x"FF",
		316844 => x"FF",
		317868 => x"FF",
		318892 => x"FF",
		319916 => x"FF",
		320940 => x"FF",
		465324 => x"FF",
		466348 => x"FF",
		467372 => x"FF",
		468396 => x"FF",
		469420 => x"FF",
		19885 => x"FF",
		20909 => x"FF",
		21933 => x"FF",
		22957 => x"FF",
		23981 => x"FF",
		168365 => x"FF",
		169389 => x"FF",
		170413 => x"FF",
		171437 => x"FF",
		172461 => x"FF",
		316845 => x"FF",
		317869 => x"FF",
		318893 => x"FF",
		319917 => x"FF",
		320941 => x"FF",
		465325 => x"FF",
		466349 => x"FF",
		467373 => x"FF",
		468397 => x"FF",
		469421 => x"FF",
		19886 => x"FF",
		20910 => x"FF",
		21934 => x"FF",
		22958 => x"FF",
		23982 => x"FF",
		168366 => x"FF",
		169390 => x"FF",
		170414 => x"FF",
		171438 => x"FF",
		172462 => x"FF",
		316846 => x"FF",
		317870 => x"FF",
		318894 => x"FF",
		319918 => x"FF",
		320942 => x"FF",
		465326 => x"FF",
		466350 => x"FF",
		467374 => x"FF",
		468398 => x"FF",
		469422 => x"FF",
		19887 => x"FF",
		20911 => x"FF",
		21935 => x"FF",
		22959 => x"FF",
		23983 => x"FF",
		168367 => x"FF",
		169391 => x"FF",
		170415 => x"FF",
		171439 => x"FF",
		172463 => x"FF",
		316847 => x"FF",
		317871 => x"FF",
		318895 => x"FF",
		319919 => x"FF",
		320943 => x"FF",
		465327 => x"FF",
		466351 => x"FF",
		467375 => x"FF",
		468399 => x"FF",
		469423 => x"FF",
		19888 => x"FF",
		20912 => x"FF",
		21936 => x"FF",
		22960 => x"FF",
		23984 => x"FF",
		168368 => x"FF",
		169392 => x"FF",
		170416 => x"FF",
		171440 => x"FF",
		172464 => x"FF",
		316848 => x"FF",
		317872 => x"FF",
		318896 => x"FF",
		319920 => x"FF",
		320944 => x"FF",
		465328 => x"FF",
		466352 => x"FF",
		467376 => x"FF",
		468400 => x"FF",
		469424 => x"FF",
		19889 => x"FF",
		20913 => x"FF",
		21937 => x"FF",
		22961 => x"FF",
		23985 => x"FF",
		168369 => x"FF",
		169393 => x"FF",
		170417 => x"FF",
		171441 => x"FF",
		172465 => x"FF",
		316849 => x"FF",
		317873 => x"FF",
		318897 => x"FF",
		319921 => x"FF",
		320945 => x"FF",
		465329 => x"FF",
		466353 => x"FF",
		467377 => x"FF",
		468401 => x"FF",
		469425 => x"FF",
		19890 => x"FF",
		20914 => x"FF",
		21938 => x"FF",
		22962 => x"FF",
		23986 => x"FF",
		168370 => x"FF",
		169394 => x"FF",
		170418 => x"FF",
		171442 => x"FF",
		172466 => x"FF",
		316850 => x"FF",
		317874 => x"FF",
		318898 => x"FF",
		319922 => x"FF",
		320946 => x"FF",
		465330 => x"FF",
		466354 => x"FF",
		467378 => x"FF",
		468402 => x"FF",
		469426 => x"FF",
		19891 => x"FF",
		20915 => x"FF",
		21939 => x"FF",
		22963 => x"FF",
		23987 => x"FF",
		168371 => x"FF",
		169395 => x"FF",
		170419 => x"FF",
		171443 => x"FF",
		172467 => x"FF",
		316851 => x"FF",
		317875 => x"FF",
		318899 => x"FF",
		319923 => x"FF",
		320947 => x"FF",
		465331 => x"FF",
		466355 => x"FF",
		467379 => x"FF",
		468403 => x"FF",
		469427 => x"FF",
		19892 => x"FF",
		20916 => x"FF",
		21940 => x"FF",
		22964 => x"FF",
		23988 => x"FF",
		168372 => x"FF",
		169396 => x"FF",
		170420 => x"FF",
		171444 => x"FF",
		172468 => x"FF",
		316852 => x"FF",
		317876 => x"FF",
		318900 => x"FF",
		319924 => x"FF",
		320948 => x"FF",
		465332 => x"FF",
		466356 => x"FF",
		467380 => x"FF",
		468404 => x"FF",
		469428 => x"FF",
		19893 => x"FF",
		20917 => x"FF",
		21941 => x"FF",
		22965 => x"FF",
		23989 => x"FF",
		168373 => x"FF",
		169397 => x"FF",
		170421 => x"FF",
		171445 => x"FF",
		172469 => x"FF",
		316853 => x"FF",
		317877 => x"FF",
		318901 => x"FF",
		319925 => x"FF",
		320949 => x"FF",
		465333 => x"FF",
		466357 => x"FF",
		467381 => x"FF",
		468405 => x"FF",
		469429 => x"FF",
		19894 => x"FF",
		20918 => x"FF",
		21942 => x"FF",
		22966 => x"FF",
		23990 => x"FF",
		168374 => x"FF",
		169398 => x"FF",
		170422 => x"FF",
		171446 => x"FF",
		172470 => x"FF",
		316854 => x"FF",
		317878 => x"FF",
		318902 => x"FF",
		319926 => x"FF",
		320950 => x"FF",
		465334 => x"FF",
		466358 => x"FF",
		467382 => x"FF",
		468406 => x"FF",
		469430 => x"FF",
		19895 => x"FF",
		20919 => x"FF",
		21943 => x"FF",
		22967 => x"FF",
		23991 => x"FF",
		168375 => x"FF",
		169399 => x"FF",
		170423 => x"FF",
		171447 => x"FF",
		172471 => x"FF",
		316855 => x"FF",
		317879 => x"FF",
		318903 => x"FF",
		319927 => x"FF",
		320951 => x"FF",
		465335 => x"FF",
		466359 => x"FF",
		467383 => x"FF",
		468407 => x"FF",
		469431 => x"FF",
		19896 => x"FF",
		20920 => x"FF",
		21944 => x"FF",
		22968 => x"FF",
		23992 => x"FF",
		168376 => x"FF",
		169400 => x"FF",
		170424 => x"FF",
		171448 => x"FF",
		172472 => x"FF",
		316856 => x"FF",
		317880 => x"FF",
		318904 => x"FF",
		319928 => x"FF",
		320952 => x"FF",
		465336 => x"FF",
		466360 => x"FF",
		467384 => x"FF",
		468408 => x"FF",
		469432 => x"FF",
		19897 => x"FF",
		20921 => x"FF",
		21945 => x"FF",
		22969 => x"FF",
		23993 => x"FF",
		168377 => x"FF",
		169401 => x"FF",
		170425 => x"FF",
		171449 => x"FF",
		172473 => x"FF",
		316857 => x"FF",
		317881 => x"FF",
		318905 => x"FF",
		319929 => x"FF",
		320953 => x"FF",
		465337 => x"FF",
		466361 => x"FF",
		467385 => x"FF",
		468409 => x"FF",
		469433 => x"FF",
		19898 => x"FF",
		20922 => x"FF",
		21946 => x"FF",
		22970 => x"FF",
		23994 => x"FF",
		168378 => x"FF",
		169402 => x"FF",
		170426 => x"FF",
		171450 => x"FF",
		172474 => x"FF",
		316858 => x"FF",
		317882 => x"FF",
		318906 => x"FF",
		319930 => x"FF",
		320954 => x"FF",
		465338 => x"FF",
		466362 => x"FF",
		467386 => x"FF",
		468410 => x"FF",
		469434 => x"FF",
		19899 => x"FF",
		20923 => x"FF",
		21947 => x"FF",
		22971 => x"FF",
		23995 => x"FF",
		168379 => x"FF",
		169403 => x"FF",
		170427 => x"FF",
		171451 => x"FF",
		172475 => x"FF",
		316859 => x"FF",
		317883 => x"FF",
		318907 => x"FF",
		319931 => x"FF",
		320955 => x"FF",
		465339 => x"FF",
		466363 => x"FF",
		467387 => x"FF",
		468411 => x"FF",
		469435 => x"FF",
		19900 => x"FF",
		20924 => x"FF",
		21948 => x"FF",
		22972 => x"FF",
		23996 => x"FF",
		168380 => x"FF",
		169404 => x"FF",
		170428 => x"FF",
		171452 => x"FF",
		172476 => x"FF",
		316860 => x"FF",
		317884 => x"FF",
		318908 => x"FF",
		319932 => x"FF",
		320956 => x"FF",
		465340 => x"FF",
		466364 => x"FF",
		467388 => x"FF",
		468412 => x"FF",
		469436 => x"FF",
		19901 => x"FF",
		20925 => x"FF",
		21949 => x"FF",
		22973 => x"FF",
		23997 => x"FF",
		168381 => x"FF",
		169405 => x"FF",
		170429 => x"FF",
		171453 => x"FF",
		172477 => x"FF",
		316861 => x"FF",
		317885 => x"FF",
		318909 => x"FF",
		319933 => x"FF",
		320957 => x"FF",
		465341 => x"FF",
		466365 => x"FF",
		467389 => x"FF",
		468413 => x"FF",
		469437 => x"FF",
		19902 => x"FF",
		20926 => x"FF",
		21950 => x"FF",
		22974 => x"FF",
		23998 => x"FF",
		168382 => x"FF",
		169406 => x"FF",
		170430 => x"FF",
		171454 => x"FF",
		172478 => x"FF",
		316862 => x"FF",
		317886 => x"FF",
		318910 => x"FF",
		319934 => x"FF",
		320958 => x"FF",
		465342 => x"FF",
		466366 => x"FF",
		467390 => x"FF",
		468414 => x"FF",
		469438 => x"FF",
		19903 => x"FF",
		20927 => x"FF",
		21951 => x"FF",
		22975 => x"FF",
		23999 => x"FF",
		168383 => x"FF",
		169407 => x"FF",
		170431 => x"FF",
		171455 => x"FF",
		172479 => x"FF",
		316863 => x"FF",
		317887 => x"FF",
		318911 => x"FF",
		319935 => x"FF",
		320959 => x"FF",
		465343 => x"FF",
		466367 => x"FF",
		467391 => x"FF",
		468415 => x"FF",
		469439 => x"FF",
		19904 => x"FF",
		20928 => x"FF",
		21952 => x"FF",
		22976 => x"FF",
		24000 => x"FF",
		168384 => x"FF",
		169408 => x"FF",
		170432 => x"FF",
		171456 => x"FF",
		172480 => x"FF",
		316864 => x"FF",
		317888 => x"FF",
		318912 => x"FF",
		319936 => x"FF",
		320960 => x"FF",
		465344 => x"FF",
		466368 => x"FF",
		467392 => x"FF",
		468416 => x"FF",
		469440 => x"FF",
		19905 => x"FF",
		20929 => x"FF",
		21953 => x"FF",
		22977 => x"FF",
		24001 => x"FF",
		168385 => x"FF",
		169409 => x"FF",
		170433 => x"FF",
		171457 => x"FF",
		172481 => x"FF",
		316865 => x"FF",
		317889 => x"FF",
		318913 => x"FF",
		319937 => x"FF",
		320961 => x"FF",
		465345 => x"FF",
		466369 => x"FF",
		467393 => x"FF",
		468417 => x"FF",
		469441 => x"FF",
		19906 => x"FF",
		20930 => x"FF",
		21954 => x"FF",
		22978 => x"FF",
		24002 => x"FF",
		168386 => x"FF",
		169410 => x"FF",
		170434 => x"FF",
		171458 => x"FF",
		172482 => x"FF",
		316866 => x"FF",
		317890 => x"FF",
		318914 => x"FF",
		319938 => x"FF",
		320962 => x"FF",
		465346 => x"FF",
		466370 => x"FF",
		467394 => x"FF",
		468418 => x"FF",
		469442 => x"FF",
		19907 => x"FF",
		20931 => x"FF",
		21955 => x"FF",
		22979 => x"FF",
		24003 => x"FF",
		168387 => x"FF",
		169411 => x"FF",
		170435 => x"FF",
		171459 => x"FF",
		172483 => x"FF",
		316867 => x"FF",
		317891 => x"FF",
		318915 => x"FF",
		319939 => x"FF",
		320963 => x"FF",
		465347 => x"FF",
		466371 => x"FF",
		467395 => x"FF",
		468419 => x"FF",
		469443 => x"FF",
		19908 => x"FF",
		20932 => x"FF",
		21956 => x"FF",
		22980 => x"FF",
		24004 => x"FF",
		168388 => x"FF",
		169412 => x"FF",
		170436 => x"FF",
		171460 => x"FF",
		172484 => x"FF",
		316868 => x"FF",
		317892 => x"FF",
		318916 => x"FF",
		319940 => x"FF",
		320964 => x"FF",
		465348 => x"FF",
		466372 => x"FF",
		467396 => x"FF",
		468420 => x"FF",
		469444 => x"FF",
		19909 => x"FF",
		20933 => x"FF",
		21957 => x"FF",
		22981 => x"FF",
		24005 => x"FF",
		168389 => x"FF",
		169413 => x"FF",
		170437 => x"FF",
		171461 => x"FF",
		172485 => x"FF",
		316869 => x"FF",
		317893 => x"FF",
		318917 => x"FF",
		319941 => x"FF",
		320965 => x"FF",
		465349 => x"FF",
		466373 => x"FF",
		467397 => x"FF",
		468421 => x"FF",
		469445 => x"FF",
		19910 => x"FF",
		20934 => x"FF",
		21958 => x"FF",
		22982 => x"FF",
		24006 => x"FF",
		168390 => x"FF",
		169414 => x"FF",
		170438 => x"FF",
		171462 => x"FF",
		172486 => x"FF",
		316870 => x"FF",
		317894 => x"FF",
		318918 => x"FF",
		319942 => x"FF",
		320966 => x"FF",
		465350 => x"FF",
		466374 => x"FF",
		467398 => x"FF",
		468422 => x"FF",
		469446 => x"FF",
		19911 => x"FF",
		20935 => x"FF",
		21959 => x"FF",
		22983 => x"FF",
		24007 => x"FF",
		168391 => x"FF",
		169415 => x"FF",
		170439 => x"FF",
		171463 => x"FF",
		172487 => x"FF",
		316871 => x"FF",
		317895 => x"FF",
		318919 => x"FF",
		319943 => x"FF",
		320967 => x"FF",
		465351 => x"FF",
		466375 => x"FF",
		467399 => x"FF",
		468423 => x"FF",
		469447 => x"FF",
		19912 => x"FF",
		20936 => x"FF",
		21960 => x"FF",
		22984 => x"FF",
		24008 => x"FF",
		168392 => x"FF",
		169416 => x"FF",
		170440 => x"FF",
		171464 => x"FF",
		172488 => x"FF",
		316872 => x"FF",
		317896 => x"FF",
		318920 => x"FF",
		319944 => x"FF",
		320968 => x"FF",
		465352 => x"FF",
		466376 => x"FF",
		467400 => x"FF",
		468424 => x"FF",
		469448 => x"FF",
		19913 => x"FF",
		20937 => x"FF",
		21961 => x"FF",
		22985 => x"FF",
		24009 => x"FF",
		168393 => x"FF",
		169417 => x"FF",
		170441 => x"FF",
		171465 => x"FF",
		172489 => x"FF",
		316873 => x"FF",
		317897 => x"FF",
		318921 => x"FF",
		319945 => x"FF",
		320969 => x"FF",
		465353 => x"FF",
		466377 => x"FF",
		467401 => x"FF",
		468425 => x"FF",
		469449 => x"FF",
		19914 => x"FF",
		20938 => x"FF",
		21962 => x"FF",
		22986 => x"FF",
		24010 => x"FF",
		168394 => x"FF",
		169418 => x"FF",
		170442 => x"FF",
		171466 => x"FF",
		172490 => x"FF",
		316874 => x"FF",
		317898 => x"FF",
		318922 => x"FF",
		319946 => x"FF",
		320970 => x"FF",
		465354 => x"FF",
		466378 => x"FF",
		467402 => x"FF",
		468426 => x"FF",
		469450 => x"FF",
		19915 => x"FF",
		20939 => x"FF",
		21963 => x"FF",
		22987 => x"FF",
		24011 => x"FF",
		168395 => x"FF",
		169419 => x"FF",
		170443 => x"FF",
		171467 => x"FF",
		172491 => x"FF",
		316875 => x"FF",
		317899 => x"FF",
		318923 => x"FF",
		319947 => x"FF",
		320971 => x"FF",
		465355 => x"FF",
		466379 => x"FF",
		467403 => x"FF",
		468427 => x"FF",
		469451 => x"FF",
		19916 => x"FF",
		20940 => x"FF",
		21964 => x"FF",
		22988 => x"FF",
		24012 => x"FF",
		168396 => x"FF",
		169420 => x"FF",
		170444 => x"FF",
		171468 => x"FF",
		172492 => x"FF",
		316876 => x"FF",
		317900 => x"FF",
		318924 => x"FF",
		319948 => x"FF",
		320972 => x"FF",
		465356 => x"FF",
		466380 => x"FF",
		467404 => x"FF",
		468428 => x"FF",
		469452 => x"FF",
		19917 => x"FF",
		20941 => x"FF",
		21965 => x"FF",
		22989 => x"FF",
		24013 => x"FF",
		168397 => x"FF",
		169421 => x"FF",
		170445 => x"FF",
		171469 => x"FF",
		172493 => x"FF",
		316877 => x"FF",
		317901 => x"FF",
		318925 => x"FF",
		319949 => x"FF",
		320973 => x"FF",
		465357 => x"FF",
		466381 => x"FF",
		467405 => x"FF",
		468429 => x"FF",
		469453 => x"FF",
		19918 => x"FF",
		20942 => x"FF",
		21966 => x"FF",
		22990 => x"FF",
		24014 => x"FF",
		168398 => x"FF",
		169422 => x"FF",
		170446 => x"FF",
		171470 => x"FF",
		172494 => x"FF",
		316878 => x"FF",
		317902 => x"FF",
		318926 => x"FF",
		319950 => x"FF",
		320974 => x"FF",
		465358 => x"FF",
		466382 => x"FF",
		467406 => x"FF",
		468430 => x"FF",
		469454 => x"FF",
		19919 => x"FF",
		20943 => x"FF",
		21967 => x"FF",
		22991 => x"FF",
		24015 => x"FF",
		168399 => x"FF",
		169423 => x"FF",
		170447 => x"FF",
		171471 => x"FF",
		172495 => x"FF",
		316879 => x"FF",
		317903 => x"FF",
		318927 => x"FF",
		319951 => x"FF",
		320975 => x"FF",
		465359 => x"FF",
		466383 => x"FF",
		467407 => x"FF",
		468431 => x"FF",
		469455 => x"FF",
		19920 => x"FF",
		20944 => x"FF",
		21968 => x"FF",
		22992 => x"FF",
		24016 => x"FF",
		168400 => x"FF",
		169424 => x"FF",
		170448 => x"FF",
		171472 => x"FF",
		172496 => x"FF",
		316880 => x"FF",
		317904 => x"FF",
		318928 => x"FF",
		319952 => x"FF",
		320976 => x"FF",
		465360 => x"FF",
		466384 => x"FF",
		467408 => x"FF",
		468432 => x"FF",
		469456 => x"FF",
		19921 => x"FF",
		20945 => x"FF",
		21969 => x"FF",
		22993 => x"FF",
		24017 => x"FF",
		168401 => x"FF",
		169425 => x"FF",
		170449 => x"FF",
		171473 => x"FF",
		172497 => x"FF",
		316881 => x"FF",
		317905 => x"FF",
		318929 => x"FF",
		319953 => x"FF",
		320977 => x"FF",
		465361 => x"FF",
		466385 => x"FF",
		467409 => x"FF",
		468433 => x"FF",
		469457 => x"FF",
		19922 => x"FF",
		20946 => x"FF",
		21970 => x"FF",
		22994 => x"FF",
		24018 => x"FF",
		168402 => x"FF",
		169426 => x"FF",
		170450 => x"FF",
		171474 => x"FF",
		172498 => x"FF",
		316882 => x"FF",
		317906 => x"FF",
		318930 => x"FF",
		319954 => x"FF",
		320978 => x"FF",
		465362 => x"FF",
		466386 => x"FF",
		467410 => x"FF",
		468434 => x"FF",
		469458 => x"FF",
		19923 => x"FF",
		20947 => x"FF",
		21971 => x"FF",
		22995 => x"FF",
		24019 => x"FF",
		168403 => x"FF",
		169427 => x"FF",
		170451 => x"FF",
		171475 => x"FF",
		172499 => x"FF",
		316883 => x"FF",
		317907 => x"FF",
		318931 => x"FF",
		319955 => x"FF",
		320979 => x"FF",
		465363 => x"FF",
		466387 => x"FF",
		467411 => x"FF",
		468435 => x"FF",
		469459 => x"FF",
		19924 => x"FF",
		20948 => x"FF",
		21972 => x"FF",
		22996 => x"FF",
		24020 => x"FF",
		168404 => x"FF",
		169428 => x"FF",
		170452 => x"FF",
		171476 => x"FF",
		172500 => x"FF",
		316884 => x"FF",
		317908 => x"FF",
		318932 => x"FF",
		319956 => x"FF",
		320980 => x"FF",
		465364 => x"FF",
		466388 => x"FF",
		467412 => x"FF",
		468436 => x"FF",
		469460 => x"FF",
		19925 => x"FF",
		20949 => x"FF",
		21973 => x"FF",
		22997 => x"FF",
		24021 => x"FF",
		168405 => x"FF",
		169429 => x"FF",
		170453 => x"FF",
		171477 => x"FF",
		172501 => x"FF",
		316885 => x"FF",
		317909 => x"FF",
		318933 => x"FF",
		319957 => x"FF",
		320981 => x"FF",
		465365 => x"FF",
		466389 => x"FF",
		467413 => x"FF",
		468437 => x"FF",
		469461 => x"FF",
		19926 => x"FF",
		20950 => x"FF",
		21974 => x"FF",
		22998 => x"FF",
		24022 => x"FF",
		168406 => x"FF",
		169430 => x"FF",
		170454 => x"FF",
		171478 => x"FF",
		172502 => x"FF",
		316886 => x"FF",
		317910 => x"FF",
		318934 => x"FF",
		319958 => x"FF",
		320982 => x"FF",
		465366 => x"FF",
		466390 => x"FF",
		467414 => x"FF",
		468438 => x"FF",
		469462 => x"FF",
		19927 => x"FF",
		20951 => x"FF",
		21975 => x"FF",
		22999 => x"FF",
		24023 => x"FF",
		168407 => x"FF",
		169431 => x"FF",
		170455 => x"FF",
		171479 => x"FF",
		172503 => x"FF",
		316887 => x"FF",
		317911 => x"FF",
		318935 => x"FF",
		319959 => x"FF",
		320983 => x"FF",
		465367 => x"FF",
		466391 => x"FF",
		467415 => x"FF",
		468439 => x"FF",
		469463 => x"FF",
		19928 => x"FF",
		20952 => x"FF",
		21976 => x"FF",
		23000 => x"FF",
		24024 => x"FF",
		168408 => x"FF",
		169432 => x"FF",
		170456 => x"FF",
		171480 => x"FF",
		172504 => x"FF",
		316888 => x"FF",
		317912 => x"FF",
		318936 => x"FF",
		319960 => x"FF",
		320984 => x"FF",
		465368 => x"FF",
		466392 => x"FF",
		467416 => x"FF",
		468440 => x"FF",
		469464 => x"FF",
		19929 => x"FF",
		20953 => x"FF",
		21977 => x"FF",
		23001 => x"FF",
		24025 => x"FF",
		168409 => x"FF",
		169433 => x"FF",
		170457 => x"FF",
		171481 => x"FF",
		172505 => x"FF",
		316889 => x"FF",
		317913 => x"FF",
		318937 => x"FF",
		319961 => x"FF",
		320985 => x"FF",
		465369 => x"FF",
		466393 => x"FF",
		467417 => x"FF",
		468441 => x"FF",
		469465 => x"FF",
		19930 => x"FF",
		20954 => x"FF",
		21978 => x"FF",
		23002 => x"FF",
		24026 => x"FF",
		168410 => x"FF",
		169434 => x"FF",
		170458 => x"FF",
		171482 => x"FF",
		172506 => x"FF",
		316890 => x"FF",
		317914 => x"FF",
		318938 => x"FF",
		319962 => x"FF",
		320986 => x"FF",
		465370 => x"FF",
		466394 => x"FF",
		467418 => x"FF",
		468442 => x"FF",
		469466 => x"FF",
		19931 => x"FF",
		20955 => x"FF",
		21979 => x"FF",
		23003 => x"FF",
		24027 => x"FF",
		168411 => x"FF",
		169435 => x"FF",
		170459 => x"FF",
		171483 => x"FF",
		172507 => x"FF",
		316891 => x"FF",
		317915 => x"FF",
		318939 => x"FF",
		319963 => x"FF",
		320987 => x"FF",
		465371 => x"FF",
		466395 => x"FF",
		467419 => x"FF",
		468443 => x"FF",
		469467 => x"FF",
		19932 => x"FF",
		20956 => x"FF",
		21980 => x"FF",
		23004 => x"FF",
		24028 => x"FF",
		168412 => x"FF",
		169436 => x"FF",
		170460 => x"FF",
		171484 => x"FF",
		172508 => x"FF",
		316892 => x"FF",
		317916 => x"FF",
		318940 => x"FF",
		319964 => x"FF",
		320988 => x"FF",
		465372 => x"FF",
		466396 => x"FF",
		467420 => x"FF",
		468444 => x"FF",
		469468 => x"FF",
		19933 => x"FF",
		20957 => x"FF",
		21981 => x"FF",
		23005 => x"FF",
		24029 => x"FF",
		168413 => x"FF",
		169437 => x"FF",
		170461 => x"FF",
		171485 => x"FF",
		172509 => x"FF",
		316893 => x"FF",
		317917 => x"FF",
		318941 => x"FF",
		319965 => x"FF",
		320989 => x"FF",
		465373 => x"FF",
		466397 => x"FF",
		467421 => x"FF",
		468445 => x"FF",
		469469 => x"FF",
		19934 => x"FF",
		20958 => x"FF",
		21982 => x"FF",
		23006 => x"FF",
		24030 => x"FF",
		168414 => x"FF",
		169438 => x"FF",
		170462 => x"FF",
		171486 => x"FF",
		172510 => x"FF",
		316894 => x"FF",
		317918 => x"FF",
		318942 => x"FF",
		319966 => x"FF",
		320990 => x"FF",
		465374 => x"FF",
		466398 => x"FF",
		467422 => x"FF",
		468446 => x"FF",
		469470 => x"FF",
		19935 => x"FF",
		20959 => x"FF",
		21983 => x"FF",
		23007 => x"FF",
		24031 => x"FF",
		168415 => x"FF",
		169439 => x"FF",
		170463 => x"FF",
		171487 => x"FF",
		172511 => x"FF",
		316895 => x"FF",
		317919 => x"FF",
		318943 => x"FF",
		319967 => x"FF",
		320991 => x"FF",
		465375 => x"FF",
		466399 => x"FF",
		467423 => x"FF",
		468447 => x"FF",
		469471 => x"FF",
		19936 => x"FF",
		20960 => x"FF",
		21984 => x"FF",
		23008 => x"FF",
		24032 => x"FF",
		168416 => x"FF",
		169440 => x"FF",
		170464 => x"FF",
		171488 => x"FF",
		172512 => x"FF",
		316896 => x"FF",
		317920 => x"FF",
		318944 => x"FF",
		319968 => x"FF",
		320992 => x"FF",
		465376 => x"FF",
		466400 => x"FF",
		467424 => x"FF",
		468448 => x"FF",
		469472 => x"FF",
		19937 => x"FF",
		20961 => x"FF",
		21985 => x"FF",
		23009 => x"FF",
		24033 => x"FF",
		168417 => x"FF",
		169441 => x"FF",
		170465 => x"FF",
		171489 => x"FF",
		172513 => x"FF",
		316897 => x"FF",
		317921 => x"FF",
		318945 => x"FF",
		319969 => x"FF",
		320993 => x"FF",
		465377 => x"FF",
		466401 => x"FF",
		467425 => x"FF",
		468449 => x"FF",
		469473 => x"FF",
		19938 => x"FF",
		20962 => x"FF",
		21986 => x"FF",
		23010 => x"FF",
		24034 => x"FF",
		168418 => x"FF",
		169442 => x"FF",
		170466 => x"FF",
		171490 => x"FF",
		172514 => x"FF",
		316898 => x"FF",
		317922 => x"FF",
		318946 => x"FF",
		319970 => x"FF",
		320994 => x"FF",
		465378 => x"FF",
		466402 => x"FF",
		467426 => x"FF",
		468450 => x"FF",
		469474 => x"FF",
		19939 => x"FF",
		20963 => x"FF",
		21987 => x"FF",
		23011 => x"FF",
		24035 => x"FF",
		168419 => x"FF",
		169443 => x"FF",
		170467 => x"FF",
		171491 => x"FF",
		172515 => x"FF",
		316899 => x"FF",
		317923 => x"FF",
		318947 => x"FF",
		319971 => x"FF",
		320995 => x"FF",
		465379 => x"FF",
		466403 => x"FF",
		467427 => x"FF",
		468451 => x"FF",
		469475 => x"FF",
		19940 => x"FF",
		20964 => x"FF",
		21988 => x"FF",
		23012 => x"FF",
		24036 => x"FF",
		168420 => x"FF",
		169444 => x"FF",
		170468 => x"FF",
		171492 => x"FF",
		172516 => x"FF",
		316900 => x"FF",
		317924 => x"FF",
		318948 => x"FF",
		319972 => x"FF",
		320996 => x"FF",
		465380 => x"FF",
		466404 => x"FF",
		467428 => x"FF",
		468452 => x"FF",
		469476 => x"FF",
		19941 => x"FF",
		20965 => x"FF",
		21989 => x"FF",
		23013 => x"FF",
		24037 => x"FF",
		168421 => x"FF",
		169445 => x"FF",
		170469 => x"FF",
		171493 => x"FF",
		172517 => x"FF",
		316901 => x"FF",
		317925 => x"FF",
		318949 => x"FF",
		319973 => x"FF",
		320997 => x"FF",
		465381 => x"FF",
		466405 => x"FF",
		467429 => x"FF",
		468453 => x"FF",
		469477 => x"FF",
		19942 => x"FF",
		20966 => x"FF",
		21990 => x"FF",
		23014 => x"FF",
		24038 => x"FF",
		168422 => x"FF",
		169446 => x"FF",
		170470 => x"FF",
		171494 => x"FF",
		172518 => x"FF",
		316902 => x"FF",
		317926 => x"FF",
		318950 => x"FF",
		319974 => x"FF",
		320998 => x"FF",
		465382 => x"FF",
		466406 => x"FF",
		467430 => x"FF",
		468454 => x"FF",
		469478 => x"FF",
		19943 => x"FF",
		20967 => x"FF",
		21991 => x"FF",
		23015 => x"FF",
		24039 => x"FF",
		168423 => x"FF",
		169447 => x"FF",
		170471 => x"FF",
		171495 => x"FF",
		172519 => x"FF",
		316903 => x"FF",
		317927 => x"FF",
		318951 => x"FF",
		319975 => x"FF",
		320999 => x"FF",
		465383 => x"FF",
		466407 => x"FF",
		467431 => x"FF",
		468455 => x"FF",
		469479 => x"FF",
		19944 => x"FF",
		20968 => x"FF",
		21992 => x"FF",
		23016 => x"FF",
		24040 => x"FF",
		168424 => x"FF",
		169448 => x"FF",
		170472 => x"FF",
		171496 => x"FF",
		172520 => x"FF",
		316904 => x"FF",
		317928 => x"FF",
		318952 => x"FF",
		319976 => x"FF",
		321000 => x"FF",
		465384 => x"FF",
		466408 => x"FF",
		467432 => x"FF",
		468456 => x"FF",
		469480 => x"FF",
		19945 => x"FF",
		20969 => x"FF",
		21993 => x"FF",
		23017 => x"FF",
		24041 => x"FF",
		168425 => x"FF",
		169449 => x"FF",
		170473 => x"FF",
		171497 => x"FF",
		172521 => x"FF",
		316905 => x"FF",
		317929 => x"FF",
		318953 => x"FF",
		319977 => x"FF",
		321001 => x"FF",
		465385 => x"FF",
		466409 => x"FF",
		467433 => x"FF",
		468457 => x"FF",
		469481 => x"FF",
		19946 => x"FF",
		20970 => x"FF",
		21994 => x"FF",
		23018 => x"FF",
		24042 => x"FF",
		168426 => x"FF",
		169450 => x"FF",
		170474 => x"FF",
		171498 => x"FF",
		172522 => x"FF",
		316906 => x"FF",
		317930 => x"FF",
		318954 => x"FF",
		319978 => x"FF",
		321002 => x"FF",
		465386 => x"FF",
		466410 => x"FF",
		467434 => x"FF",
		468458 => x"FF",
		469482 => x"FF",
		19947 => x"FF",
		20971 => x"FF",
		21995 => x"FF",
		23019 => x"FF",
		24043 => x"FF",
		168427 => x"FF",
		169451 => x"FF",
		170475 => x"FF",
		171499 => x"FF",
		172523 => x"FF",
		316907 => x"FF",
		317931 => x"FF",
		318955 => x"FF",
		319979 => x"FF",
		321003 => x"FF",
		465387 => x"FF",
		466411 => x"FF",
		467435 => x"FF",
		468459 => x"FF",
		469483 => x"FF",
		19948 => x"FF",
		20972 => x"FF",
		21996 => x"FF",
		23020 => x"FF",
		24044 => x"FF",
		168428 => x"FF",
		169452 => x"FF",
		170476 => x"FF",
		171500 => x"FF",
		172524 => x"FF",
		316908 => x"FF",
		317932 => x"FF",
		318956 => x"FF",
		319980 => x"FF",
		321004 => x"FF",
		465388 => x"FF",
		466412 => x"FF",
		467436 => x"FF",
		468460 => x"FF",
		469484 => x"FF",
		19949 => x"FF",
		20973 => x"FF",
		21997 => x"FF",
		23021 => x"FF",
		24045 => x"FF",
		168429 => x"FF",
		169453 => x"FF",
		170477 => x"FF",
		171501 => x"FF",
		172525 => x"FF",
		316909 => x"FF",
		317933 => x"FF",
		318957 => x"FF",
		319981 => x"FF",
		321005 => x"FF",
		465389 => x"FF",
		466413 => x"FF",
		467437 => x"FF",
		468461 => x"FF",
		469485 => x"FF",
		19950 => x"FF",
		20974 => x"FF",
		21998 => x"FF",
		23022 => x"FF",
		24046 => x"FF",
		168430 => x"FF",
		169454 => x"FF",
		170478 => x"FF",
		171502 => x"FF",
		172526 => x"FF",
		316910 => x"FF",
		317934 => x"FF",
		318958 => x"FF",
		319982 => x"FF",
		321006 => x"FF",
		465390 => x"FF",
		466414 => x"FF",
		467438 => x"FF",
		468462 => x"FF",
		469486 => x"FF",
		19951 => x"FF",
		20975 => x"FF",
		21999 => x"FF",
		23023 => x"FF",
		24047 => x"FF",
		168431 => x"FF",
		169455 => x"FF",
		170479 => x"FF",
		171503 => x"FF",
		172527 => x"FF",
		316911 => x"FF",
		317935 => x"FF",
		318959 => x"FF",
		319983 => x"FF",
		321007 => x"FF",
		465391 => x"FF",
		466415 => x"FF",
		467439 => x"FF",
		468463 => x"FF",
		469487 => x"FF",
		19952 => x"FF",
		20976 => x"FF",
		22000 => x"FF",
		23024 => x"FF",
		24048 => x"FF",
		168432 => x"FF",
		169456 => x"FF",
		170480 => x"FF",
		171504 => x"FF",
		172528 => x"FF",
		316912 => x"FF",
		317936 => x"FF",
		318960 => x"FF",
		319984 => x"FF",
		321008 => x"FF",
		465392 => x"FF",
		466416 => x"FF",
		467440 => x"FF",
		468464 => x"FF",
		469488 => x"FF",
		19953 => x"FF",
		20977 => x"FF",
		22001 => x"FF",
		23025 => x"FF",
		24049 => x"FF",
		168433 => x"FF",
		169457 => x"FF",
		170481 => x"FF",
		171505 => x"FF",
		172529 => x"FF",
		316913 => x"FF",
		317937 => x"FF",
		318961 => x"FF",
		319985 => x"FF",
		321009 => x"FF",
		465393 => x"FF",
		466417 => x"FF",
		467441 => x"FF",
		468465 => x"FF",
		469489 => x"FF",
		19954 => x"FF",
		20978 => x"FF",
		22002 => x"FF",
		23026 => x"FF",
		24050 => x"FF",
		168434 => x"FF",
		169458 => x"FF",
		170482 => x"FF",
		171506 => x"FF",
		172530 => x"FF",
		316914 => x"FF",
		317938 => x"FF",
		318962 => x"FF",
		319986 => x"FF",
		321010 => x"FF",
		465394 => x"FF",
		466418 => x"FF",
		467442 => x"FF",
		468466 => x"FF",
		469490 => x"FF",
		19955 => x"FF",
		20979 => x"FF",
		22003 => x"FF",
		23027 => x"FF",
		24051 => x"FF",
		168435 => x"FF",
		169459 => x"FF",
		170483 => x"FF",
		171507 => x"FF",
		172531 => x"FF",
		316915 => x"FF",
		317939 => x"FF",
		318963 => x"FF",
		319987 => x"FF",
		321011 => x"FF",
		465395 => x"FF",
		466419 => x"FF",
		467443 => x"FF",
		468467 => x"FF",
		469491 => x"FF",
		19956 => x"FF",
		20980 => x"FF",
		22004 => x"FF",
		23028 => x"FF",
		24052 => x"FF",
		168436 => x"FF",
		169460 => x"FF",
		170484 => x"FF",
		171508 => x"FF",
		172532 => x"FF",
		316916 => x"FF",
		317940 => x"FF",
		318964 => x"FF",
		319988 => x"FF",
		321012 => x"FF",
		465396 => x"FF",
		466420 => x"FF",
		467444 => x"FF",
		468468 => x"FF",
		469492 => x"FF",
		19957 => x"FF",
		20981 => x"FF",
		22005 => x"FF",
		23029 => x"FF",
		24053 => x"FF",
		168437 => x"FF",
		169461 => x"FF",
		170485 => x"FF",
		171509 => x"FF",
		172533 => x"FF",
		316917 => x"FF",
		317941 => x"FF",
		318965 => x"FF",
		319989 => x"FF",
		321013 => x"FF",
		465397 => x"FF",
		466421 => x"FF",
		467445 => x"FF",
		468469 => x"FF",
		469493 => x"FF",
		19958 => x"FF",
		20982 => x"FF",
		22006 => x"FF",
		23030 => x"FF",
		24054 => x"FF",
		168438 => x"FF",
		169462 => x"FF",
		170486 => x"FF",
		171510 => x"FF",
		172534 => x"FF",
		316918 => x"FF",
		317942 => x"FF",
		318966 => x"FF",
		319990 => x"FF",
		321014 => x"FF",
		465398 => x"FF",
		466422 => x"FF",
		467446 => x"FF",
		468470 => x"FF",
		469494 => x"FF",
		19959 => x"FF",
		20983 => x"FF",
		22007 => x"FF",
		23031 => x"FF",
		24055 => x"FF",
		168439 => x"FF",
		169463 => x"FF",
		170487 => x"FF",
		171511 => x"FF",
		172535 => x"FF",
		316919 => x"FF",
		317943 => x"FF",
		318967 => x"FF",
		319991 => x"FF",
		321015 => x"FF",
		465399 => x"FF",
		466423 => x"FF",
		467447 => x"FF",
		468471 => x"FF",
		469495 => x"FF",
		19960 => x"FF",
		20984 => x"FF",
		22008 => x"FF",
		23032 => x"FF",
		24056 => x"FF",
		168440 => x"FF",
		169464 => x"FF",
		170488 => x"FF",
		171512 => x"FF",
		172536 => x"FF",
		316920 => x"FF",
		317944 => x"FF",
		318968 => x"FF",
		319992 => x"FF",
		321016 => x"FF",
		465400 => x"FF",
		466424 => x"FF",
		467448 => x"FF",
		468472 => x"FF",
		469496 => x"FF",
		19961 => x"FF",
		20985 => x"FF",
		22009 => x"FF",
		23033 => x"FF",
		24057 => x"FF",
		168441 => x"FF",
		169465 => x"FF",
		170489 => x"FF",
		171513 => x"FF",
		172537 => x"FF",
		316921 => x"FF",
		317945 => x"FF",
		318969 => x"FF",
		319993 => x"FF",
		321017 => x"FF",
		465401 => x"FF",
		466425 => x"FF",
		467449 => x"FF",
		468473 => x"FF",
		469497 => x"FF",
		19962 => x"FF",
		20986 => x"FF",
		22010 => x"FF",
		23034 => x"FF",
		24058 => x"FF",
		168442 => x"FF",
		169466 => x"FF",
		170490 => x"FF",
		171514 => x"FF",
		172538 => x"FF",
		316922 => x"FF",
		317946 => x"FF",
		318970 => x"FF",
		319994 => x"FF",
		321018 => x"FF",
		465402 => x"FF",
		466426 => x"FF",
		467450 => x"FF",
		468474 => x"FF",
		469498 => x"FF",
		19963 => x"FF",
		20987 => x"FF",
		22011 => x"FF",
		23035 => x"FF",
		24059 => x"FF",
		168443 => x"FF",
		169467 => x"FF",
		170491 => x"FF",
		171515 => x"FF",
		172539 => x"FF",
		316923 => x"FF",
		317947 => x"FF",
		318971 => x"FF",
		319995 => x"FF",
		321019 => x"FF",
		465403 => x"FF",
		466427 => x"FF",
		467451 => x"FF",
		468475 => x"FF",
		469499 => x"FF",
		19964 => x"FF",
		20988 => x"FF",
		22012 => x"FF",
		23036 => x"FF",
		24060 => x"FF",
		168444 => x"FF",
		169468 => x"FF",
		170492 => x"FF",
		171516 => x"FF",
		172540 => x"FF",
		316924 => x"FF",
		317948 => x"FF",
		318972 => x"FF",
		319996 => x"FF",
		321020 => x"FF",
		465404 => x"FF",
		466428 => x"FF",
		467452 => x"FF",
		468476 => x"FF",
		469500 => x"FF",
		19965 => x"FF",
		20989 => x"FF",
		22013 => x"FF",
		23037 => x"FF",
		24061 => x"FF",
		168445 => x"FF",
		169469 => x"FF",
		170493 => x"FF",
		171517 => x"FF",
		172541 => x"FF",
		316925 => x"FF",
		317949 => x"FF",
		318973 => x"FF",
		319997 => x"FF",
		321021 => x"FF",
		465405 => x"FF",
		466429 => x"FF",
		467453 => x"FF",
		468477 => x"FF",
		469501 => x"FF",
		19966 => x"FF",
		20990 => x"FF",
		22014 => x"FF",
		23038 => x"FF",
		24062 => x"FF",
		168446 => x"FF",
		169470 => x"FF",
		170494 => x"FF",
		171518 => x"FF",
		172542 => x"FF",
		316926 => x"FF",
		317950 => x"FF",
		318974 => x"FF",
		319998 => x"FF",
		321022 => x"FF",
		465406 => x"FF",
		466430 => x"FF",
		467454 => x"FF",
		468478 => x"FF",
		469502 => x"FF",
		19967 => x"FF",
		20991 => x"FF",
		22015 => x"FF",
		23039 => x"FF",
		24063 => x"FF",
		168447 => x"FF",
		169471 => x"FF",
		170495 => x"FF",
		171519 => x"FF",
		172543 => x"FF",
		316927 => x"FF",
		317951 => x"FF",
		318975 => x"FF",
		319999 => x"FF",
		321023 => x"FF",
		465407 => x"FF",
		466431 => x"FF",
		467455 => x"FF",
		468479 => x"FF",
		469503 => x"FF",
		19968 => x"FF",
		20992 => x"FF",
		22016 => x"FF",
		23040 => x"FF",
		24064 => x"FF",
		168448 => x"FF",
		169472 => x"FF",
		170496 => x"FF",
		171520 => x"FF",
		172544 => x"FF",
		316928 => x"FF",
		317952 => x"FF",
		318976 => x"FF",
		320000 => x"FF",
		321024 => x"FF",
		465408 => x"FF",
		466432 => x"FF",
		467456 => x"FF",
		468480 => x"FF",
		469504 => x"FF",
		19969 => x"FF",
		20993 => x"FF",
		22017 => x"FF",
		23041 => x"FF",
		24065 => x"FF",
		168449 => x"FF",
		169473 => x"FF",
		170497 => x"FF",
		171521 => x"FF",
		172545 => x"FF",
		316929 => x"FF",
		317953 => x"FF",
		318977 => x"FF",
		320001 => x"FF",
		321025 => x"FF",
		465409 => x"FF",
		466433 => x"FF",
		467457 => x"FF",
		468481 => x"FF",
		469505 => x"FF",
		19970 => x"FF",
		20994 => x"FF",
		22018 => x"FF",
		23042 => x"FF",
		24066 => x"FF",
		168450 => x"FF",
		169474 => x"FF",
		170498 => x"FF",
		171522 => x"FF",
		172546 => x"FF",
		316930 => x"FF",
		317954 => x"FF",
		318978 => x"FF",
		320002 => x"FF",
		321026 => x"FF",
		465410 => x"FF",
		466434 => x"FF",
		467458 => x"FF",
		468482 => x"FF",
		469506 => x"FF",
		19971 => x"FF",
		20995 => x"FF",
		22019 => x"FF",
		23043 => x"FF",
		24067 => x"FF",
		168451 => x"FF",
		169475 => x"FF",
		170499 => x"FF",
		171523 => x"FF",
		172547 => x"FF",
		316931 => x"FF",
		317955 => x"FF",
		318979 => x"FF",
		320003 => x"FF",
		321027 => x"FF",
		465411 => x"FF",
		466435 => x"FF",
		467459 => x"FF",
		468483 => x"FF",
		469507 => x"FF",
		19972 => x"FF",
		20996 => x"FF",
		22020 => x"FF",
		23044 => x"FF",
		24068 => x"FF",
		168452 => x"FF",
		169476 => x"FF",
		170500 => x"FF",
		171524 => x"FF",
		172548 => x"FF",
		316932 => x"FF",
		317956 => x"FF",
		318980 => x"FF",
		320004 => x"FF",
		321028 => x"FF",
		465412 => x"FF",
		466436 => x"FF",
		467460 => x"FF",
		468484 => x"FF",
		469508 => x"FF",
		19973 => x"FF",
		20997 => x"FF",
		22021 => x"FF",
		23045 => x"FF",
		24069 => x"FF",
		168453 => x"FF",
		169477 => x"FF",
		170501 => x"FF",
		171525 => x"FF",
		172549 => x"FF",
		316933 => x"FF",
		317957 => x"FF",
		318981 => x"FF",
		320005 => x"FF",
		321029 => x"FF",
		465413 => x"FF",
		466437 => x"FF",
		467461 => x"FF",
		468485 => x"FF",
		469509 => x"FF",
		19974 => x"FF",
		20998 => x"FF",
		22022 => x"FF",
		23046 => x"FF",
		24070 => x"FF",
		168454 => x"FF",
		169478 => x"FF",
		170502 => x"FF",
		171526 => x"FF",
		172550 => x"FF",
		316934 => x"FF",
		317958 => x"FF",
		318982 => x"FF",
		320006 => x"FF",
		321030 => x"FF",
		465414 => x"FF",
		466438 => x"FF",
		467462 => x"FF",
		468486 => x"FF",
		469510 => x"FF",
		19975 => x"FF",
		20999 => x"FF",
		22023 => x"FF",
		23047 => x"FF",
		24071 => x"FF",
		168455 => x"FF",
		169479 => x"FF",
		170503 => x"FF",
		171527 => x"FF",
		172551 => x"FF",
		316935 => x"FF",
		317959 => x"FF",
		318983 => x"FF",
		320007 => x"FF",
		321031 => x"FF",
		465415 => x"FF",
		466439 => x"FF",
		467463 => x"FF",
		468487 => x"FF",
		469511 => x"FF",
		19976 => x"FF",
		21000 => x"FF",
		22024 => x"FF",
		23048 => x"FF",
		24072 => x"FF",
		168456 => x"FF",
		169480 => x"FF",
		170504 => x"FF",
		171528 => x"FF",
		172552 => x"FF",
		316936 => x"FF",
		317960 => x"FF",
		318984 => x"FF",
		320008 => x"FF",
		321032 => x"FF",
		465416 => x"FF",
		466440 => x"FF",
		467464 => x"FF",
		468488 => x"FF",
		469512 => x"FF",
		19977 => x"FF",
		21001 => x"FF",
		22025 => x"FF",
		23049 => x"FF",
		24073 => x"FF",
		168457 => x"FF",
		169481 => x"FF",
		170505 => x"FF",
		171529 => x"FF",
		172553 => x"FF",
		316937 => x"FF",
		317961 => x"FF",
		318985 => x"FF",
		320009 => x"FF",
		321033 => x"FF",
		465417 => x"FF",
		466441 => x"FF",
		467465 => x"FF",
		468489 => x"FF",
		469513 => x"FF",
		19978 => x"FF",
		21002 => x"FF",
		22026 => x"FF",
		23050 => x"FF",
		24074 => x"FF",
		168458 => x"FF",
		169482 => x"FF",
		170506 => x"FF",
		171530 => x"FF",
		172554 => x"FF",
		316938 => x"FF",
		317962 => x"FF",
		318986 => x"FF",
		320010 => x"FF",
		321034 => x"FF",
		465418 => x"FF",
		466442 => x"FF",
		467466 => x"FF",
		468490 => x"FF",
		469514 => x"FF",
		19979 => x"FF",
		21003 => x"FF",
		22027 => x"FF",
		23051 => x"FF",
		24075 => x"FF",
		168459 => x"FF",
		169483 => x"FF",
		170507 => x"FF",
		171531 => x"FF",
		172555 => x"FF",
		316939 => x"FF",
		317963 => x"FF",
		318987 => x"FF",
		320011 => x"FF",
		321035 => x"FF",
		465419 => x"FF",
		466443 => x"FF",
		467467 => x"FF",
		468491 => x"FF",
		469515 => x"FF",
		19980 => x"FF",
		21004 => x"FF",
		22028 => x"FF",
		23052 => x"FF",
		24076 => x"FF",
		168460 => x"FF",
		169484 => x"FF",
		170508 => x"FF",
		171532 => x"FF",
		172556 => x"FF",
		316940 => x"FF",
		317964 => x"FF",
		318988 => x"FF",
		320012 => x"FF",
		321036 => x"FF",
		465420 => x"FF",
		466444 => x"FF",
		467468 => x"FF",
		468492 => x"FF",
		469516 => x"FF",
		19981 => x"FF",
		21005 => x"FF",
		22029 => x"FF",
		23053 => x"FF",
		24077 => x"FF",
		168461 => x"FF",
		169485 => x"FF",
		170509 => x"FF",
		171533 => x"FF",
		172557 => x"FF",
		316941 => x"FF",
		317965 => x"FF",
		318989 => x"FF",
		320013 => x"FF",
		321037 => x"FF",
		465421 => x"FF",
		466445 => x"FF",
		467469 => x"FF",
		468493 => x"FF",
		469517 => x"FF",
		19982 => x"FF",
		21006 => x"FF",
		22030 => x"FF",
		23054 => x"FF",
		24078 => x"FF",
		168462 => x"FF",
		169486 => x"FF",
		170510 => x"FF",
		171534 => x"FF",
		172558 => x"FF",
		316942 => x"FF",
		317966 => x"FF",
		318990 => x"FF",
		320014 => x"FF",
		321038 => x"FF",
		465422 => x"FF",
		466446 => x"FF",
		467470 => x"FF",
		468494 => x"FF",
		469518 => x"FF",
		19983 => x"FF",
		21007 => x"FF",
		22031 => x"FF",
		23055 => x"FF",
		24079 => x"FF",
		168463 => x"FF",
		169487 => x"FF",
		170511 => x"FF",
		171535 => x"FF",
		172559 => x"FF",
		316943 => x"FF",
		317967 => x"FF",
		318991 => x"FF",
		320015 => x"FF",
		321039 => x"FF",
		465423 => x"FF",
		466447 => x"FF",
		467471 => x"FF",
		468495 => x"FF",
		469519 => x"FF",
		19984 => x"FF",
		21008 => x"FF",
		22032 => x"FF",
		23056 => x"FF",
		24080 => x"FF",
		168464 => x"FF",
		169488 => x"FF",
		170512 => x"FF",
		171536 => x"FF",
		172560 => x"FF",
		316944 => x"FF",
		317968 => x"FF",
		318992 => x"FF",
		320016 => x"FF",
		321040 => x"FF",
		465424 => x"FF",
		466448 => x"FF",
		467472 => x"FF",
		468496 => x"FF",
		469520 => x"FF",
		19985 => x"FF",
		21009 => x"FF",
		22033 => x"FF",
		23057 => x"FF",
		24081 => x"FF",
		168465 => x"FF",
		169489 => x"FF",
		170513 => x"FF",
		171537 => x"FF",
		172561 => x"FF",
		316945 => x"FF",
		317969 => x"FF",
		318993 => x"FF",
		320017 => x"FF",
		321041 => x"FF",
		465425 => x"FF",
		466449 => x"FF",
		467473 => x"FF",
		468497 => x"FF",
		469521 => x"FF",
		19986 => x"FF",
		21010 => x"FF",
		22034 => x"FF",
		23058 => x"FF",
		24082 => x"FF",
		168466 => x"FF",
		169490 => x"FF",
		170514 => x"FF",
		171538 => x"FF",
		172562 => x"FF",
		316946 => x"FF",
		317970 => x"FF",
		318994 => x"FF",
		320018 => x"FF",
		321042 => x"FF",
		465426 => x"FF",
		466450 => x"FF",
		467474 => x"FF",
		468498 => x"FF",
		469522 => x"FF",
		19987 => x"FF",
		21011 => x"FF",
		22035 => x"FF",
		23059 => x"FF",
		24083 => x"FF",
		168467 => x"FF",
		169491 => x"FF",
		170515 => x"FF",
		171539 => x"FF",
		172563 => x"FF",
		316947 => x"FF",
		317971 => x"FF",
		318995 => x"FF",
		320019 => x"FF",
		321043 => x"FF",
		465427 => x"FF",
		466451 => x"FF",
		467475 => x"FF",
		468499 => x"FF",
		469523 => x"FF",
		19988 => x"FF",
		21012 => x"FF",
		22036 => x"FF",
		23060 => x"FF",
		24084 => x"FF",
		168468 => x"FF",
		169492 => x"FF",
		170516 => x"FF",
		171540 => x"FF",
		172564 => x"FF",
		316948 => x"FF",
		317972 => x"FF",
		318996 => x"FF",
		320020 => x"FF",
		321044 => x"FF",
		465428 => x"FF",
		466452 => x"FF",
		467476 => x"FF",
		468500 => x"FF",
		469524 => x"FF",
		19989 => x"FF",
		21013 => x"FF",
		22037 => x"FF",
		23061 => x"FF",
		24085 => x"FF",
		168469 => x"FF",
		169493 => x"FF",
		170517 => x"FF",
		171541 => x"FF",
		172565 => x"FF",
		316949 => x"FF",
		317973 => x"FF",
		318997 => x"FF",
		320021 => x"FF",
		321045 => x"FF",
		465429 => x"FF",
		466453 => x"FF",
		467477 => x"FF",
		468501 => x"FF",
		469525 => x"FF",
		19990 => x"FF",
		21014 => x"FF",
		22038 => x"FF",
		23062 => x"FF",
		24086 => x"FF",
		25110 => x"FF",
		26134 => x"FF",
		27158 => x"FF",
		28182 => x"FF",
		29206 => x"FF",
		30230 => x"FF",
		31254 => x"FF",
		32278 => x"FF",
		33302 => x"FF",
		34326 => x"FF",
		35350 => x"FF",
		36374 => x"FF",
		37398 => x"FF",
		38422 => x"FF",
		39446 => x"FF",
		40470 => x"FF",
		41494 => x"FF",
		42518 => x"FF",
		43542 => x"FF",
		44566 => x"FF",
		45590 => x"FF",
		46614 => x"FF",
		47638 => x"FF",
		48662 => x"FF",
		49686 => x"FF",
		50710 => x"FF",
		51734 => x"FF",
		52758 => x"FF",
		53782 => x"FF",
		54806 => x"FF",
		55830 => x"FF",
		56854 => x"FF",
		57878 => x"FF",
		58902 => x"FF",
		59926 => x"FF",
		60950 => x"FF",
		61974 => x"FF",
		62998 => x"FF",
		64022 => x"FF",
		65046 => x"FF",
		66070 => x"FF",
		67094 => x"FF",
		68118 => x"FF",
		69142 => x"FF",
		70166 => x"FF",
		71190 => x"FF",
		72214 => x"FF",
		73238 => x"FF",
		74262 => x"FF",
		75286 => x"FF",
		76310 => x"FF",
		77334 => x"FF",
		78358 => x"FF",
		79382 => x"FF",
		80406 => x"FF",
		81430 => x"FF",
		82454 => x"FF",
		83478 => x"FF",
		84502 => x"FF",
		85526 => x"FF",
		86550 => x"FF",
		87574 => x"FF",
		88598 => x"FF",
		89622 => x"FF",
		90646 => x"FF",
		91670 => x"FF",
		92694 => x"FF",
		93718 => x"FF",
		94742 => x"FF",
		95766 => x"FF",
		96790 => x"FF",
		97814 => x"FF",
		98838 => x"FF",
		99862 => x"FF",
		100886 => x"FF",
		101910 => x"FF",
		102934 => x"FF",
		103958 => x"FF",
		104982 => x"FF",
		106006 => x"FF",
		107030 => x"FF",
		108054 => x"FF",
		109078 => x"FF",
		110102 => x"FF",
		111126 => x"FF",
		112150 => x"FF",
		113174 => x"FF",
		114198 => x"FF",
		115222 => x"FF",
		116246 => x"FF",
		117270 => x"FF",
		118294 => x"FF",
		119318 => x"FF",
		120342 => x"FF",
		121366 => x"FF",
		122390 => x"FF",
		123414 => x"FF",
		124438 => x"FF",
		125462 => x"FF",
		126486 => x"FF",
		127510 => x"FF",
		128534 => x"FF",
		129558 => x"FF",
		130582 => x"FF",
		131606 => x"FF",
		132630 => x"FF",
		133654 => x"FF",
		134678 => x"FF",
		135702 => x"FF",
		136726 => x"FF",
		137750 => x"FF",
		138774 => x"FF",
		139798 => x"FF",
		140822 => x"FF",
		141846 => x"FF",
		142870 => x"FF",
		143894 => x"FF",
		144918 => x"FF",
		145942 => x"FF",
		146966 => x"FF",
		147990 => x"FF",
		149014 => x"FF",
		150038 => x"FF",
		151062 => x"FF",
		152086 => x"FF",
		153110 => x"FF",
		154134 => x"FF",
		155158 => x"FF",
		156182 => x"FF",
		157206 => x"FF",
		158230 => x"FF",
		159254 => x"FF",
		160278 => x"FF",
		161302 => x"FF",
		162326 => x"FF",
		163350 => x"FF",
		164374 => x"FF",
		165398 => x"FF",
		166422 => x"FF",
		167446 => x"FF",
		168470 => x"FF",
		169494 => x"FF",
		170518 => x"FF",
		171542 => x"FF",
		172566 => x"FF",
		173590 => x"FF",
		174614 => x"FF",
		175638 => x"FF",
		176662 => x"FF",
		177686 => x"FF",
		178710 => x"FF",
		179734 => x"FF",
		180758 => x"FF",
		181782 => x"FF",
		182806 => x"FF",
		183830 => x"FF",
		184854 => x"FF",
		185878 => x"FF",
		186902 => x"FF",
		187926 => x"FF",
		188950 => x"FF",
		189974 => x"FF",
		190998 => x"FF",
		192022 => x"FF",
		193046 => x"FF",
		194070 => x"FF",
		195094 => x"FF",
		196118 => x"FF",
		197142 => x"FF",
		198166 => x"FF",
		199190 => x"FF",
		200214 => x"FF",
		201238 => x"FF",
		202262 => x"FF",
		203286 => x"FF",
		204310 => x"FF",
		205334 => x"FF",
		206358 => x"FF",
		207382 => x"FF",
		208406 => x"FF",
		209430 => x"FF",
		210454 => x"FF",
		211478 => x"FF",
		212502 => x"FF",
		213526 => x"FF",
		214550 => x"FF",
		215574 => x"FF",
		216598 => x"FF",
		217622 => x"FF",
		218646 => x"FF",
		219670 => x"FF",
		220694 => x"FF",
		221718 => x"FF",
		222742 => x"FF",
		223766 => x"FF",
		224790 => x"FF",
		225814 => x"FF",
		226838 => x"FF",
		227862 => x"FF",
		228886 => x"FF",
		229910 => x"FF",
		230934 => x"FF",
		231958 => x"FF",
		232982 => x"FF",
		234006 => x"FF",
		235030 => x"FF",
		236054 => x"FF",
		237078 => x"FF",
		238102 => x"FF",
		239126 => x"FF",
		240150 => x"FF",
		241174 => x"FF",
		242198 => x"FF",
		243222 => x"FF",
		244246 => x"FF",
		245270 => x"FF",
		246294 => x"FF",
		247318 => x"FF",
		248342 => x"FF",
		249366 => x"FF",
		250390 => x"FF",
		251414 => x"FF",
		252438 => x"FF",
		253462 => x"FF",
		254486 => x"FF",
		255510 => x"FF",
		256534 => x"FF",
		257558 => x"FF",
		258582 => x"FF",
		259606 => x"FF",
		260630 => x"FF",
		261654 => x"FF",
		262678 => x"FF",
		263702 => x"FF",
		264726 => x"FF",
		265750 => x"FF",
		266774 => x"FF",
		267798 => x"FF",
		268822 => x"FF",
		269846 => x"FF",
		270870 => x"FF",
		271894 => x"FF",
		272918 => x"FF",
		273942 => x"FF",
		274966 => x"FF",
		275990 => x"FF",
		277014 => x"FF",
		278038 => x"FF",
		279062 => x"FF",
		280086 => x"FF",
		281110 => x"FF",
		282134 => x"FF",
		283158 => x"FF",
		284182 => x"FF",
		285206 => x"FF",
		286230 => x"FF",
		287254 => x"FF",
		288278 => x"FF",
		289302 => x"FF",
		290326 => x"FF",
		291350 => x"FF",
		292374 => x"FF",
		293398 => x"FF",
		294422 => x"FF",
		295446 => x"FF",
		296470 => x"FF",
		297494 => x"FF",
		298518 => x"FF",
		299542 => x"FF",
		300566 => x"FF",
		301590 => x"FF",
		302614 => x"FF",
		303638 => x"FF",
		304662 => x"FF",
		305686 => x"FF",
		306710 => x"FF",
		307734 => x"FF",
		308758 => x"FF",
		309782 => x"FF",
		310806 => x"FF",
		311830 => x"FF",
		312854 => x"FF",
		313878 => x"FF",
		314902 => x"FF",
		315926 => x"FF",
		316950 => x"FF",
		317974 => x"FF",
		318998 => x"FF",
		320022 => x"FF",
		321046 => x"FF",
		322070 => x"FF",
		323094 => x"FF",
		324118 => x"FF",
		325142 => x"FF",
		326166 => x"FF",
		327190 => x"FF",
		328214 => x"FF",
		329238 => x"FF",
		330262 => x"FF",
		331286 => x"FF",
		332310 => x"FF",
		333334 => x"FF",
		334358 => x"FF",
		335382 => x"FF",
		336406 => x"FF",
		337430 => x"FF",
		338454 => x"FF",
		339478 => x"FF",
		340502 => x"FF",
		341526 => x"FF",
		342550 => x"FF",
		343574 => x"FF",
		344598 => x"FF",
		345622 => x"FF",
		346646 => x"FF",
		347670 => x"FF",
		348694 => x"FF",
		349718 => x"FF",
		350742 => x"FF",
		351766 => x"FF",
		352790 => x"FF",
		353814 => x"FF",
		354838 => x"FF",
		355862 => x"FF",
		356886 => x"FF",
		357910 => x"FF",
		358934 => x"FF",
		359958 => x"FF",
		360982 => x"FF",
		362006 => x"FF",
		363030 => x"FF",
		364054 => x"FF",
		365078 => x"FF",
		366102 => x"FF",
		367126 => x"FF",
		368150 => x"FF",
		369174 => x"FF",
		370198 => x"FF",
		371222 => x"FF",
		372246 => x"FF",
		373270 => x"FF",
		374294 => x"FF",
		375318 => x"FF",
		376342 => x"FF",
		377366 => x"FF",
		378390 => x"FF",
		379414 => x"FF",
		380438 => x"FF",
		381462 => x"FF",
		382486 => x"FF",
		383510 => x"FF",
		384534 => x"FF",
		385558 => x"FF",
		386582 => x"FF",
		387606 => x"FF",
		388630 => x"FF",
		389654 => x"FF",
		390678 => x"FF",
		391702 => x"FF",
		392726 => x"FF",
		393750 => x"FF",
		394774 => x"FF",
		395798 => x"FF",
		396822 => x"FF",
		397846 => x"FF",
		398870 => x"FF",
		399894 => x"FF",
		400918 => x"FF",
		401942 => x"FF",
		402966 => x"FF",
		403990 => x"FF",
		405014 => x"FF",
		406038 => x"FF",
		407062 => x"FF",
		408086 => x"FF",
		409110 => x"FF",
		410134 => x"FF",
		411158 => x"FF",
		412182 => x"FF",
		413206 => x"FF",
		414230 => x"FF",
		415254 => x"FF",
		416278 => x"FF",
		417302 => x"FF",
		418326 => x"FF",
		419350 => x"FF",
		420374 => x"FF",
		421398 => x"FF",
		422422 => x"FF",
		423446 => x"FF",
		424470 => x"FF",
		425494 => x"FF",
		426518 => x"FF",
		427542 => x"FF",
		428566 => x"FF",
		429590 => x"FF",
		430614 => x"FF",
		431638 => x"FF",
		432662 => x"FF",
		433686 => x"FF",
		434710 => x"FF",
		435734 => x"FF",
		436758 => x"FF",
		437782 => x"FF",
		438806 => x"FF",
		439830 => x"FF",
		440854 => x"FF",
		441878 => x"FF",
		442902 => x"FF",
		443926 => x"FF",
		444950 => x"FF",
		445974 => x"FF",
		446998 => x"FF",
		448022 => x"FF",
		449046 => x"FF",
		450070 => x"FF",
		451094 => x"FF",
		452118 => x"FF",
		453142 => x"FF",
		454166 => x"FF",
		455190 => x"FF",
		456214 => x"FF",
		457238 => x"FF",
		458262 => x"FF",
		459286 => x"FF",
		460310 => x"FF",
		461334 => x"FF",
		462358 => x"FF",
		463382 => x"FF",
		464406 => x"FF",
		465430 => x"FF",
		466454 => x"FF",
		467478 => x"FF",
		468502 => x"FF",
		469526 => x"FF",
		19991 => x"FF",
		21015 => x"FF",
		22039 => x"FF",
		23063 => x"FF",
		24087 => x"FF",
		25111 => x"FF",
		26135 => x"FF",
		27159 => x"FF",
		28183 => x"FF",
		29207 => x"FF",
		30231 => x"FF",
		31255 => x"FF",
		32279 => x"FF",
		33303 => x"FF",
		34327 => x"FF",
		35351 => x"FF",
		36375 => x"FF",
		37399 => x"FF",
		38423 => x"FF",
		39447 => x"FF",
		40471 => x"FF",
		41495 => x"FF",
		42519 => x"FF",
		43543 => x"FF",
		44567 => x"FF",
		45591 => x"FF",
		46615 => x"FF",
		47639 => x"FF",
		48663 => x"FF",
		49687 => x"FF",
		50711 => x"FF",
		51735 => x"FF",
		52759 => x"FF",
		53783 => x"FF",
		54807 => x"FF",
		55831 => x"FF",
		56855 => x"FF",
		57879 => x"FF",
		58903 => x"FF",
		59927 => x"FF",
		60951 => x"FF",
		61975 => x"FF",
		62999 => x"FF",
		64023 => x"FF",
		65047 => x"FF",
		66071 => x"FF",
		67095 => x"FF",
		68119 => x"FF",
		69143 => x"FF",
		70167 => x"FF",
		71191 => x"FF",
		72215 => x"FF",
		73239 => x"FF",
		74263 => x"FF",
		75287 => x"FF",
		76311 => x"FF",
		77335 => x"FF",
		78359 => x"FF",
		79383 => x"FF",
		80407 => x"FF",
		81431 => x"FF",
		82455 => x"FF",
		83479 => x"FF",
		84503 => x"FF",
		85527 => x"FF",
		86551 => x"FF",
		87575 => x"FF",
		88599 => x"FF",
		89623 => x"FF",
		90647 => x"FF",
		91671 => x"FF",
		92695 => x"FF",
		93719 => x"FF",
		94743 => x"FF",
		95767 => x"FF",
		96791 => x"FF",
		97815 => x"FF",
		98839 => x"FF",
		99863 => x"FF",
		100887 => x"FF",
		101911 => x"FF",
		102935 => x"FF",
		103959 => x"FF",
		104983 => x"FF",
		106007 => x"FF",
		107031 => x"FF",
		108055 => x"FF",
		109079 => x"FF",
		110103 => x"FF",
		111127 => x"FF",
		112151 => x"FF",
		113175 => x"FF",
		114199 => x"FF",
		115223 => x"FF",
		116247 => x"FF",
		117271 => x"FF",
		118295 => x"FF",
		119319 => x"FF",
		120343 => x"FF",
		121367 => x"FF",
		122391 => x"FF",
		123415 => x"FF",
		124439 => x"FF",
		125463 => x"FF",
		126487 => x"FF",
		127511 => x"FF",
		128535 => x"FF",
		129559 => x"FF",
		130583 => x"FF",
		131607 => x"FF",
		132631 => x"FF",
		133655 => x"FF",
		134679 => x"FF",
		135703 => x"FF",
		136727 => x"FF",
		137751 => x"FF",
		138775 => x"FF",
		139799 => x"FF",
		140823 => x"FF",
		141847 => x"FF",
		142871 => x"FF",
		143895 => x"FF",
		144919 => x"FF",
		145943 => x"FF",
		146967 => x"FF",
		147991 => x"FF",
		149015 => x"FF",
		150039 => x"FF",
		151063 => x"FF",
		152087 => x"FF",
		153111 => x"FF",
		154135 => x"FF",
		155159 => x"FF",
		156183 => x"FF",
		157207 => x"FF",
		158231 => x"FF",
		159255 => x"FF",
		160279 => x"FF",
		161303 => x"FF",
		162327 => x"FF",
		163351 => x"FF",
		164375 => x"FF",
		165399 => x"FF",
		166423 => x"FF",
		167447 => x"FF",
		168471 => x"FF",
		169495 => x"FF",
		170519 => x"FF",
		171543 => x"FF",
		172567 => x"FF",
		173591 => x"FF",
		174615 => x"FF",
		175639 => x"FF",
		176663 => x"FF",
		177687 => x"FF",
		178711 => x"FF",
		179735 => x"FF",
		180759 => x"FF",
		181783 => x"FF",
		182807 => x"FF",
		183831 => x"FF",
		184855 => x"FF",
		185879 => x"FF",
		186903 => x"FF",
		187927 => x"FF",
		188951 => x"FF",
		189975 => x"FF",
		190999 => x"FF",
		192023 => x"FF",
		193047 => x"FF",
		194071 => x"FF",
		195095 => x"FF",
		196119 => x"FF",
		197143 => x"FF",
		198167 => x"FF",
		199191 => x"FF",
		200215 => x"FF",
		201239 => x"FF",
		202263 => x"FF",
		203287 => x"FF",
		204311 => x"FF",
		205335 => x"FF",
		206359 => x"FF",
		207383 => x"FF",
		208407 => x"FF",
		209431 => x"FF",
		210455 => x"FF",
		211479 => x"FF",
		212503 => x"FF",
		213527 => x"FF",
		214551 => x"FF",
		215575 => x"FF",
		216599 => x"FF",
		217623 => x"FF",
		218647 => x"FF",
		219671 => x"FF",
		220695 => x"FF",
		221719 => x"FF",
		222743 => x"FF",
		223767 => x"FF",
		224791 => x"FF",
		225815 => x"FF",
		226839 => x"FF",
		227863 => x"FF",
		228887 => x"FF",
		229911 => x"FF",
		230935 => x"FF",
		231959 => x"FF",
		232983 => x"FF",
		234007 => x"FF",
		235031 => x"FF",
		236055 => x"FF",
		237079 => x"FF",
		238103 => x"FF",
		239127 => x"FF",
		240151 => x"FF",
		241175 => x"FF",
		242199 => x"FF",
		243223 => x"FF",
		244247 => x"FF",
		245271 => x"FF",
		246295 => x"FF",
		247319 => x"FF",
		248343 => x"FF",
		249367 => x"FF",
		250391 => x"FF",
		251415 => x"FF",
		252439 => x"FF",
		253463 => x"FF",
		254487 => x"FF",
		255511 => x"FF",
		256535 => x"FF",
		257559 => x"FF",
		258583 => x"FF",
		259607 => x"FF",
		260631 => x"FF",
		261655 => x"FF",
		262679 => x"FF",
		263703 => x"FF",
		264727 => x"FF",
		265751 => x"FF",
		266775 => x"FF",
		267799 => x"FF",
		268823 => x"FF",
		269847 => x"FF",
		270871 => x"FF",
		271895 => x"FF",
		272919 => x"FF",
		273943 => x"FF",
		274967 => x"FF",
		275991 => x"FF",
		277015 => x"FF",
		278039 => x"FF",
		279063 => x"FF",
		280087 => x"FF",
		281111 => x"FF",
		282135 => x"FF",
		283159 => x"FF",
		284183 => x"FF",
		285207 => x"FF",
		286231 => x"FF",
		287255 => x"FF",
		288279 => x"FF",
		289303 => x"FF",
		290327 => x"FF",
		291351 => x"FF",
		292375 => x"FF",
		293399 => x"FF",
		294423 => x"FF",
		295447 => x"FF",
		296471 => x"FF",
		297495 => x"FF",
		298519 => x"FF",
		299543 => x"FF",
		300567 => x"FF",
		301591 => x"FF",
		302615 => x"FF",
		303639 => x"FF",
		304663 => x"FF",
		305687 => x"FF",
		306711 => x"FF",
		307735 => x"FF",
		308759 => x"FF",
		309783 => x"FF",
		310807 => x"FF",
		311831 => x"FF",
		312855 => x"FF",
		313879 => x"FF",
		314903 => x"FF",
		315927 => x"FF",
		316951 => x"FF",
		317975 => x"FF",
		318999 => x"FF",
		320023 => x"FF",
		321047 => x"FF",
		322071 => x"FF",
		323095 => x"FF",
		324119 => x"FF",
		325143 => x"FF",
		326167 => x"FF",
		327191 => x"FF",
		328215 => x"FF",
		329239 => x"FF",
		330263 => x"FF",
		331287 => x"FF",
		332311 => x"FF",
		333335 => x"FF",
		334359 => x"FF",
		335383 => x"FF",
		336407 => x"FF",
		337431 => x"FF",
		338455 => x"FF",
		339479 => x"FF",
		340503 => x"FF",
		341527 => x"FF",
		342551 => x"FF",
		343575 => x"FF",
		344599 => x"FF",
		345623 => x"FF",
		346647 => x"FF",
		347671 => x"FF",
		348695 => x"FF",
		349719 => x"FF",
		350743 => x"FF",
		351767 => x"FF",
		352791 => x"FF",
		353815 => x"FF",
		354839 => x"FF",
		355863 => x"FF",
		356887 => x"FF",
		357911 => x"FF",
		358935 => x"FF",
		359959 => x"FF",
		360983 => x"FF",
		362007 => x"FF",
		363031 => x"FF",
		364055 => x"FF",
		365079 => x"FF",
		366103 => x"FF",
		367127 => x"FF",
		368151 => x"FF",
		369175 => x"FF",
		370199 => x"FF",
		371223 => x"FF",
		372247 => x"FF",
		373271 => x"FF",
		374295 => x"FF",
		375319 => x"FF",
		376343 => x"FF",
		377367 => x"FF",
		378391 => x"FF",
		379415 => x"FF",
		380439 => x"FF",
		381463 => x"FF",
		382487 => x"FF",
		383511 => x"FF",
		384535 => x"FF",
		385559 => x"FF",
		386583 => x"FF",
		387607 => x"FF",
		388631 => x"FF",
		389655 => x"FF",
		390679 => x"FF",
		391703 => x"FF",
		392727 => x"FF",
		393751 => x"FF",
		394775 => x"FF",
		395799 => x"FF",
		396823 => x"FF",
		397847 => x"FF",
		398871 => x"FF",
		399895 => x"FF",
		400919 => x"FF",
		401943 => x"FF",
		402967 => x"FF",
		403991 => x"FF",
		405015 => x"FF",
		406039 => x"FF",
		407063 => x"FF",
		408087 => x"FF",
		409111 => x"FF",
		410135 => x"FF",
		411159 => x"FF",
		412183 => x"FF",
		413207 => x"FF",
		414231 => x"FF",
		415255 => x"FF",
		416279 => x"FF",
		417303 => x"FF",
		418327 => x"FF",
		419351 => x"FF",
		420375 => x"FF",
		421399 => x"FF",
		422423 => x"FF",
		423447 => x"FF",
		424471 => x"FF",
		425495 => x"FF",
		426519 => x"FF",
		427543 => x"FF",
		428567 => x"FF",
		429591 => x"FF",
		430615 => x"FF",
		431639 => x"FF",
		432663 => x"FF",
		433687 => x"FF",
		434711 => x"FF",
		435735 => x"FF",
		436759 => x"FF",
		437783 => x"FF",
		438807 => x"FF",
		439831 => x"FF",
		440855 => x"FF",
		441879 => x"FF",
		442903 => x"FF",
		443927 => x"FF",
		444951 => x"FF",
		445975 => x"FF",
		446999 => x"FF",
		448023 => x"FF",
		449047 => x"FF",
		450071 => x"FF",
		451095 => x"FF",
		452119 => x"FF",
		453143 => x"FF",
		454167 => x"FF",
		455191 => x"FF",
		456215 => x"FF",
		457239 => x"FF",
		458263 => x"FF",
		459287 => x"FF",
		460311 => x"FF",
		461335 => x"FF",
		462359 => x"FF",
		463383 => x"FF",
		464407 => x"FF",
		465431 => x"FF",
		466455 => x"FF",
		467479 => x"FF",
		468503 => x"FF",
		469527 => x"FF",
		19992 => x"FF",
		21016 => x"FF",
		22040 => x"FF",
		23064 => x"FF",
		24088 => x"FF",
		25112 => x"FF",
		26136 => x"FF",
		27160 => x"FF",
		28184 => x"FF",
		29208 => x"FF",
		30232 => x"FF",
		31256 => x"FF",
		32280 => x"FF",
		33304 => x"FF",
		34328 => x"FF",
		35352 => x"FF",
		36376 => x"FF",
		37400 => x"FF",
		38424 => x"FF",
		39448 => x"FF",
		40472 => x"FF",
		41496 => x"FF",
		42520 => x"FF",
		43544 => x"FF",
		44568 => x"FF",
		45592 => x"FF",
		46616 => x"FF",
		47640 => x"FF",
		48664 => x"FF",
		49688 => x"FF",
		50712 => x"FF",
		51736 => x"FF",
		52760 => x"FF",
		53784 => x"FF",
		54808 => x"FF",
		55832 => x"FF",
		56856 => x"FF",
		57880 => x"FF",
		58904 => x"FF",
		59928 => x"FF",
		60952 => x"FF",
		61976 => x"FF",
		63000 => x"FF",
		64024 => x"FF",
		65048 => x"FF",
		66072 => x"FF",
		67096 => x"FF",
		68120 => x"FF",
		69144 => x"FF",
		70168 => x"FF",
		71192 => x"FF",
		72216 => x"FF",
		73240 => x"FF",
		74264 => x"FF",
		75288 => x"FF",
		76312 => x"FF",
		77336 => x"FF",
		78360 => x"FF",
		79384 => x"FF",
		80408 => x"FF",
		81432 => x"FF",
		82456 => x"FF",
		83480 => x"FF",
		84504 => x"FF",
		85528 => x"FF",
		86552 => x"FF",
		87576 => x"FF",
		88600 => x"FF",
		89624 => x"FF",
		90648 => x"FF",
		91672 => x"FF",
		92696 => x"FF",
		93720 => x"FF",
		94744 => x"FF",
		95768 => x"FF",
		96792 => x"FF",
		97816 => x"FF",
		98840 => x"FF",
		99864 => x"FF",
		100888 => x"FF",
		101912 => x"FF",
		102936 => x"FF",
		103960 => x"FF",
		104984 => x"FF",
		106008 => x"FF",
		107032 => x"FF",
		108056 => x"FF",
		109080 => x"FF",
		110104 => x"FF",
		111128 => x"FF",
		112152 => x"FF",
		113176 => x"FF",
		114200 => x"FF",
		115224 => x"FF",
		116248 => x"FF",
		117272 => x"FF",
		118296 => x"FF",
		119320 => x"FF",
		120344 => x"FF",
		121368 => x"FF",
		122392 => x"FF",
		123416 => x"FF",
		124440 => x"FF",
		125464 => x"FF",
		126488 => x"FF",
		127512 => x"FF",
		128536 => x"FF",
		129560 => x"FF",
		130584 => x"FF",
		131608 => x"FF",
		132632 => x"FF",
		133656 => x"FF",
		134680 => x"FF",
		135704 => x"FF",
		136728 => x"FF",
		137752 => x"FF",
		138776 => x"FF",
		139800 => x"FF",
		140824 => x"FF",
		141848 => x"FF",
		142872 => x"FF",
		143896 => x"FF",
		144920 => x"FF",
		145944 => x"FF",
		146968 => x"FF",
		147992 => x"FF",
		149016 => x"FF",
		150040 => x"FF",
		151064 => x"FF",
		152088 => x"FF",
		153112 => x"FF",
		154136 => x"FF",
		155160 => x"FF",
		156184 => x"FF",
		157208 => x"FF",
		158232 => x"FF",
		159256 => x"FF",
		160280 => x"FF",
		161304 => x"FF",
		162328 => x"FF",
		163352 => x"FF",
		164376 => x"FF",
		165400 => x"FF",
		166424 => x"FF",
		167448 => x"FF",
		168472 => x"FF",
		169496 => x"FF",
		170520 => x"FF",
		171544 => x"FF",
		172568 => x"FF",
		173592 => x"FF",
		174616 => x"FF",
		175640 => x"FF",
		176664 => x"FF",
		177688 => x"FF",
		178712 => x"FF",
		179736 => x"FF",
		180760 => x"FF",
		181784 => x"FF",
		182808 => x"FF",
		183832 => x"FF",
		184856 => x"FF",
		185880 => x"FF",
		186904 => x"FF",
		187928 => x"FF",
		188952 => x"FF",
		189976 => x"FF",
		191000 => x"FF",
		192024 => x"FF",
		193048 => x"FF",
		194072 => x"FF",
		195096 => x"FF",
		196120 => x"FF",
		197144 => x"FF",
		198168 => x"FF",
		199192 => x"FF",
		200216 => x"FF",
		201240 => x"FF",
		202264 => x"FF",
		203288 => x"FF",
		204312 => x"FF",
		205336 => x"FF",
		206360 => x"FF",
		207384 => x"FF",
		208408 => x"FF",
		209432 => x"FF",
		210456 => x"FF",
		211480 => x"FF",
		212504 => x"FF",
		213528 => x"FF",
		214552 => x"FF",
		215576 => x"FF",
		216600 => x"FF",
		217624 => x"FF",
		218648 => x"FF",
		219672 => x"FF",
		220696 => x"FF",
		221720 => x"FF",
		222744 => x"FF",
		223768 => x"FF",
		224792 => x"FF",
		225816 => x"FF",
		226840 => x"FF",
		227864 => x"FF",
		228888 => x"FF",
		229912 => x"FF",
		230936 => x"FF",
		231960 => x"FF",
		232984 => x"FF",
		234008 => x"FF",
		235032 => x"FF",
		236056 => x"FF",
		237080 => x"FF",
		238104 => x"FF",
		239128 => x"FF",
		240152 => x"FF",
		241176 => x"FF",
		242200 => x"FF",
		243224 => x"FF",
		244248 => x"FF",
		245272 => x"FF",
		246296 => x"FF",
		247320 => x"FF",
		248344 => x"FF",
		249368 => x"FF",
		250392 => x"FF",
		251416 => x"FF",
		252440 => x"FF",
		253464 => x"FF",
		254488 => x"FF",
		255512 => x"FF",
		256536 => x"FF",
		257560 => x"FF",
		258584 => x"FF",
		259608 => x"FF",
		260632 => x"FF",
		261656 => x"FF",
		262680 => x"FF",
		263704 => x"FF",
		264728 => x"FF",
		265752 => x"FF",
		266776 => x"FF",
		267800 => x"FF",
		268824 => x"FF",
		269848 => x"FF",
		270872 => x"FF",
		271896 => x"FF",
		272920 => x"FF",
		273944 => x"FF",
		274968 => x"FF",
		275992 => x"FF",
		277016 => x"FF",
		278040 => x"FF",
		279064 => x"FF",
		280088 => x"FF",
		281112 => x"FF",
		282136 => x"FF",
		283160 => x"FF",
		284184 => x"FF",
		285208 => x"FF",
		286232 => x"FF",
		287256 => x"FF",
		288280 => x"FF",
		289304 => x"FF",
		290328 => x"FF",
		291352 => x"FF",
		292376 => x"FF",
		293400 => x"FF",
		294424 => x"FF",
		295448 => x"FF",
		296472 => x"FF",
		297496 => x"FF",
		298520 => x"FF",
		299544 => x"FF",
		300568 => x"FF",
		301592 => x"FF",
		302616 => x"FF",
		303640 => x"FF",
		304664 => x"FF",
		305688 => x"FF",
		306712 => x"FF",
		307736 => x"FF",
		308760 => x"FF",
		309784 => x"FF",
		310808 => x"FF",
		311832 => x"FF",
		312856 => x"FF",
		313880 => x"FF",
		314904 => x"FF",
		315928 => x"FF",
		316952 => x"FF",
		317976 => x"FF",
		319000 => x"FF",
		320024 => x"FF",
		321048 => x"FF",
		322072 => x"FF",
		323096 => x"FF",
		324120 => x"FF",
		325144 => x"FF",
		326168 => x"FF",
		327192 => x"FF",
		328216 => x"FF",
		329240 => x"FF",
		330264 => x"FF",
		331288 => x"FF",
		332312 => x"FF",
		333336 => x"FF",
		334360 => x"FF",
		335384 => x"FF",
		336408 => x"FF",
		337432 => x"FF",
		338456 => x"FF",
		339480 => x"FF",
		340504 => x"FF",
		341528 => x"FF",
		342552 => x"FF",
		343576 => x"FF",
		344600 => x"FF",
		345624 => x"FF",
		346648 => x"FF",
		347672 => x"FF",
		348696 => x"FF",
		349720 => x"FF",
		350744 => x"FF",
		351768 => x"FF",
		352792 => x"FF",
		353816 => x"FF",
		354840 => x"FF",
		355864 => x"FF",
		356888 => x"FF",
		357912 => x"FF",
		358936 => x"FF",
		359960 => x"FF",
		360984 => x"FF",
		362008 => x"FF",
		363032 => x"FF",
		364056 => x"FF",
		365080 => x"FF",
		366104 => x"FF",
		367128 => x"FF",
		368152 => x"FF",
		369176 => x"FF",
		370200 => x"FF",
		371224 => x"FF",
		372248 => x"FF",
		373272 => x"FF",
		374296 => x"FF",
		375320 => x"FF",
		376344 => x"FF",
		377368 => x"FF",
		378392 => x"FF",
		379416 => x"FF",
		380440 => x"FF",
		381464 => x"FF",
		382488 => x"FF",
		383512 => x"FF",
		384536 => x"FF",
		385560 => x"FF",
		386584 => x"FF",
		387608 => x"FF",
		388632 => x"FF",
		389656 => x"FF",
		390680 => x"FF",
		391704 => x"FF",
		392728 => x"FF",
		393752 => x"FF",
		394776 => x"FF",
		395800 => x"FF",
		396824 => x"FF",
		397848 => x"FF",
		398872 => x"FF",
		399896 => x"FF",
		400920 => x"FF",
		401944 => x"FF",
		402968 => x"FF",
		403992 => x"FF",
		405016 => x"FF",
		406040 => x"FF",
		407064 => x"FF",
		408088 => x"FF",
		409112 => x"FF",
		410136 => x"FF",
		411160 => x"FF",
		412184 => x"FF",
		413208 => x"FF",
		414232 => x"FF",
		415256 => x"FF",
		416280 => x"FF",
		417304 => x"FF",
		418328 => x"FF",
		419352 => x"FF",
		420376 => x"FF",
		421400 => x"FF",
		422424 => x"FF",
		423448 => x"FF",
		424472 => x"FF",
		425496 => x"FF",
		426520 => x"FF",
		427544 => x"FF",
		428568 => x"FF",
		429592 => x"FF",
		430616 => x"FF",
		431640 => x"FF",
		432664 => x"FF",
		433688 => x"FF",
		434712 => x"FF",
		435736 => x"FF",
		436760 => x"FF",
		437784 => x"FF",
		438808 => x"FF",
		439832 => x"FF",
		440856 => x"FF",
		441880 => x"FF",
		442904 => x"FF",
		443928 => x"FF",
		444952 => x"FF",
		445976 => x"FF",
		447000 => x"FF",
		448024 => x"FF",
		449048 => x"FF",
		450072 => x"FF",
		451096 => x"FF",
		452120 => x"FF",
		453144 => x"FF",
		454168 => x"FF",
		455192 => x"FF",
		456216 => x"FF",
		457240 => x"FF",
		458264 => x"FF",
		459288 => x"FF",
		460312 => x"FF",
		461336 => x"FF",
		462360 => x"FF",
		463384 => x"FF",
		464408 => x"FF",
		465432 => x"FF",
		466456 => x"FF",
		467480 => x"FF",
		468504 => x"FF",
		469528 => x"FF",
		19993 => x"FF",
		21017 => x"FF",
		22041 => x"FF",
		23065 => x"FF",
		24089 => x"FF",
		25113 => x"FF",
		26137 => x"FF",
		27161 => x"FF",
		28185 => x"FF",
		29209 => x"FF",
		30233 => x"FF",
		31257 => x"FF",
		32281 => x"FF",
		33305 => x"FF",
		34329 => x"FF",
		35353 => x"FF",
		36377 => x"FF",
		37401 => x"FF",
		38425 => x"FF",
		39449 => x"FF",
		40473 => x"FF",
		41497 => x"FF",
		42521 => x"FF",
		43545 => x"FF",
		44569 => x"FF",
		45593 => x"FF",
		46617 => x"FF",
		47641 => x"FF",
		48665 => x"FF",
		49689 => x"FF",
		50713 => x"FF",
		51737 => x"FF",
		52761 => x"FF",
		53785 => x"FF",
		54809 => x"FF",
		55833 => x"FF",
		56857 => x"FF",
		57881 => x"FF",
		58905 => x"FF",
		59929 => x"FF",
		60953 => x"FF",
		61977 => x"FF",
		63001 => x"FF",
		64025 => x"FF",
		65049 => x"FF",
		66073 => x"FF",
		67097 => x"FF",
		68121 => x"FF",
		69145 => x"FF",
		70169 => x"FF",
		71193 => x"FF",
		72217 => x"FF",
		73241 => x"FF",
		74265 => x"FF",
		75289 => x"FF",
		76313 => x"FF",
		77337 => x"FF",
		78361 => x"FF",
		79385 => x"FF",
		80409 => x"FF",
		81433 => x"FF",
		82457 => x"FF",
		83481 => x"FF",
		84505 => x"FF",
		85529 => x"FF",
		86553 => x"FF",
		87577 => x"FF",
		88601 => x"FF",
		89625 => x"FF",
		90649 => x"FF",
		91673 => x"FF",
		92697 => x"FF",
		93721 => x"FF",
		94745 => x"FF",
		95769 => x"FF",
		96793 => x"FF",
		97817 => x"FF",
		98841 => x"FF",
		99865 => x"FF",
		100889 => x"FF",
		101913 => x"FF",
		102937 => x"FF",
		103961 => x"FF",
		104985 => x"FF",
		106009 => x"FF",
		107033 => x"FF",
		108057 => x"FF",
		109081 => x"FF",
		110105 => x"FF",
		111129 => x"FF",
		112153 => x"FF",
		113177 => x"FF",
		114201 => x"FF",
		115225 => x"FF",
		116249 => x"FF",
		117273 => x"FF",
		118297 => x"FF",
		119321 => x"FF",
		120345 => x"FF",
		121369 => x"FF",
		122393 => x"FF",
		123417 => x"FF",
		124441 => x"FF",
		125465 => x"FF",
		126489 => x"FF",
		127513 => x"FF",
		128537 => x"FF",
		129561 => x"FF",
		130585 => x"FF",
		131609 => x"FF",
		132633 => x"FF",
		133657 => x"FF",
		134681 => x"FF",
		135705 => x"FF",
		136729 => x"FF",
		137753 => x"FF",
		138777 => x"FF",
		139801 => x"FF",
		140825 => x"FF",
		141849 => x"FF",
		142873 => x"FF",
		143897 => x"FF",
		144921 => x"FF",
		145945 => x"FF",
		146969 => x"FF",
		147993 => x"FF",
		149017 => x"FF",
		150041 => x"FF",
		151065 => x"FF",
		152089 => x"FF",
		153113 => x"FF",
		154137 => x"FF",
		155161 => x"FF",
		156185 => x"FF",
		157209 => x"FF",
		158233 => x"FF",
		159257 => x"FF",
		160281 => x"FF",
		161305 => x"FF",
		162329 => x"FF",
		163353 => x"FF",
		164377 => x"FF",
		165401 => x"FF",
		166425 => x"FF",
		167449 => x"FF",
		168473 => x"FF",
		169497 => x"FF",
		170521 => x"FF",
		171545 => x"FF",
		172569 => x"FF",
		173593 => x"FF",
		174617 => x"FF",
		175641 => x"FF",
		176665 => x"FF",
		177689 => x"FF",
		178713 => x"FF",
		179737 => x"FF",
		180761 => x"FF",
		181785 => x"FF",
		182809 => x"FF",
		183833 => x"FF",
		184857 => x"FF",
		185881 => x"FF",
		186905 => x"FF",
		187929 => x"FF",
		188953 => x"FF",
		189977 => x"FF",
		191001 => x"FF",
		192025 => x"FF",
		193049 => x"FF",
		194073 => x"FF",
		195097 => x"FF",
		196121 => x"FF",
		197145 => x"FF",
		198169 => x"FF",
		199193 => x"FF",
		200217 => x"FF",
		201241 => x"FF",
		202265 => x"FF",
		203289 => x"FF",
		204313 => x"FF",
		205337 => x"FF",
		206361 => x"FF",
		207385 => x"FF",
		208409 => x"FF",
		209433 => x"FF",
		210457 => x"FF",
		211481 => x"FF",
		212505 => x"FF",
		213529 => x"FF",
		214553 => x"FF",
		215577 => x"FF",
		216601 => x"FF",
		217625 => x"FF",
		218649 => x"FF",
		219673 => x"FF",
		220697 => x"FF",
		221721 => x"FF",
		222745 => x"FF",
		223769 => x"FF",
		224793 => x"FF",
		225817 => x"FF",
		226841 => x"FF",
		227865 => x"FF",
		228889 => x"FF",
		229913 => x"FF",
		230937 => x"FF",
		231961 => x"FF",
		232985 => x"FF",
		234009 => x"FF",
		235033 => x"FF",
		236057 => x"FF",
		237081 => x"FF",
		238105 => x"FF",
		239129 => x"FF",
		240153 => x"FF",
		241177 => x"FF",
		242201 => x"FF",
		243225 => x"FF",
		244249 => x"FF",
		245273 => x"FF",
		246297 => x"FF",
		247321 => x"FF",
		248345 => x"FF",
		249369 => x"FF",
		250393 => x"FF",
		251417 => x"FF",
		252441 => x"FF",
		253465 => x"FF",
		254489 => x"FF",
		255513 => x"FF",
		256537 => x"FF",
		257561 => x"FF",
		258585 => x"FF",
		259609 => x"FF",
		260633 => x"FF",
		261657 => x"FF",
		262681 => x"FF",
		263705 => x"FF",
		264729 => x"FF",
		265753 => x"FF",
		266777 => x"FF",
		267801 => x"FF",
		268825 => x"FF",
		269849 => x"FF",
		270873 => x"FF",
		271897 => x"FF",
		272921 => x"FF",
		273945 => x"FF",
		274969 => x"FF",
		275993 => x"FF",
		277017 => x"FF",
		278041 => x"FF",
		279065 => x"FF",
		280089 => x"FF",
		281113 => x"FF",
		282137 => x"FF",
		283161 => x"FF",
		284185 => x"FF",
		285209 => x"FF",
		286233 => x"FF",
		287257 => x"FF",
		288281 => x"FF",
		289305 => x"FF",
		290329 => x"FF",
		291353 => x"FF",
		292377 => x"FF",
		293401 => x"FF",
		294425 => x"FF",
		295449 => x"FF",
		296473 => x"FF",
		297497 => x"FF",
		298521 => x"FF",
		299545 => x"FF",
		300569 => x"FF",
		301593 => x"FF",
		302617 => x"FF",
		303641 => x"FF",
		304665 => x"FF",
		305689 => x"FF",
		306713 => x"FF",
		307737 => x"FF",
		308761 => x"FF",
		309785 => x"FF",
		310809 => x"FF",
		311833 => x"FF",
		312857 => x"FF",
		313881 => x"FF",
		314905 => x"FF",
		315929 => x"FF",
		316953 => x"FF",
		317977 => x"FF",
		319001 => x"FF",
		320025 => x"FF",
		321049 => x"FF",
		322073 => x"FF",
		323097 => x"FF",
		324121 => x"FF",
		325145 => x"FF",
		326169 => x"FF",
		327193 => x"FF",
		328217 => x"FF",
		329241 => x"FF",
		330265 => x"FF",
		331289 => x"FF",
		332313 => x"FF",
		333337 => x"FF",
		334361 => x"FF",
		335385 => x"FF",
		336409 => x"FF",
		337433 => x"FF",
		338457 => x"FF",
		339481 => x"FF",
		340505 => x"FF",
		341529 => x"FF",
		342553 => x"FF",
		343577 => x"FF",
		344601 => x"FF",
		345625 => x"FF",
		346649 => x"FF",
		347673 => x"FF",
		348697 => x"FF",
		349721 => x"FF",
		350745 => x"FF",
		351769 => x"FF",
		352793 => x"FF",
		353817 => x"FF",
		354841 => x"FF",
		355865 => x"FF",
		356889 => x"FF",
		357913 => x"FF",
		358937 => x"FF",
		359961 => x"FF",
		360985 => x"FF",
		362009 => x"FF",
		363033 => x"FF",
		364057 => x"FF",
		365081 => x"FF",
		366105 => x"FF",
		367129 => x"FF",
		368153 => x"FF",
		369177 => x"FF",
		370201 => x"FF",
		371225 => x"FF",
		372249 => x"FF",
		373273 => x"FF",
		374297 => x"FF",
		375321 => x"FF",
		376345 => x"FF",
		377369 => x"FF",
		378393 => x"FF",
		379417 => x"FF",
		380441 => x"FF",
		381465 => x"FF",
		382489 => x"FF",
		383513 => x"FF",
		384537 => x"FF",
		385561 => x"FF",
		386585 => x"FF",
		387609 => x"FF",
		388633 => x"FF",
		389657 => x"FF",
		390681 => x"FF",
		391705 => x"FF",
		392729 => x"FF",
		393753 => x"FF",
		394777 => x"FF",
		395801 => x"FF",
		396825 => x"FF",
		397849 => x"FF",
		398873 => x"FF",
		399897 => x"FF",
		400921 => x"FF",
		401945 => x"FF",
		402969 => x"FF",
		403993 => x"FF",
		405017 => x"FF",
		406041 => x"FF",
		407065 => x"FF",
		408089 => x"FF",
		409113 => x"FF",
		410137 => x"FF",
		411161 => x"FF",
		412185 => x"FF",
		413209 => x"FF",
		414233 => x"FF",
		415257 => x"FF",
		416281 => x"FF",
		417305 => x"FF",
		418329 => x"FF",
		419353 => x"FF",
		420377 => x"FF",
		421401 => x"FF",
		422425 => x"FF",
		423449 => x"FF",
		424473 => x"FF",
		425497 => x"FF",
		426521 => x"FF",
		427545 => x"FF",
		428569 => x"FF",
		429593 => x"FF",
		430617 => x"FF",
		431641 => x"FF",
		432665 => x"FF",
		433689 => x"FF",
		434713 => x"FF",
		435737 => x"FF",
		436761 => x"FF",
		437785 => x"FF",
		438809 => x"FF",
		439833 => x"FF",
		440857 => x"FF",
		441881 => x"FF",
		442905 => x"FF",
		443929 => x"FF",
		444953 => x"FF",
		445977 => x"FF",
		447001 => x"FF",
		448025 => x"FF",
		449049 => x"FF",
		450073 => x"FF",
		451097 => x"FF",
		452121 => x"FF",
		453145 => x"FF",
		454169 => x"FF",
		455193 => x"FF",
		456217 => x"FF",
		457241 => x"FF",
		458265 => x"FF",
		459289 => x"FF",
		460313 => x"FF",
		461337 => x"FF",
		462361 => x"FF",
		463385 => x"FF",
		464409 => x"FF",
		465433 => x"FF",
		466457 => x"FF",
		467481 => x"FF",
		468505 => x"FF",
		469529 => x"FF",
		19994 => x"FF",
		21018 => x"FF",
		22042 => x"FF",
		23066 => x"FF",
		24090 => x"FF",
		25114 => x"FF",
		26138 => x"FF",
		27162 => x"FF",
		28186 => x"FF",
		29210 => x"FF",
		30234 => x"FF",
		31258 => x"FF",
		32282 => x"FF",
		33306 => x"FF",
		34330 => x"FF",
		35354 => x"FF",
		36378 => x"FF",
		37402 => x"FF",
		38426 => x"FF",
		39450 => x"FF",
		40474 => x"FF",
		41498 => x"FF",
		42522 => x"FF",
		43546 => x"FF",
		44570 => x"FF",
		45594 => x"FF",
		46618 => x"FF",
		47642 => x"FF",
		48666 => x"FF",
		49690 => x"FF",
		50714 => x"FF",
		51738 => x"FF",
		52762 => x"FF",
		53786 => x"FF",
		54810 => x"FF",
		55834 => x"FF",
		56858 => x"FF",
		57882 => x"FF",
		58906 => x"FF",
		59930 => x"FF",
		60954 => x"FF",
		61978 => x"FF",
		63002 => x"FF",
		64026 => x"FF",
		65050 => x"FF",
		66074 => x"FF",
		67098 => x"FF",
		68122 => x"FF",
		69146 => x"FF",
		70170 => x"FF",
		71194 => x"FF",
		72218 => x"FF",
		73242 => x"FF",
		74266 => x"FF",
		75290 => x"FF",
		76314 => x"FF",
		77338 => x"FF",
		78362 => x"FF",
		79386 => x"FF",
		80410 => x"FF",
		81434 => x"FF",
		82458 => x"FF",
		83482 => x"FF",
		84506 => x"FF",
		85530 => x"FF",
		86554 => x"FF",
		87578 => x"FF",
		88602 => x"FF",
		89626 => x"FF",
		90650 => x"FF",
		91674 => x"FF",
		92698 => x"FF",
		93722 => x"FF",
		94746 => x"FF",
		95770 => x"FF",
		96794 => x"FF",
		97818 => x"FF",
		98842 => x"FF",
		99866 => x"FF",
		100890 => x"FF",
		101914 => x"FF",
		102938 => x"FF",
		103962 => x"FF",
		104986 => x"FF",
		106010 => x"FF",
		107034 => x"FF",
		108058 => x"FF",
		109082 => x"FF",
		110106 => x"FF",
		111130 => x"FF",
		112154 => x"FF",
		113178 => x"FF",
		114202 => x"FF",
		115226 => x"FF",
		116250 => x"FF",
		117274 => x"FF",
		118298 => x"FF",
		119322 => x"FF",
		120346 => x"FF",
		121370 => x"FF",
		122394 => x"FF",
		123418 => x"FF",
		124442 => x"FF",
		125466 => x"FF",
		126490 => x"FF",
		127514 => x"FF",
		128538 => x"FF",
		129562 => x"FF",
		130586 => x"FF",
		131610 => x"FF",
		132634 => x"FF",
		133658 => x"FF",
		134682 => x"FF",
		135706 => x"FF",
		136730 => x"FF",
		137754 => x"FF",
		138778 => x"FF",
		139802 => x"FF",
		140826 => x"FF",
		141850 => x"FF",
		142874 => x"FF",
		143898 => x"FF",
		144922 => x"FF",
		145946 => x"FF",
		146970 => x"FF",
		147994 => x"FF",
		149018 => x"FF",
		150042 => x"FF",
		151066 => x"FF",
		152090 => x"FF",
		153114 => x"FF",
		154138 => x"FF",
		155162 => x"FF",
		156186 => x"FF",
		157210 => x"FF",
		158234 => x"FF",
		159258 => x"FF",
		160282 => x"FF",
		161306 => x"FF",
		162330 => x"FF",
		163354 => x"FF",
		164378 => x"FF",
		165402 => x"FF",
		166426 => x"FF",
		167450 => x"FF",
		168474 => x"FF",
		169498 => x"FF",
		170522 => x"FF",
		171546 => x"FF",
		172570 => x"FF",
		173594 => x"FF",
		174618 => x"FF",
		175642 => x"FF",
		176666 => x"FF",
		177690 => x"FF",
		178714 => x"FF",
		179738 => x"FF",
		180762 => x"FF",
		181786 => x"FF",
		182810 => x"FF",
		183834 => x"FF",
		184858 => x"FF",
		185882 => x"FF",
		186906 => x"FF",
		187930 => x"FF",
		188954 => x"FF",
		189978 => x"FF",
		191002 => x"FF",
		192026 => x"FF",
		193050 => x"FF",
		194074 => x"FF",
		195098 => x"FF",
		196122 => x"FF",
		197146 => x"FF",
		198170 => x"FF",
		199194 => x"FF",
		200218 => x"FF",
		201242 => x"FF",
		202266 => x"FF",
		203290 => x"FF",
		204314 => x"FF",
		205338 => x"FF",
		206362 => x"FF",
		207386 => x"FF",
		208410 => x"FF",
		209434 => x"FF",
		210458 => x"FF",
		211482 => x"FF",
		212506 => x"FF",
		213530 => x"FF",
		214554 => x"FF",
		215578 => x"FF",
		216602 => x"FF",
		217626 => x"FF",
		218650 => x"FF",
		219674 => x"FF",
		220698 => x"FF",
		221722 => x"FF",
		222746 => x"FF",
		223770 => x"FF",
		224794 => x"FF",
		225818 => x"FF",
		226842 => x"FF",
		227866 => x"FF",
		228890 => x"FF",
		229914 => x"FF",
		230938 => x"FF",
		231962 => x"FF",
		232986 => x"FF",
		234010 => x"FF",
		235034 => x"FF",
		236058 => x"FF",
		237082 => x"FF",
		238106 => x"FF",
		239130 => x"FF",
		240154 => x"FF",
		241178 => x"FF",
		242202 => x"FF",
		243226 => x"FF",
		244250 => x"FF",
		245274 => x"FF",
		246298 => x"FF",
		247322 => x"FF",
		248346 => x"FF",
		249370 => x"FF",
		250394 => x"FF",
		251418 => x"FF",
		252442 => x"FF",
		253466 => x"FF",
		254490 => x"FF",
		255514 => x"FF",
		256538 => x"FF",
		257562 => x"FF",
		258586 => x"FF",
		259610 => x"FF",
		260634 => x"FF",
		261658 => x"FF",
		262682 => x"FF",
		263706 => x"FF",
		264730 => x"FF",
		265754 => x"FF",
		266778 => x"FF",
		267802 => x"FF",
		268826 => x"FF",
		269850 => x"FF",
		270874 => x"FF",
		271898 => x"FF",
		272922 => x"FF",
		273946 => x"FF",
		274970 => x"FF",
		275994 => x"FF",
		277018 => x"FF",
		278042 => x"FF",
		279066 => x"FF",
		280090 => x"FF",
		281114 => x"FF",
		282138 => x"FF",
		283162 => x"FF",
		284186 => x"FF",
		285210 => x"FF",
		286234 => x"FF",
		287258 => x"FF",
		288282 => x"FF",
		289306 => x"FF",
		290330 => x"FF",
		291354 => x"FF",
		292378 => x"FF",
		293402 => x"FF",
		294426 => x"FF",
		295450 => x"FF",
		296474 => x"FF",
		297498 => x"FF",
		298522 => x"FF",
		299546 => x"FF",
		300570 => x"FF",
		301594 => x"FF",
		302618 => x"FF",
		303642 => x"FF",
		304666 => x"FF",
		305690 => x"FF",
		306714 => x"FF",
		307738 => x"FF",
		308762 => x"FF",
		309786 => x"FF",
		310810 => x"FF",
		311834 => x"FF",
		312858 => x"FF",
		313882 => x"FF",
		314906 => x"FF",
		315930 => x"FF",
		316954 => x"FF",
		317978 => x"FF",
		319002 => x"FF",
		320026 => x"FF",
		321050 => x"FF",
		322074 => x"FF",
		323098 => x"FF",
		324122 => x"FF",
		325146 => x"FF",
		326170 => x"FF",
		327194 => x"FF",
		328218 => x"FF",
		329242 => x"FF",
		330266 => x"FF",
		331290 => x"FF",
		332314 => x"FF",
		333338 => x"FF",
		334362 => x"FF",
		335386 => x"FF",
		336410 => x"FF",
		337434 => x"FF",
		338458 => x"FF",
		339482 => x"FF",
		340506 => x"FF",
		341530 => x"FF",
		342554 => x"FF",
		343578 => x"FF",
		344602 => x"FF",
		345626 => x"FF",
		346650 => x"FF",
		347674 => x"FF",
		348698 => x"FF",
		349722 => x"FF",
		350746 => x"FF",
		351770 => x"FF",
		352794 => x"FF",
		353818 => x"FF",
		354842 => x"FF",
		355866 => x"FF",
		356890 => x"FF",
		357914 => x"FF",
		358938 => x"FF",
		359962 => x"FF",
		360986 => x"FF",
		362010 => x"FF",
		363034 => x"FF",
		364058 => x"FF",
		365082 => x"FF",
		366106 => x"FF",
		367130 => x"FF",
		368154 => x"FF",
		369178 => x"FF",
		370202 => x"FF",
		371226 => x"FF",
		372250 => x"FF",
		373274 => x"FF",
		374298 => x"FF",
		375322 => x"FF",
		376346 => x"FF",
		377370 => x"FF",
		378394 => x"FF",
		379418 => x"FF",
		380442 => x"FF",
		381466 => x"FF",
		382490 => x"FF",
		383514 => x"FF",
		384538 => x"FF",
		385562 => x"FF",
		386586 => x"FF",
		387610 => x"FF",
		388634 => x"FF",
		389658 => x"FF",
		390682 => x"FF",
		391706 => x"FF",
		392730 => x"FF",
		393754 => x"FF",
		394778 => x"FF",
		395802 => x"FF",
		396826 => x"FF",
		397850 => x"FF",
		398874 => x"FF",
		399898 => x"FF",
		400922 => x"FF",
		401946 => x"FF",
		402970 => x"FF",
		403994 => x"FF",
		405018 => x"FF",
		406042 => x"FF",
		407066 => x"FF",
		408090 => x"FF",
		409114 => x"FF",
		410138 => x"FF",
		411162 => x"FF",
		412186 => x"FF",
		413210 => x"FF",
		414234 => x"FF",
		415258 => x"FF",
		416282 => x"FF",
		417306 => x"FF",
		418330 => x"FF",
		419354 => x"FF",
		420378 => x"FF",
		421402 => x"FF",
		422426 => x"FF",
		423450 => x"FF",
		424474 => x"FF",
		425498 => x"FF",
		426522 => x"FF",
		427546 => x"FF",
		428570 => x"FF",
		429594 => x"FF",
		430618 => x"FF",
		431642 => x"FF",
		432666 => x"FF",
		433690 => x"FF",
		434714 => x"FF",
		435738 => x"FF",
		436762 => x"FF",
		437786 => x"FF",
		438810 => x"FF",
		439834 => x"FF",
		440858 => x"FF",
		441882 => x"FF",
		442906 => x"FF",
		443930 => x"FF",
		444954 => x"FF",
		445978 => x"FF",
		447002 => x"FF",
		448026 => x"FF",
		449050 => x"FF",
		450074 => x"FF",
		451098 => x"FF",
		452122 => x"FF",
		453146 => x"FF",
		454170 => x"FF",
		455194 => x"FF",
		456218 => x"FF",
		457242 => x"FF",
		458266 => x"FF",
		459290 => x"FF",
		460314 => x"FF",
		461338 => x"FF",
		462362 => x"FF",
		463386 => x"FF",
		464410 => x"FF",
		465434 => x"FF",
		466458 => x"FF",
		467482 => x"FF",
		468506 => x"FF",
		469530 => x"FF",
		others=> "00000000");
begin

	process (Clk)
	begin
		if (Clk'event and Clk = '1') then
			if (CE = '1') then
				if (Enable_w = '1') then
					VRAM (to_integer(unsigned(Addr_w))) <= Data_in;
				end if;
				Data_out <= VRAM(to_integer(unsigned(Addr_r)));
			else
				NULL;
			end if;
		end if;
	end process;

end Behavioral;

					
