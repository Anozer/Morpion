0 => x"2B",
2 => x"6D",
3 => x"C5",
4 => x"C0",
5 => x"2C",
6 => x"6B",
7 => x"D4",
8 => x"6B",
9 => x"DC",
10 => x"CB",
11 => x"2B",
12 => x"70",
14 => x"2B",
15 => x"71",
16 => x"2C",
17 => x"B1",
19 => x"C0",
20 => x"2B",
21 => x"70",
22 => x"6D",
23 => x"B0",
24 => x"6E",
25 => x"E7",
26 => x"B0",
27 => x"E7",
28 => x"6D",
29 => x"2B",
30 => x"70",
31 => x"6B",
32 => x"C0",
33 => x"B0",
34 => x"6D",
35 => x"E7",
36 => x"6F",
37 => x"B0",
38 => x"E7",
39 => x"2B",
40 => x"70",
42 => x"C0",
43 => x"FF",
44 => x"00",
45 => x"01",
46 => x"F7",
47 => x"08",
48 => x"00",
49 => x"00",
others => x"00"