library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM_X is
	port (CLK : in std_logic;
		  EN : in std_logic;
		  ADDR : in std_logic_vector(13 downto 0);
		  DATA : out std_logic_vector(7 downto 0));
end ROM_X;

architecture Behavioral of ROM_X is

type zone_memoire is array ((2**14)-1 downto 0) of std_logic_vector (7 downto 0);
constant ROM: zone_memoire := (
	0 => "00000000",
	1 => "00000000",
	2 => "00000000",
	3 => "00000000",
	4 => "00000000",
	5 => "00000000",
	6 => "00000000",
	7 => "00000000",
	8 => "00000000",
	9 => "00000000",
	10 => "00000000",
	11 => "00000000",
	12 => "00000000",
	13 => "00000000",
	14 => "00000000",
	15 => "00000000",
	16 => "00000000",
	17 => "00000000",
	18 => "00000000",
	19 => "00000000",
	20 => "00000000",
	21 => "00000000",
	22 => "00000000",
	23 => "00000000",
	24 => "00000000",
	25 => "00000000",
	26 => "00000000",
	27 => "00000000",
	28 => "00000000",
	29 => "00000000",
	30 => "00000000",
	31 => "00000000",
	32 => "00000000",
	33 => "00000000",
	34 => "00000000",
	35 => "00000000",
	36 => "00000000",
	37 => "00000000",
	38 => "00000000",
	39 => "00000000",
	40 => "00000000",
	41 => "00000000",
	42 => "00000000",
	43 => "00000000",
	44 => "00000000",
	45 => "00000000",
	46 => "00000000",
	47 => "00000000",
	48 => "00000000",
	49 => "00000000",
	50 => "00000000",
	51 => "00000000",
	52 => "00000000",
	53 => "00000000",
	54 => "00000000",
	55 => "00000000",
	56 => "00000000",
	57 => "00000000",
	58 => "00000000",
	59 => "00000000",
	60 => "00000000",
	61 => "00000000",
	62 => "00000000",
	63 => "00000000",
	64 => "00000000",
	65 => "00000000",
	66 => "00000000",
	67 => "00000000",
	68 => "00000000",
	69 => "00000000",
	70 => "00000000",
	71 => "00000000",
	72 => "00000000",
	73 => "00000000",
	74 => "00000000",
	75 => "00000000",
	76 => "00000000",
	77 => "00000000",
	78 => "00000000",
	79 => "00000000",
	80 => "00000000",
	81 => "00000000",
	82 => "00000000",
	83 => "00000000",
	84 => "00000000",
	85 => "00000000",
	86 => "00000000",
	87 => "00000000",
	88 => "00000000",
	89 => "00000000",
	90 => "00000000",
	91 => "00000000",
	92 => "00000000",
	93 => "00000000",
	94 => "00000000",
	95 => "00000000",
	96 => "00000000",
	97 => "00000000",
	98 => "00000000",
	99 => "00000000",
	100 => "00000000",
	101 => "00000000",
	102 => "00000000",
	103 => "00000000",
	104 => "00000000",
	105 => "00000000",
	106 => "00000000",
	107 => "00000000",
	108 => "00000000",
	109 => "00000000",
	110 => "00000000",
	111 => "00000000",
	112 => "00000000",
	113 => "00000000",
	114 => "00000000",
	115 => "00000000",
	116 => "00000000",
	117 => "00000000",
	118 => "00000000",
	119 => "00000000",
	128 => "00000000",
	129 => "00000000",
	130 => "00000000",
	131 => "00000000",
	132 => "00000000",
	133 => "00000000",
	134 => "00000000",
	135 => "00000000",
	136 => "00000000",
	137 => "00000000",
	138 => "00000000",
	139 => "00000000",
	140 => "00000000",
	141 => "00000000",
	142 => "00000000",
	143 => "00000000",
	144 => "00000000",
	145 => "00000000",
	146 => "00000000",
	147 => "00000000",
	148 => "00000000",
	149 => "00000000",
	150 => "00000000",
	151 => "00000000",
	152 => "00000000",
	153 => "00000000",
	154 => "00000000",
	155 => "00000000",
	156 => "00000000",
	157 => "00000000",
	158 => "00000000",
	159 => "00000000",
	160 => "00000000",
	161 => "00000000",
	162 => "00000000",
	163 => "00000000",
	164 => "00000000",
	165 => "00000000",
	166 => "00000000",
	167 => "00000000",
	168 => "00000000",
	169 => "00000000",
	170 => "00000000",
	171 => "00000000",
	172 => "00000000",
	173 => "00000000",
	174 => "00000000",
	175 => "00000000",
	176 => "00000000",
	177 => "00000000",
	178 => "00000000",
	179 => "00000000",
	180 => "00000000",
	181 => "00000000",
	182 => "00000000",
	183 => "00000000",
	184 => "00000000",
	185 => "00000000",
	186 => "00000000",
	187 => "00000000",
	188 => "00000000",
	189 => "00000000",
	190 => "00000000",
	191 => "00000000",
	192 => "00000000",
	193 => "00000000",
	194 => "00000000",
	195 => "00000000",
	196 => "00000000",
	197 => "00000000",
	198 => "00000000",
	199 => "00000000",
	200 => "00000000",
	201 => "00000000",
	202 => "00000000",
	203 => "00000000",
	204 => "00000000",
	205 => "00000000",
	206 => "00000000",
	207 => "00000000",
	208 => "00000000",
	209 => "00000000",
	210 => "00000000",
	211 => "00000000",
	212 => "00000000",
	213 => "00000000",
	214 => "00000000",
	215 => "00000000",
	216 => "00000000",
	217 => "00000000",
	218 => "00000000",
	219 => "00000000",
	220 => "00000000",
	221 => "00000000",
	222 => "00000000",
	223 => "00000000",
	224 => "00000000",
	225 => "00000000",
	226 => "00000000",
	227 => "00000000",
	228 => "00000000",
	229 => "00000000",
	230 => "00000000",
	231 => "00000000",
	232 => "00000000",
	233 => "00000000",
	234 => "00000000",
	235 => "00000000",
	236 => "00000000",
	237 => "00000000",
	238 => "00000000",
	239 => "00000000",
	240 => "00000000",
	241 => "00000000",
	242 => "00000000",
	243 => "00000000",
	244 => "00000000",
	245 => "00000000",
	246 => "00000000",
	247 => "00000000",
	256 => "00000000",
	257 => "00000000",
	258 => "00000000",
	259 => "00000000",
	260 => "00000000",
	261 => "00000000",
	262 => "00000000",
	263 => "00000000",
	264 => "00000000",
	265 => "00000000",
	266 => "00000000",
	267 => "00000000",
	268 => "00000000",
	269 => "00000000",
	270 => "00000000",
	271 => "00000000",
	272 => "00000000",
	273 => "00000000",
	274 => "00000000",
	275 => "00000000",
	276 => "00000000",
	277 => "00000000",
	278 => "00000000",
	279 => "00000000",
	280 => "00000000",
	281 => "00000000",
	282 => "00000000",
	283 => "00000000",
	284 => "00000000",
	285 => "00000000",
	286 => "00000000",
	287 => "00000000",
	288 => "00000000",
	289 => "00000000",
	290 => "00000000",
	291 => "00000000",
	292 => "00000000",
	293 => "00000000",
	294 => "00000000",
	295 => "00000000",
	296 => "00000000",
	297 => "00000000",
	298 => "00000000",
	299 => "00000000",
	300 => "00000000",
	301 => "00000000",
	302 => "00000000",
	303 => "00000000",
	304 => "00000000",
	305 => "00000000",
	306 => "00000000",
	307 => "00000000",
	308 => "00000000",
	309 => "00000000",
	310 => "00000000",
	311 => "00000000",
	312 => "00000000",
	313 => "00000000",
	314 => "00000000",
	315 => "00000000",
	316 => "00000000",
	317 => "00000000",
	318 => "00000000",
	319 => "00000000",
	320 => "00000000",
	321 => "00000000",
	322 => "00000000",
	323 => "00000000",
	324 => "00000000",
	325 => "00000000",
	326 => "00000000",
	327 => "00000000",
	328 => "00000000",
	329 => "00000000",
	330 => "00000000",
	331 => "00000000",
	332 => "00000000",
	333 => "00000000",
	334 => "00000000",
	335 => "00000000",
	336 => "00000000",
	337 => "00000000",
	338 => "00000000",
	339 => "00000000",
	340 => "00000000",
	341 => "00000000",
	342 => "00000000",
	343 => "00000000",
	344 => "00000000",
	345 => "00000000",
	346 => "00000000",
	347 => "00000000",
	348 => "00000000",
	349 => "00000000",
	350 => "00000000",
	351 => "00000000",
	352 => "00000000",
	353 => "00000000",
	354 => "00000000",
	355 => "00000000",
	356 => "00000000",
	357 => "00000000",
	358 => "00000000",
	359 => "00000000",
	360 => "00000000",
	361 => "00000000",
	362 => "00000000",
	363 => "00000000",
	364 => "00000000",
	365 => "00000000",
	366 => "00000000",
	367 => "00000000",
	368 => "00000000",
	369 => "00000000",
	370 => "00000000",
	371 => "00000000",
	372 => "00000000",
	373 => "00000000",
	374 => "00000000",
	375 => "00000000",
	384 => "00000000",
	385 => "00000000",
	386 => "00000000",
	387 => "00000000",
	388 => "00000000",
	389 => "00000000",
	390 => "00000000",
	391 => "00000000",
	392 => "00000000",
	393 => "00000000",
	394 => "00000000",
	395 => "00000000",
	396 => "00000000",
	397 => "00000000",
	398 => "00000000",
	399 => "00000000",
	400 => "00000000",
	401 => "00000000",
	402 => "00000000",
	403 => "00000000",
	404 => "00000000",
	405 => "00000000",
	406 => "00000000",
	407 => "00000000",
	408 => "00000000",
	409 => "00000000",
	410 => "00000000",
	411 => "00000000",
	412 => "00000000",
	413 => "00000000",
	414 => "00000000",
	415 => "00000000",
	416 => "00000000",
	417 => "00000000",
	418 => "00000000",
	419 => "00000000",
	420 => "00000000",
	421 => "00000000",
	422 => "00000000",
	423 => "00000000",
	424 => "00000000",
	425 => "00000000",
	426 => "00000000",
	427 => "00000000",
	428 => "00000000",
	429 => "00000000",
	430 => "00000000",
	431 => "00000000",
	432 => "00000000",
	433 => "00000000",
	434 => "00000000",
	435 => "00000000",
	436 => "00000000",
	437 => "00000000",
	438 => "00000000",
	439 => "00000000",
	440 => "00000000",
	441 => "00000000",
	442 => "00000000",
	443 => "00000000",
	444 => "00000000",
	445 => "00000000",
	446 => "00000000",
	447 => "00000000",
	448 => "00000000",
	449 => "00000000",
	450 => "00000000",
	451 => "00000000",
	452 => "00000000",
	453 => "00000000",
	454 => "00000000",
	455 => "00000000",
	456 => "00000000",
	457 => "00000000",
	458 => "00000000",
	459 => "00000000",
	460 => "00000000",
	461 => "00000000",
	462 => "00000000",
	463 => "00000000",
	464 => "00000000",
	465 => "00000000",
	466 => "00000000",
	467 => "00000000",
	468 => "00000000",
	469 => "00000000",
	470 => "00000000",
	471 => "00000000",
	472 => "00000000",
	473 => "00000000",
	474 => "00000000",
	475 => "00000000",
	476 => "00000000",
	477 => "00000000",
	478 => "00000000",
	479 => "00000000",
	480 => "00000000",
	481 => "00000000",
	482 => "00000000",
	483 => "00000000",
	484 => "00000000",
	485 => "00000000",
	486 => "00000000",
	487 => "00000000",
	488 => "00000000",
	489 => "00000000",
	490 => "00000000",
	491 => "00000000",
	492 => "00000000",
	493 => "00000000",
	494 => "00000000",
	495 => "00000000",
	496 => "00000000",
	497 => "00000000",
	498 => "00000000",
	499 => "00000000",
	500 => "00000000",
	501 => "00000000",
	502 => "00000000",
	503 => "00000000",
	512 => "00000000",
	513 => "00000000",
	514 => "00000000",
	515 => "00000000",
	516 => "00000000",
	517 => "00000000",
	518 => "00000000",
	519 => "00000000",
	520 => "00000000",
	521 => "00000000",
	522 => "00000000",
	523 => "00000000",
	524 => "00000000",
	525 => "00000000",
	526 => "00000000",
	527 => "00000000",
	528 => "00000000",
	529 => "00000000",
	530 => "00000000",
	531 => "00000000",
	532 => "00000000",
	533 => "00000000",
	534 => "00000000",
	535 => "00000000",
	536 => "00000000",
	537 => "00000000",
	538 => "00000000",
	539 => "00000000",
	540 => "00000000",
	541 => "00000000",
	542 => "00000000",
	543 => "00000000",
	544 => "00000000",
	545 => "00000000",
	546 => "00000000",
	547 => "00000000",
	548 => "00000000",
	549 => "00000000",
	550 => "00000000",
	551 => "00000000",
	552 => "00000000",
	553 => "00000000",
	554 => "00000000",
	555 => "00000000",
	556 => "00000000",
	557 => "00000000",
	558 => "00000000",
	559 => "00000000",
	560 => "00000000",
	561 => "00000000",
	562 => "00000000",
	563 => "00000000",
	564 => "00000000",
	565 => "00000000",
	566 => "00000000",
	567 => "00000000",
	568 => "00000000",
	569 => "00000000",
	570 => "00000000",
	571 => "00000000",
	572 => "00000000",
	573 => "00000000",
	574 => "00000000",
	575 => "00000000",
	576 => "00000000",
	577 => "00000000",
	578 => "00000000",
	579 => "00000000",
	580 => "00000000",
	581 => "00000000",
	582 => "00000000",
	583 => "00000000",
	584 => "00000000",
	585 => "00000000",
	586 => "00000000",
	587 => "00000000",
	588 => "00000000",
	589 => "00000000",
	590 => "00000000",
	591 => "00000000",
	592 => "00000000",
	593 => "00000000",
	594 => "00000000",
	595 => "00000000",
	596 => "00000000",
	597 => "00000000",
	598 => "00000000",
	599 => "00000000",
	600 => "00000000",
	601 => "00000000",
	602 => "00000000",
	603 => "00000000",
	604 => "00000000",
	605 => "00000000",
	606 => "00000000",
	607 => "00000000",
	608 => "00000000",
	609 => "00000000",
	610 => "00000000",
	611 => "00000000",
	612 => "00000000",
	613 => "00000000",
	614 => "00000000",
	615 => "00000000",
	616 => "00000000",
	617 => "00000000",
	618 => "00000000",
	619 => "00000000",
	620 => "00000000",
	621 => "00000000",
	622 => "00000000",
	623 => "00000000",
	624 => "00000000",
	625 => "00000000",
	626 => "00000000",
	627 => "00000000",
	628 => "00000000",
	629 => "00000000",
	630 => "00000000",
	631 => "00000000",
	640 => "00000000",
	641 => "00000000",
	642 => "00000000",
	643 => "00000000",
	644 => "00000000",
	645 => "00000000",
	646 => "00000000",
	647 => "00000000",
	648 => "00000000",
	649 => "00000000",
	650 => "00000000",
	651 => "00000000",
	652 => "00000000",
	653 => "00000000",
	654 => "00000000",
	655 => "00000000",
	656 => "00000000",
	657 => "00000000",
	658 => "00000000",
	659 => "00000000",
	660 => "00000000",
	661 => "00000000",
	662 => "00000000",
	663 => "00000000",
	664 => "00000000",
	665 => "00000000",
	666 => "00000000",
	667 => "00000000",
	668 => "00000000",
	669 => "00000000",
	670 => "00000000",
	671 => "00000000",
	672 => "00000000",
	673 => "00000000",
	674 => "00000000",
	675 => "00000000",
	676 => "00000000",
	677 => "00000000",
	678 => "00000000",
	679 => "00000000",
	680 => "00000000",
	681 => "00000000",
	682 => "00000000",
	683 => "00000000",
	684 => "00000000",
	685 => "00000000",
	686 => "00000000",
	687 => "00000000",
	688 => "00000000",
	689 => "00000000",
	690 => "00000000",
	691 => "00000000",
	692 => "00000000",
	693 => "00000000",
	694 => "00000000",
	695 => "00000000",
	696 => "00000000",
	697 => "00000000",
	698 => "00000000",
	699 => "00000000",
	700 => "00000000",
	701 => "00000000",
	702 => "00000000",
	703 => "00000000",
	704 => "00000000",
	705 => "00000000",
	706 => "00000000",
	707 => "00000000",
	708 => "00000000",
	709 => "00000000",
	710 => "00000000",
	711 => "00000000",
	712 => "00000000",
	713 => "00000000",
	714 => "00000000",
	715 => "00000000",
	716 => "00000000",
	717 => "00000000",
	718 => "00000000",
	719 => "00000000",
	720 => "00000000",
	721 => "00000000",
	722 => "00000000",
	723 => "00000000",
	724 => "00000000",
	725 => "00000000",
	726 => "00000000",
	727 => "00000000",
	728 => "00000000",
	729 => "00000000",
	730 => "00000000",
	731 => "00000000",
	732 => "00000000",
	733 => "00000000",
	734 => "00000000",
	735 => "00000000",
	736 => "00000000",
	737 => "00000000",
	738 => "00000000",
	739 => "00000000",
	740 => "00000000",
	741 => "00000000",
	742 => "00000000",
	743 => "00000000",
	744 => "00000000",
	745 => "00000000",
	746 => "00000000",
	747 => "00000000",
	748 => "00000000",
	749 => "00000000",
	750 => "00000000",
	751 => "00000000",
	752 => "00000000",
	753 => "00000000",
	754 => "00000000",
	755 => "00000000",
	756 => "00000000",
	757 => "00000000",
	758 => "00000000",
	759 => "00000000",
	768 => "00000000",
	769 => "00000000",
	770 => "00000000",
	771 => "00000000",
	772 => "00000000",
	773 => "00000000",
	774 => "00000000",
	775 => "00000000",
	776 => "00000000",
	777 => "00000000",
	778 => "00000000",
	779 => "00000000",
	780 => "00000000",
	781 => "00000000",
	782 => "00000000",
	783 => "00000000",
	784 => "00000000",
	785 => "00000000",
	786 => "00000000",
	787 => "00000000",
	788 => "00000000",
	789 => "00000000",
	790 => "00000000",
	791 => "00000000",
	792 => "00000000",
	793 => "00000000",
	794 => "00000000",
	795 => "00000000",
	796 => "00000000",
	797 => "00000000",
	798 => "00000000",
	799 => "00000000",
	800 => "00000000",
	801 => "00000000",
	802 => "00000000",
	803 => "00000000",
	804 => "00000000",
	805 => "00000000",
	806 => "00000000",
	807 => "00000000",
	808 => "00000000",
	809 => "00000000",
	810 => "00000000",
	811 => "00000000",
	812 => "00000000",
	813 => "00000000",
	814 => "00000000",
	815 => "00000000",
	816 => "00000000",
	817 => "00000000",
	818 => "00000000",
	819 => "00000000",
	820 => "00000000",
	821 => "00000000",
	822 => "00000000",
	823 => "00000000",
	824 => "00000000",
	825 => "00000000",
	826 => "00000000",
	827 => "00000000",
	828 => "00000000",
	829 => "00000000",
	830 => "00000000",
	831 => "00000000",
	832 => "00000000",
	833 => "00000000",
	834 => "00000000",
	835 => "00000000",
	836 => "00000000",
	837 => "00000000",
	838 => "00000000",
	839 => "00000000",
	840 => "00000000",
	841 => "00000000",
	842 => "00000000",
	843 => "00000000",
	844 => "00000000",
	845 => "00000000",
	846 => "00000000",
	847 => "00000000",
	848 => "00000000",
	849 => "00000000",
	850 => "00000000",
	851 => "00000000",
	852 => "00000000",
	853 => "00000000",
	854 => "00000000",
	855 => "00000000",
	856 => "00000000",
	857 => "00000000",
	858 => "00000000",
	859 => "00000000",
	860 => "00000000",
	861 => "00000000",
	862 => "00000000",
	863 => "00000000",
	864 => "00000000",
	865 => "00000000",
	866 => "00000000",
	867 => "00000000",
	868 => "00000000",
	869 => "00000000",
	870 => "00000000",
	871 => "00000000",
	872 => "00000000",
	873 => "00000000",
	874 => "00000000",
	875 => "00000000",
	876 => "00000000",
	877 => "00000000",
	878 => "00000000",
	879 => "00000000",
	880 => "00000000",
	881 => "00000000",
	882 => "00000000",
	883 => "00000000",
	884 => "00000000",
	885 => "00000000",
	886 => "00000000",
	887 => "00000000",
	896 => "00000000",
	897 => "00000000",
	898 => "00000000",
	899 => "00000000",
	900 => "00000000",
	901 => "00000000",
	902 => "00000000",
	903 => "00000000",
	904 => "00000000",
	905 => "00000000",
	906 => "00000000",
	907 => "00000000",
	908 => "00000000",
	909 => "00000000",
	910 => "00000000",
	911 => "00000000",
	912 => "00000000",
	913 => "00000000",
	914 => "00000000",
	915 => "00000000",
	916 => "00000000",
	917 => "00000000",
	918 => "00000000",
	919 => "00000000",
	920 => "00000000",
	921 => "00000000",
	922 => "00000000",
	923 => "00000000",
	924 => "00000000",
	925 => "00000000",
	926 => "00000000",
	927 => "00000000",
	928 => "00000000",
	929 => "00000000",
	930 => "00000000",
	931 => "00000000",
	932 => "00000000",
	933 => "00000000",
	934 => "00000000",
	935 => "00000000",
	936 => "00000000",
	937 => "00000000",
	938 => "00000000",
	939 => "00000000",
	940 => "00000000",
	941 => "00000000",
	942 => "00000000",
	943 => "00000000",
	944 => "00000000",
	945 => "00000000",
	946 => "00000000",
	947 => "00000000",
	948 => "00000000",
	949 => "00000000",
	950 => "00000000",
	951 => "00000000",
	952 => "00000000",
	953 => "00000000",
	954 => "00000000",
	955 => "00000000",
	956 => "00000000",
	957 => "00000000",
	958 => "00000000",
	959 => "00000000",
	960 => "00000000",
	961 => "00000000",
	962 => "00000000",
	963 => "00000000",
	964 => "00000000",
	965 => "00000000",
	966 => "00000000",
	967 => "00000000",
	968 => "00000000",
	969 => "00000000",
	970 => "00000000",
	971 => "00000000",
	972 => "00000000",
	973 => "00000000",
	974 => "00000000",
	975 => "00000000",
	976 => "00000000",
	977 => "00000000",
	978 => "00000000",
	979 => "00000000",
	980 => "00000000",
	981 => "00000000",
	982 => "00000000",
	983 => "00000000",
	984 => "00000000",
	985 => "00000000",
	986 => "00000000",
	987 => "00000000",
	988 => "00000000",
	989 => "00000000",
	990 => "00000000",
	991 => "00000000",
	992 => "00000000",
	993 => "00000000",
	994 => "00000000",
	995 => "00000000",
	996 => "00000000",
	997 => "00000000",
	998 => "00000000",
	999 => "00000000",
	1000 => "00000000",
	1001 => "00000000",
	1002 => "00000000",
	1003 => "00000000",
	1004 => "00000000",
	1005 => "00000000",
	1006 => "00000000",
	1007 => "00000000",
	1008 => "00000000",
	1009 => "00000000",
	1010 => "00000000",
	1011 => "00000000",
	1012 => "00000000",
	1013 => "00000000",
	1014 => "00000000",
	1015 => "00000000",
	1024 => "00000000",
	1025 => "00000000",
	1026 => "00000000",
	1027 => "00000000",
	1028 => "00000000",
	1029 => "00000000",
	1030 => "00000000",
	1031 => "00000000",
	1032 => "00000000",
	1033 => "00000000",
	1034 => "00000000",
	1035 => "00000000",
	1036 => "00000000",
	1037 => "00000000",
	1038 => "00000000",
	1039 => "00000000",
	1040 => "00000000",
	1041 => "00000000",
	1042 => "00000000",
	1043 => "00000000",
	1044 => "00000000",
	1045 => "00000000",
	1046 => "00000000",
	1047 => "00000000",
	1048 => "00000000",
	1049 => "00000000",
	1050 => "00000000",
	1051 => "00000000",
	1052 => "00000000",
	1053 => "00000000",
	1054 => "00000000",
	1055 => "00000000",
	1056 => "00000000",
	1057 => "00000000",
	1058 => "00000000",
	1059 => "00000000",
	1060 => "00000000",
	1061 => "00000000",
	1062 => "00000000",
	1063 => "00000000",
	1064 => "00000000",
	1065 => "00000000",
	1066 => "00000000",
	1067 => "00000000",
	1068 => "00000000",
	1069 => "00000000",
	1070 => "00000000",
	1071 => "00000000",
	1072 => "00000000",
	1073 => "00000000",
	1074 => "00000000",
	1075 => "00000000",
	1076 => "00000000",
	1077 => "00000000",
	1078 => "00000000",
	1079 => "00000000",
	1080 => "00000000",
	1081 => "00000000",
	1082 => "00000000",
	1083 => "00000000",
	1084 => "00000000",
	1085 => "00000000",
	1086 => "00000000",
	1087 => "00000000",
	1088 => "00000000",
	1089 => "00000000",
	1090 => "00000000",
	1091 => "00000000",
	1092 => "00000000",
	1093 => "00000000",
	1094 => "00000000",
	1095 => "00000000",
	1096 => "00000000",
	1097 => "00000000",
	1098 => "00000000",
	1099 => "00000000",
	1100 => "00000000",
	1101 => "00000000",
	1102 => "00000000",
	1103 => "00000000",
	1104 => "00000000",
	1105 => "00000000",
	1106 => "00000000",
	1107 => "00000000",
	1108 => "00000000",
	1109 => "00000000",
	1110 => "00000000",
	1111 => "00000000",
	1112 => "00000000",
	1113 => "00000000",
	1114 => "00000000",
	1115 => "00000000",
	1116 => "00000000",
	1117 => "00000000",
	1118 => "00000000",
	1119 => "00000000",
	1120 => "00000000",
	1121 => "00000000",
	1122 => "00000000",
	1123 => "00000000",
	1124 => "00000000",
	1125 => "00000000",
	1126 => "00000000",
	1127 => "00000000",
	1128 => "00000000",
	1129 => "00000000",
	1130 => "00000000",
	1131 => "00000000",
	1132 => "00000000",
	1133 => "00000000",
	1134 => "00000000",
	1135 => "00000000",
	1136 => "00000000",
	1137 => "00000000",
	1138 => "00000000",
	1139 => "00000000",
	1140 => "00000000",
	1141 => "00000000",
	1142 => "00000000",
	1143 => "00000000",
	1152 => "00000000",
	1153 => "00000000",
	1154 => "00000000",
	1155 => "00000000",
	1156 => "00000000",
	1157 => "00000000",
	1158 => "00000000",
	1159 => "00000000",
	1160 => "00000000",
	1161 => "00000000",
	1162 => "00000000",
	1163 => "00000000",
	1164 => "00000000",
	1165 => "00000000",
	1166 => "00000000",
	1167 => "00000000",
	1168 => "00000000",
	1169 => "00000000",
	1170 => "00000000",
	1171 => "00000000",
	1172 => "00000000",
	1173 => "00000000",
	1174 => "00000000",
	1175 => "00000000",
	1176 => "00000000",
	1177 => "00000000",
	1178 => "00000000",
	1179 => "00000000",
	1180 => "00000000",
	1181 => "00000000",
	1182 => "00000000",
	1183 => "00000000",
	1184 => "00000000",
	1185 => "00000000",
	1186 => "00000000",
	1187 => "00000000",
	1188 => "00000000",
	1189 => "00000000",
	1190 => "00000000",
	1191 => "00000000",
	1192 => "00000000",
	1193 => "00000000",
	1194 => "00000000",
	1195 => "00000000",
	1196 => "00000000",
	1197 => "00000000",
	1198 => "00000000",
	1199 => "00000000",
	1200 => "00000000",
	1201 => "00000000",
	1202 => "00000000",
	1203 => "00000000",
	1204 => "00000000",
	1205 => "00000000",
	1206 => "00000000",
	1207 => "00000000",
	1208 => "00000000",
	1209 => "00000000",
	1210 => "00000000",
	1211 => "00000000",
	1212 => "00000000",
	1213 => "00000000",
	1214 => "00000000",
	1215 => "00000000",
	1216 => "00000000",
	1217 => "00000000",
	1218 => "00000000",
	1219 => "00000000",
	1220 => "00000000",
	1221 => "00000000",
	1222 => "00000000",
	1223 => "00000000",
	1224 => "00000000",
	1225 => "00000000",
	1226 => "00000000",
	1227 => "00000000",
	1228 => "00000000",
	1229 => "00000000",
	1230 => "00000000",
	1231 => "00000000",
	1232 => "00000000",
	1233 => "00000000",
	1234 => "00000000",
	1235 => "00000000",
	1236 => "00000000",
	1237 => "00000000",
	1238 => "00000000",
	1239 => "00000000",
	1240 => "00000000",
	1241 => "00000000",
	1242 => "00000000",
	1243 => "00000000",
	1244 => "00000000",
	1245 => "00000000",
	1246 => "00000000",
	1247 => "00000000",
	1248 => "00000000",
	1249 => "00000000",
	1250 => "00000000",
	1251 => "00000000",
	1252 => "00000000",
	1253 => "00000000",
	1254 => "00000000",
	1255 => "00000000",
	1256 => "00000000",
	1257 => "00000000",
	1258 => "00000000",
	1259 => "00000000",
	1260 => "00000000",
	1261 => "00000000",
	1262 => "00000000",
	1263 => "00000000",
	1264 => "00000000",
	1265 => "00000000",
	1266 => "00000000",
	1267 => "00000000",
	1268 => "00000000",
	1269 => "00000000",
	1270 => "00000000",
	1271 => "00000000",
	1280 => "00000000",
	1281 => "00000000",
	1282 => "00000000",
	1283 => "00000000",
	1284 => "00000000",
	1285 => "00000000",
	1286 => "00000000",
	1287 => "00000000",
	1288 => "00000000",
	1289 => "00000000",
	1290 => "00000000",
	1291 => "00000000",
	1292 => "00000000",
	1293 => "00000000",
	1294 => "00000000",
	1295 => "00000000",
	1296 => "00000000",
	1297 => "00000000",
	1298 => "00000000",
	1299 => "00000000",
	1300 => "00000000",
	1301 => "00000000",
	1302 => "00000000",
	1303 => "00000000",
	1304 => "00000000",
	1305 => "00000000",
	1306 => "00000000",
	1307 => "00000000",
	1308 => "00000000",
	1309 => "00000000",
	1310 => "00000000",
	1311 => "00000000",
	1312 => "00000000",
	1313 => "00000000",
	1314 => "00000000",
	1315 => "00000000",
	1316 => "00000000",
	1317 => "00000000",
	1318 => "00000000",
	1319 => "00000000",
	1320 => "00000000",
	1321 => "00000000",
	1322 => "00000000",
	1323 => "00000000",
	1324 => "00000000",
	1325 => "00000000",
	1326 => "00000000",
	1327 => "00000000",
	1328 => "00000000",
	1329 => "00000000",
	1330 => "00000000",
	1331 => "00000000",
	1332 => "00000000",
	1333 => "00000000",
	1334 => "00000000",
	1335 => "00000000",
	1336 => "00000000",
	1337 => "00000000",
	1338 => "00000000",
	1339 => "00000000",
	1340 => "00000000",
	1341 => "00000000",
	1342 => "00000000",
	1343 => "00000000",
	1344 => "00000000",
	1345 => "00000000",
	1346 => "00000000",
	1347 => "00000000",
	1348 => "00000000",
	1349 => "00000000",
	1350 => "00000000",
	1351 => "00000000",
	1352 => "00000000",
	1353 => "00000000",
	1354 => "00000000",
	1355 => "00000000",
	1356 => "00000000",
	1357 => "00000000",
	1358 => "00000000",
	1359 => "00000000",
	1360 => "00000000",
	1361 => "00000000",
	1362 => "00000000",
	1363 => "00000000",
	1364 => "00000000",
	1365 => "00000000",
	1366 => "00000000",
	1367 => "00000000",
	1368 => "00000000",
	1369 => "00000000",
	1370 => "00000000",
	1371 => "00000000",
	1372 => "00000000",
	1373 => "00000000",
	1374 => "00000000",
	1375 => "00000000",
	1376 => "00000000",
	1377 => "00000000",
	1378 => "00000000",
	1379 => "00000000",
	1380 => "00000000",
	1381 => "00000000",
	1382 => "00000000",
	1383 => "00000000",
	1384 => "00000000",
	1385 => "00000000",
	1386 => "00000000",
	1387 => "00000000",
	1388 => "00000000",
	1389 => "00000000",
	1390 => "00000000",
	1391 => "00000000",
	1392 => "00000000",
	1393 => "00000000",
	1394 => "00000000",
	1395 => "00000000",
	1396 => "00000000",
	1397 => "00000000",
	1398 => "00000000",
	1399 => "00000000",
	1408 => "00000000",
	1409 => "00000000",
	1410 => "00000000",
	1411 => "00000000",
	1412 => "00000000",
	1413 => "00000000",
	1414 => "00000000",
	1415 => "00000000",
	1416 => "00000000",
	1417 => "00000000",
	1418 => "00000000",
	1419 => "00000000",
	1420 => "00000000",
	1421 => "00000000",
	1422 => "00000000",
	1423 => "00000000",
	1424 => "00000000",
	1425 => "00000000",
	1426 => "00000000",
	1427 => "00000000",
	1428 => "00000000",
	1429 => "00000000",
	1430 => "00000000",
	1431 => "00000000",
	1432 => "00000000",
	1433 => "00000000",
	1434 => "00000000",
	1435 => "00000000",
	1436 => "00000000",
	1437 => "00000000",
	1438 => "00000000",
	1439 => "00000000",
	1440 => "00000000",
	1441 => "00000000",
	1442 => "00000000",
	1443 => "00000000",
	1444 => "00000000",
	1445 => "00000000",
	1446 => "00000000",
	1447 => "00000000",
	1448 => "00000000",
	1449 => "00000000",
	1450 => "00000000",
	1451 => "00000000",
	1452 => "00000000",
	1453 => "00000000",
	1454 => "00000000",
	1455 => "00000000",
	1456 => "00000000",
	1457 => "00000000",
	1458 => "00000000",
	1459 => "00000000",
	1460 => "00000000",
	1461 => "00000000",
	1462 => "00000000",
	1463 => "00000000",
	1464 => "00000000",
	1465 => "00000000",
	1466 => "00000000",
	1467 => "00000000",
	1468 => "00000000",
	1469 => "00000000",
	1470 => "00000000",
	1471 => "00000000",
	1472 => "00000000",
	1473 => "00000000",
	1474 => "00000000",
	1475 => "00000000",
	1476 => "00000000",
	1477 => "00000000",
	1478 => "00000000",
	1479 => "00000000",
	1480 => "00000000",
	1481 => "00000000",
	1482 => "00000000",
	1483 => "00000000",
	1484 => "00000000",
	1485 => "00000000",
	1486 => "00000000",
	1487 => "00000000",
	1488 => "00000000",
	1489 => "00000000",
	1490 => "00000000",
	1491 => "00000000",
	1492 => "00000000",
	1493 => "00000000",
	1494 => "00000000",
	1495 => "00000000",
	1496 => "00000000",
	1497 => "00000000",
	1498 => "00000000",
	1499 => "00000000",
	1500 => "00000000",
	1501 => "00000000",
	1502 => "00000000",
	1503 => "00000000",
	1504 => "00000000",
	1505 => "00000000",
	1506 => "00000000",
	1507 => "00000000",
	1508 => "00000000",
	1509 => "00000000",
	1510 => "00000000",
	1511 => "00000000",
	1512 => "00000000",
	1513 => "00000000",
	1514 => "00000000",
	1515 => "00000000",
	1516 => "00000000",
	1517 => "00000000",
	1518 => "00000000",
	1519 => "00000000",
	1520 => "00000000",
	1521 => "00000000",
	1522 => "00000000",
	1523 => "00000000",
	1524 => "00000000",
	1525 => "00000000",
	1526 => "00000000",
	1527 => "00000000",
	1536 => "00000000",
	1537 => "00000000",
	1538 => "00000000",
	1539 => "00000000",
	1540 => "00000000",
	1541 => "00000000",
	1542 => "00000000",
	1543 => "00000000",
	1544 => "00000000",
	1545 => "00000000",
	1546 => "00000000",
	1547 => "00000000",
	1548 => "00000000",
	1549 => "00000000",
	1550 => "00000000",
	1551 => "00000000",
	1552 => "00000000",
	1553 => "00000000",
	1554 => "00000000",
	1555 => "00000000",
	1556 => "00000000",
	1557 => "00000000",
	1558 => "00000000",
	1559 => "00000000",
	1560 => "00000000",
	1561 => "00000000",
	1562 => "00000000",
	1563 => "00000000",
	1564 => "00000000",
	1565 => "00000000",
	1566 => "00000000",
	1567 => "00000000",
	1568 => "00000000",
	1569 => "00000000",
	1570 => "00000000",
	1571 => "00000000",
	1572 => "00000000",
	1573 => "00000000",
	1574 => "00000000",
	1575 => "00000000",
	1576 => "00000000",
	1577 => "00000000",
	1578 => "00000000",
	1579 => "00000000",
	1580 => "00000000",
	1581 => "00000000",
	1582 => "00000000",
	1583 => "00000000",
	1584 => "00000000",
	1585 => "00000000",
	1586 => "00000000",
	1587 => "00000000",
	1588 => "00000000",
	1589 => "00000000",
	1590 => "00000000",
	1591 => "00000000",
	1592 => "00000000",
	1593 => "00000000",
	1594 => "00000000",
	1595 => "00000000",
	1596 => "00000000",
	1597 => "00000000",
	1598 => "00000000",
	1599 => "00000000",
	1600 => "00000000",
	1601 => "00000000",
	1602 => "00000000",
	1603 => "00000000",
	1604 => "00000000",
	1605 => "00000000",
	1606 => "00000000",
	1607 => "00000000",
	1608 => "00000000",
	1609 => "00000000",
	1610 => "00000000",
	1611 => "00000000",
	1612 => "00000000",
	1613 => "00000000",
	1614 => "00000000",
	1615 => "00000000",
	1616 => "00000000",
	1617 => "00000000",
	1618 => "00000000",
	1619 => "00000000",
	1620 => "00000000",
	1621 => "00000000",
	1622 => "00000000",
	1623 => "00000000",
	1624 => "00000000",
	1625 => "00000000",
	1626 => "00000000",
	1627 => "00000000",
	1628 => "00000000",
	1629 => "00000000",
	1630 => "00000000",
	1631 => "00000000",
	1632 => "00000000",
	1633 => "00000000",
	1634 => "00000000",
	1635 => "00000000",
	1636 => "00000000",
	1637 => "00000000",
	1638 => "00000000",
	1639 => "00000000",
	1640 => "00000000",
	1641 => "00000000",
	1642 => "00000000",
	1643 => "00000000",
	1644 => "00000000",
	1645 => "00000000",
	1646 => "00000000",
	1647 => "00000000",
	1648 => "00000000",
	1649 => "00000000",
	1650 => "00000000",
	1651 => "00000000",
	1652 => "00000000",
	1653 => "00000000",
	1654 => "00000000",
	1655 => "00000000",
	1664 => "00000000",
	1665 => "00000000",
	1666 => "00000000",
	1667 => "00000000",
	1668 => "00000000",
	1669 => "00000000",
	1670 => "00000000",
	1671 => "00000000",
	1672 => "00000000",
	1673 => "00000000",
	1674 => "00000000",
	1675 => "00000000",
	1676 => "00000000",
	1677 => "00000000",
	1678 => "00000000",
	1679 => "00000000",
	1680 => "00000000",
	1681 => "00000000",
	1682 => "00000000",
	1683 => "00000000",
	1684 => "00000000",
	1685 => "00000000",
	1686 => "00000000",
	1687 => "00000000",
	1688 => "00000000",
	1689 => "00000000",
	1690 => "00000000",
	1691 => "00000000",
	1692 => "00000000",
	1693 => "00000000",
	1694 => "00000000",
	1695 => "00000000",
	1696 => "00000000",
	1697 => "00000000",
	1698 => "00000000",
	1699 => "00000000",
	1700 => "00000000",
	1701 => "00000000",
	1702 => "00000000",
	1703 => "00000000",
	1704 => "00000000",
	1705 => "00000000",
	1706 => "00000000",
	1707 => "00000000",
	1708 => "00000000",
	1709 => "00000000",
	1710 => "00000000",
	1711 => "00000000",
	1712 => "00000000",
	1713 => "00000000",
	1714 => "00000000",
	1715 => "00000000",
	1716 => "00000000",
	1717 => "00000000",
	1718 => "00000000",
	1719 => "00000000",
	1720 => "00000000",
	1721 => "00000000",
	1722 => "00000000",
	1723 => "00000000",
	1724 => "00000000",
	1725 => "00000000",
	1726 => "00000000",
	1727 => "00000000",
	1728 => "00000000",
	1729 => "00000000",
	1730 => "00000000",
	1731 => "00000000",
	1732 => "00000000",
	1733 => "00000000",
	1734 => "00000000",
	1735 => "00000000",
	1736 => "00000000",
	1737 => "00000000",
	1738 => "00000000",
	1739 => "00000000",
	1740 => "00000000",
	1741 => "00000000",
	1742 => "00000000",
	1743 => "00000000",
	1744 => "00000000",
	1745 => "00000000",
	1746 => "00000000",
	1747 => "00000000",
	1748 => "00000000",
	1749 => "00000000",
	1750 => "00000000",
	1751 => "00000000",
	1752 => "00000000",
	1753 => "00000000",
	1754 => "00000000",
	1755 => "00000000",
	1756 => "00000000",
	1757 => "00000000",
	1758 => "00000000",
	1759 => "00000000",
	1760 => "00000000",
	1761 => "00000000",
	1762 => "00000000",
	1763 => "00000000",
	1764 => "00000000",
	1765 => "00000000",
	1766 => "00000000",
	1767 => "00000000",
	1768 => "00000000",
	1769 => "00000000",
	1770 => "00000000",
	1771 => "00000000",
	1772 => "00000000",
	1773 => "00000000",
	1774 => "00000000",
	1775 => "00000000",
	1776 => "00000000",
	1777 => "00000000",
	1778 => "00000000",
	1779 => "00000000",
	1780 => "00000000",
	1781 => "00000000",
	1782 => "00000000",
	1783 => "00000000",
	1792 => "00000000",
	1793 => "00000000",
	1794 => "00000000",
	1795 => "00000000",
	1796 => "00000000",
	1797 => "00000000",
	1798 => "00000000",
	1799 => "00000000",
	1800 => "00000000",
	1801 => "00000000",
	1802 => "00000000",
	1803 => "00000000",
	1804 => "00000000",
	1805 => "00000000",
	1806 => "00000000",
	1807 => "00000000",
	1808 => "00000000",
	1809 => "00000000",
	1810 => "00000000",
	1811 => "00000000",
	1812 => "00000000",
	1813 => "00000000",
	1814 => "00000000",
	1815 => "00000000",
	1816 => "00000000",
	1817 => "00000000",
	1818 => "00000000",
	1819 => "00000000",
	1820 => "00000000",
	1821 => "00000000",
	1822 => "00000000",
	1823 => "00000000",
	1824 => "00000000",
	1825 => "00000000",
	1826 => "00000000",
	1827 => "00000000",
	1828 => "00000000",
	1829 => "00000000",
	1830 => "00000000",
	1831 => "00000000",
	1832 => "00000000",
	1833 => "00000000",
	1834 => "00000000",
	1835 => "00000000",
	1836 => "00000000",
	1837 => "00000000",
	1838 => "00000000",
	1839 => "00000000",
	1840 => "00000000",
	1841 => "00000000",
	1842 => "00000000",
	1843 => "00000000",
	1844 => "00000000",
	1845 => "00000000",
	1846 => "00000000",
	1847 => "00000000",
	1848 => "00000000",
	1849 => "00000000",
	1850 => "00000000",
	1851 => "00000000",
	1852 => "00000000",
	1853 => "00000000",
	1854 => "00000000",
	1855 => "00000000",
	1856 => "00000000",
	1857 => "00000000",
	1858 => "00000000",
	1859 => "00000000",
	1860 => "00000000",
	1861 => "00000000",
	1862 => "00000000",
	1863 => "00000000",
	1864 => "00000000",
	1865 => "00000000",
	1866 => "00000000",
	1867 => "00000000",
	1868 => "00000000",
	1869 => "00000000",
	1870 => "00000000",
	1871 => "00000000",
	1872 => "00000000",
	1873 => "00000000",
	1874 => "00000000",
	1875 => "00000000",
	1876 => "00000000",
	1877 => "00000000",
	1878 => "00000000",
	1879 => "00000000",
	1880 => "00000000",
	1881 => "00000000",
	1882 => "00000000",
	1883 => "00000000",
	1884 => "00000000",
	1885 => "00000000",
	1886 => "00000000",
	1887 => "00000000",
	1888 => "00000000",
	1889 => "00000000",
	1890 => "00000000",
	1891 => "00000000",
	1892 => "00000000",
	1893 => "00000000",
	1894 => "00000000",
	1895 => "00000000",
	1896 => "00000000",
	1897 => "00000000",
	1898 => "00000000",
	1899 => "00000000",
	1900 => "00000000",
	1901 => "00000000",
	1902 => "00000000",
	1903 => "00000000",
	1904 => "00000000",
	1905 => "00000000",
	1906 => "00000000",
	1907 => "00000000",
	1908 => "00000000",
	1909 => "00000000",
	1910 => "00000000",
	1911 => "00000000",
	1920 => "00000000",
	1921 => "00000000",
	1922 => "00000000",
	1923 => "00000000",
	1924 => "00000000",
	1925 => "00000000",
	1926 => "00000000",
	1927 => "00000000",
	1928 => "00000000",
	1929 => "00000000",
	1930 => "00000000",
	1931 => "00000000",
	1932 => "00000000",
	1933 => "00000000",
	1934 => "00000000",
	1935 => "00000000",
	1936 => "00000000",
	1937 => "00000000",
	1938 => "00000000",
	1939 => "00000000",
	1940 => "00000000",
	1941 => "00000000",
	1942 => "00000000",
	1943 => "00000000",
	1944 => "00000000",
	1945 => "00000000",
	1946 => "00000000",
	1947 => "00000000",
	1948 => "00000000",
	1949 => "00000000",
	1950 => "00000000",
	1951 => "00000000",
	1952 => "00000000",
	1953 => "00000000",
	1954 => "00000000",
	1955 => "00000000",
	1956 => "00000000",
	1957 => "00000000",
	1958 => "00000000",
	1959 => "00000000",
	1960 => "00000000",
	1961 => "00000000",
	1962 => "00000000",
	1963 => "00000000",
	1964 => "00000000",
	1965 => "00000000",
	1966 => "00000000",
	1967 => "00000000",
	1968 => "00000000",
	1969 => "00000000",
	1970 => "00000000",
	1971 => "00000000",
	1972 => "00000000",
	1973 => "00000000",
	1974 => "00000000",
	1975 => "00000000",
	1976 => "00000000",
	1977 => "00000000",
	1978 => "00000000",
	1979 => "00000000",
	1980 => "00000000",
	1981 => "00000000",
	1982 => "00000000",
	1983 => "00000000",
	1984 => "00000000",
	1985 => "00000000",
	1986 => "00000000",
	1987 => "00000000",
	1988 => "00000000",
	1989 => "00000000",
	1990 => "00000000",
	1991 => "00000000",
	1992 => "00000000",
	1993 => "00000000",
	1994 => "00000000",
	1995 => "00000000",
	1996 => "00000000",
	1997 => "00000000",
	1998 => "00000000",
	1999 => "00000000",
	2000 => "00000000",
	2001 => "00000000",
	2002 => "00000000",
	2003 => "00000000",
	2004 => "00000000",
	2005 => "00000000",
	2006 => "00000000",
	2007 => "00000000",
	2008 => "00000000",
	2009 => "00000000",
	2010 => "00000000",
	2011 => "00000000",
	2012 => "00000000",
	2013 => "00000000",
	2014 => "00000000",
	2015 => "00000000",
	2016 => "00000000",
	2017 => "00000000",
	2018 => "00000000",
	2019 => "00000000",
	2020 => "00000000",
	2021 => "00000000",
	2022 => "00000000",
	2023 => "00000000",
	2024 => "00000000",
	2025 => "00000000",
	2026 => "00000000",
	2027 => "00000000",
	2028 => "00000000",
	2029 => "00000000",
	2030 => "00000000",
	2031 => "00000000",
	2032 => "00000000",
	2033 => "00000000",
	2034 => "00000000",
	2035 => "00000000",
	2036 => "00000000",
	2037 => "00000000",
	2038 => "00000000",
	2039 => "00000000",
	2048 => "00000000",
	2049 => "00000000",
	2050 => "00000000",
	2051 => "00000000",
	2052 => "00000000",
	2053 => "00000000",
	2054 => "00000000",
	2055 => "00000000",
	2056 => "00000000",
	2057 => "00000000",
	2058 => "00000000",
	2059 => "00000000",
	2060 => "00000000",
	2061 => "00000000",
	2062 => "00000000",
	2063 => "00000000",
	2064 => "00000000",
	2065 => "00000000",
	2066 => "00000000",
	2067 => "00000000",
	2068 => "00000000",
	2069 => "00000000",
	2070 => "00000000",
	2071 => "00000000",
	2072 => "00000000",
	2073 => "00000000",
	2074 => "00000000",
	2075 => "00000000",
	2076 => "00000000",
	2077 => "00000000",
	2078 => "00000000",
	2079 => "00000000",
	2080 => "00000000",
	2081 => "00000000",
	2082 => "00000000",
	2083 => "00000000",
	2084 => "00000000",
	2085 => "00000000",
	2086 => "00000000",
	2087 => "00000000",
	2088 => "00000000",
	2089 => "00000000",
	2090 => "00000000",
	2091 => "00000000",
	2092 => "00000000",
	2093 => "00000000",
	2094 => "00000000",
	2095 => "00000000",
	2096 => "00000000",
	2097 => "00000000",
	2098 => "00000000",
	2099 => "00000000",
	2100 => "00000000",
	2101 => "00000000",
	2102 => "00000000",
	2103 => "00000000",
	2104 => "00000000",
	2105 => "00000000",
	2106 => "00000000",
	2107 => "00000000",
	2108 => "00000000",
	2109 => "00000000",
	2110 => "00000000",
	2111 => "00000000",
	2112 => "00000000",
	2113 => "00000000",
	2114 => "00000000",
	2115 => "00000000",
	2116 => "00000000",
	2117 => "00000000",
	2118 => "00000000",
	2119 => "00000000",
	2120 => "00000000",
	2121 => "00000000",
	2122 => "00000000",
	2123 => "00000000",
	2124 => "00000000",
	2125 => "00000000",
	2126 => "00000000",
	2127 => "00000000",
	2128 => "00000000",
	2129 => "00000000",
	2130 => "00000000",
	2131 => "00000000",
	2132 => "00000000",
	2133 => "00000000",
	2134 => "00000000",
	2135 => "00000000",
	2136 => "00000000",
	2137 => "00000000",
	2138 => "00000000",
	2139 => "00000000",
	2140 => "00000000",
	2141 => "00000000",
	2142 => "00000000",
	2143 => "00000000",
	2144 => "00000000",
	2145 => "00000000",
	2146 => "00000000",
	2147 => "00000000",
	2148 => "00000000",
	2149 => "00000000",
	2150 => "00000000",
	2151 => "00000000",
	2152 => "00000000",
	2153 => "00000000",
	2154 => "00000000",
	2155 => "00000000",
	2156 => "00000000",
	2157 => "00000000",
	2158 => "00000000",
	2159 => "00000000",
	2160 => "00000000",
	2161 => "00000000",
	2162 => "00000000",
	2163 => "00000000",
	2164 => "00000000",
	2165 => "00000000",
	2166 => "00000000",
	2167 => "00000000",
	2176 => "00000000",
	2177 => "00000000",
	2178 => "00000000",
	2179 => "00000000",
	2180 => "00000000",
	2181 => "00000000",
	2182 => "00000000",
	2183 => "00000000",
	2184 => "00000000",
	2185 => "00000000",
	2186 => "00000000",
	2187 => "00000000",
	2188 => "00000000",
	2189 => "00000000",
	2190 => "00000000",
	2191 => "00000000",
	2192 => "00000000",
	2193 => "00000000",
	2194 => "11111111",
	2195 => "11111111",
	2196 => "11111111",
	2197 => "11111111",
	2198 => "11111111",
	2199 => "00000000",
	2200 => "00000000",
	2201 => "00000000",
	2202 => "00000000",
	2203 => "00000000",
	2204 => "00000000",
	2205 => "00000000",
	2206 => "00000000",
	2207 => "00000000",
	2208 => "00000000",
	2209 => "00000000",
	2210 => "00000000",
	2211 => "00000000",
	2212 => "00000000",
	2213 => "00000000",
	2214 => "00000000",
	2215 => "00000000",
	2216 => "00000000",
	2217 => "00000000",
	2218 => "00000000",
	2219 => "00000000",
	2220 => "00000000",
	2221 => "00000000",
	2222 => "00000000",
	2223 => "00000000",
	2224 => "00000000",
	2225 => "00000000",
	2226 => "00000000",
	2227 => "00000000",
	2228 => "00000000",
	2229 => "00000000",
	2230 => "00000000",
	2231 => "00000000",
	2232 => "00000000",
	2233 => "00000000",
	2234 => "00000000",
	2235 => "00000000",
	2236 => "00000000",
	2237 => "00000000",
	2238 => "00000000",
	2239 => "00000000",
	2240 => "00000000",
	2241 => "00000000",
	2242 => "00000000",
	2243 => "00000000",
	2244 => "00000000",
	2245 => "00000000",
	2246 => "00000000",
	2247 => "00000000",
	2248 => "00000000",
	2249 => "00000000",
	2250 => "00000000",
	2251 => "00000000",
	2252 => "00000000",
	2253 => "00000000",
	2254 => "00000000",
	2255 => "00000000",
	2256 => "00000000",
	2257 => "00000000",
	2258 => "00000000",
	2259 => "00000000",
	2260 => "00000000",
	2261 => "00000000",
	2262 => "00000000",
	2263 => "00000000",
	2264 => "00000000",
	2265 => "00000000",
	2266 => "00000000",
	2267 => "00000000",
	2268 => "00000000",
	2269 => "00000000",
	2270 => "00000000",
	2271 => "00000000",
	2272 => "00000000",
	2273 => "00000000",
	2274 => "11111111",
	2275 => "11111111",
	2276 => "11111111",
	2277 => "11111111",
	2278 => "11111111",
	2279 => "00000000",
	2280 => "00000000",
	2281 => "00000000",
	2282 => "00000000",
	2283 => "00000000",
	2284 => "00000000",
	2285 => "00000000",
	2286 => "00000000",
	2287 => "00000000",
	2288 => "00000000",
	2289 => "00000000",
	2290 => "00000000",
	2291 => "00000000",
	2292 => "00000000",
	2293 => "00000000",
	2294 => "00000000",
	2295 => "00000000",
	2304 => "00000000",
	2305 => "00000000",
	2306 => "00000000",
	2307 => "00000000",
	2308 => "00000000",
	2309 => "00000000",
	2310 => "00000000",
	2311 => "00000000",
	2312 => "00000000",
	2313 => "00000000",
	2314 => "00000000",
	2315 => "00000000",
	2316 => "00000000",
	2317 => "00000000",
	2318 => "00000000",
	2319 => "00000000",
	2320 => "00000000",
	2321 => "11111111",
	2322 => "11111111",
	2323 => "11111111",
	2324 => "11111111",
	2325 => "11111111",
	2326 => "11111111",
	2327 => "11111111",
	2328 => "00000000",
	2329 => "00000000",
	2330 => "00000000",
	2331 => "00000000",
	2332 => "00000000",
	2333 => "00000000",
	2334 => "00000000",
	2335 => "00000000",
	2336 => "00000000",
	2337 => "00000000",
	2338 => "00000000",
	2339 => "00000000",
	2340 => "00000000",
	2341 => "00000000",
	2342 => "00000000",
	2343 => "00000000",
	2344 => "00000000",
	2345 => "00000000",
	2346 => "00000000",
	2347 => "00000000",
	2348 => "00000000",
	2349 => "00000000",
	2350 => "00000000",
	2351 => "00000000",
	2352 => "00000000",
	2353 => "00000000",
	2354 => "00000000",
	2355 => "00000000",
	2356 => "00000000",
	2357 => "00000000",
	2358 => "00000000",
	2359 => "00000000",
	2360 => "00000000",
	2361 => "00000000",
	2362 => "00000000",
	2363 => "00000000",
	2364 => "00000000",
	2365 => "00000000",
	2366 => "00000000",
	2367 => "00000000",
	2368 => "00000000",
	2369 => "00000000",
	2370 => "00000000",
	2371 => "00000000",
	2372 => "00000000",
	2373 => "00000000",
	2374 => "00000000",
	2375 => "00000000",
	2376 => "00000000",
	2377 => "00000000",
	2378 => "00000000",
	2379 => "00000000",
	2380 => "00000000",
	2381 => "00000000",
	2382 => "00000000",
	2383 => "00000000",
	2384 => "00000000",
	2385 => "00000000",
	2386 => "00000000",
	2387 => "00000000",
	2388 => "00000000",
	2389 => "00000000",
	2390 => "00000000",
	2391 => "00000000",
	2392 => "00000000",
	2393 => "00000000",
	2394 => "00000000",
	2395 => "00000000",
	2396 => "00000000",
	2397 => "00000000",
	2398 => "00000000",
	2399 => "00000000",
	2400 => "00000000",
	2401 => "11111111",
	2402 => "11111111",
	2403 => "11111111",
	2404 => "11111111",
	2405 => "11111111",
	2406 => "11111111",
	2407 => "11111111",
	2408 => "00000000",
	2409 => "00000000",
	2410 => "00000000",
	2411 => "00000000",
	2412 => "00000000",
	2413 => "00000000",
	2414 => "00000000",
	2415 => "00000000",
	2416 => "00000000",
	2417 => "00000000",
	2418 => "00000000",
	2419 => "00000000",
	2420 => "00000000",
	2421 => "00000000",
	2422 => "00000000",
	2423 => "00000000",
	2432 => "00000000",
	2433 => "00000000",
	2434 => "00000000",
	2435 => "00000000",
	2436 => "00000000",
	2437 => "00000000",
	2438 => "00000000",
	2439 => "00000000",
	2440 => "00000000",
	2441 => "00000000",
	2442 => "00000000",
	2443 => "00000000",
	2444 => "00000000",
	2445 => "00000000",
	2446 => "00000000",
	2447 => "00000000",
	2448 => "00000000",
	2449 => "11111111",
	2450 => "11111111",
	2451 => "11111111",
	2452 => "11111111",
	2453 => "11111111",
	2454 => "11111111",
	2455 => "11111111",
	2456 => "11111111",
	2457 => "00000000",
	2458 => "00000000",
	2459 => "00000000",
	2460 => "00000000",
	2461 => "00000000",
	2462 => "00000000",
	2463 => "00000000",
	2464 => "00000000",
	2465 => "00000000",
	2466 => "00000000",
	2467 => "00000000",
	2468 => "00000000",
	2469 => "00000000",
	2470 => "00000000",
	2471 => "00000000",
	2472 => "00000000",
	2473 => "00000000",
	2474 => "00000000",
	2475 => "00000000",
	2476 => "00000000",
	2477 => "00000000",
	2478 => "00000000",
	2479 => "00000000",
	2480 => "00000000",
	2481 => "00000000",
	2482 => "00000000",
	2483 => "00000000",
	2484 => "00000000",
	2485 => "00000000",
	2486 => "00000000",
	2487 => "00000000",
	2488 => "00000000",
	2489 => "00000000",
	2490 => "00000000",
	2491 => "00000000",
	2492 => "00000000",
	2493 => "00000000",
	2494 => "00000000",
	2495 => "00000000",
	2496 => "00000000",
	2497 => "00000000",
	2498 => "00000000",
	2499 => "00000000",
	2500 => "00000000",
	2501 => "00000000",
	2502 => "00000000",
	2503 => "00000000",
	2504 => "00000000",
	2505 => "00000000",
	2506 => "00000000",
	2507 => "00000000",
	2508 => "00000000",
	2509 => "00000000",
	2510 => "00000000",
	2511 => "00000000",
	2512 => "00000000",
	2513 => "00000000",
	2514 => "00000000",
	2515 => "00000000",
	2516 => "00000000",
	2517 => "00000000",
	2518 => "00000000",
	2519 => "00000000",
	2520 => "00000000",
	2521 => "00000000",
	2522 => "00000000",
	2523 => "00000000",
	2524 => "00000000",
	2525 => "00000000",
	2526 => "00000000",
	2527 => "00000000",
	2528 => "11111111",
	2529 => "11111111",
	2530 => "11111111",
	2531 => "11111111",
	2532 => "11111111",
	2533 => "11111111",
	2534 => "11111111",
	2535 => "11111111",
	2536 => "00000000",
	2537 => "00000000",
	2538 => "00000000",
	2539 => "00000000",
	2540 => "00000000",
	2541 => "00000000",
	2542 => "00000000",
	2543 => "00000000",
	2544 => "00000000",
	2545 => "00000000",
	2546 => "00000000",
	2547 => "00000000",
	2548 => "00000000",
	2549 => "00000000",
	2550 => "00000000",
	2551 => "00000000",
	2560 => "00000000",
	2561 => "00000000",
	2562 => "00000000",
	2563 => "00000000",
	2564 => "00000000",
	2565 => "00000000",
	2566 => "00000000",
	2567 => "00000000",
	2568 => "00000000",
	2569 => "00000000",
	2570 => "00000000",
	2571 => "00000000",
	2572 => "00000000",
	2573 => "00000000",
	2574 => "00000000",
	2575 => "00000000",
	2576 => "00000000",
	2577 => "11111111",
	2578 => "11111111",
	2579 => "11111111",
	2580 => "11111111",
	2581 => "11111111",
	2582 => "11111111",
	2583 => "11111111",
	2584 => "11111111",
	2585 => "11111111",
	2586 => "00000000",
	2587 => "00000000",
	2588 => "00000000",
	2589 => "00000000",
	2590 => "00000000",
	2591 => "00000000",
	2592 => "00000000",
	2593 => "00000000",
	2594 => "00000000",
	2595 => "00000000",
	2596 => "00000000",
	2597 => "00000000",
	2598 => "00000000",
	2599 => "00000000",
	2600 => "00000000",
	2601 => "00000000",
	2602 => "00000000",
	2603 => "00000000",
	2604 => "00000000",
	2605 => "00000000",
	2606 => "00000000",
	2607 => "00000000",
	2608 => "00000000",
	2609 => "00000000",
	2610 => "00000000",
	2611 => "00000000",
	2612 => "00000000",
	2613 => "00000000",
	2614 => "00000000",
	2615 => "00000000",
	2616 => "00000000",
	2617 => "00000000",
	2618 => "00000000",
	2619 => "00000000",
	2620 => "00000000",
	2621 => "00000000",
	2622 => "00000000",
	2623 => "00000000",
	2624 => "00000000",
	2625 => "00000000",
	2626 => "00000000",
	2627 => "00000000",
	2628 => "00000000",
	2629 => "00000000",
	2630 => "00000000",
	2631 => "00000000",
	2632 => "00000000",
	2633 => "00000000",
	2634 => "00000000",
	2635 => "00000000",
	2636 => "00000000",
	2637 => "00000000",
	2638 => "00000000",
	2639 => "00000000",
	2640 => "00000000",
	2641 => "00000000",
	2642 => "00000000",
	2643 => "00000000",
	2644 => "00000000",
	2645 => "00000000",
	2646 => "00000000",
	2647 => "00000000",
	2648 => "00000000",
	2649 => "00000000",
	2650 => "00000000",
	2651 => "00000000",
	2652 => "00000000",
	2653 => "00000000",
	2654 => "00000000",
	2655 => "11111111",
	2656 => "11111111",
	2657 => "11111111",
	2658 => "11111111",
	2659 => "11111111",
	2660 => "11111111",
	2661 => "11111111",
	2662 => "11111111",
	2663 => "11111111",
	2664 => "11111111",
	2665 => "00000000",
	2666 => "00000000",
	2667 => "00000000",
	2668 => "00000000",
	2669 => "00000000",
	2670 => "00000000",
	2671 => "00000000",
	2672 => "00000000",
	2673 => "00000000",
	2674 => "00000000",
	2675 => "00000000",
	2676 => "00000000",
	2677 => "00000000",
	2678 => "00000000",
	2679 => "00000000",
	2688 => "00000000",
	2689 => "00000000",
	2690 => "00000000",
	2691 => "00000000",
	2692 => "00000000",
	2693 => "00000000",
	2694 => "00000000",
	2695 => "00000000",
	2696 => "00000000",
	2697 => "00000000",
	2698 => "00000000",
	2699 => "00000000",
	2700 => "00000000",
	2701 => "00000000",
	2702 => "00000000",
	2703 => "00000000",
	2704 => "00000000",
	2705 => "11111111",
	2706 => "11111111",
	2707 => "11111111",
	2708 => "11111111",
	2709 => "11111111",
	2710 => "11111111",
	2711 => "11111111",
	2712 => "11111111",
	2713 => "11111111",
	2714 => "11111111",
	2715 => "00000000",
	2716 => "00000000",
	2717 => "00000000",
	2718 => "00000000",
	2719 => "00000000",
	2720 => "00000000",
	2721 => "00000000",
	2722 => "00000000",
	2723 => "00000000",
	2724 => "00000000",
	2725 => "00000000",
	2726 => "00000000",
	2727 => "00000000",
	2728 => "00000000",
	2729 => "00000000",
	2730 => "00000000",
	2731 => "00000000",
	2732 => "00000000",
	2733 => "00000000",
	2734 => "00000000",
	2735 => "00000000",
	2736 => "00000000",
	2737 => "00000000",
	2738 => "00000000",
	2739 => "00000000",
	2740 => "00000000",
	2741 => "00000000",
	2742 => "00000000",
	2743 => "00000000",
	2744 => "00000000",
	2745 => "00000000",
	2746 => "00000000",
	2747 => "00000000",
	2748 => "00000000",
	2749 => "00000000",
	2750 => "00000000",
	2751 => "00000000",
	2752 => "00000000",
	2753 => "00000000",
	2754 => "00000000",
	2755 => "00000000",
	2756 => "00000000",
	2757 => "00000000",
	2758 => "00000000",
	2759 => "00000000",
	2760 => "00000000",
	2761 => "00000000",
	2762 => "00000000",
	2763 => "00000000",
	2764 => "00000000",
	2765 => "00000000",
	2766 => "00000000",
	2767 => "00000000",
	2768 => "00000000",
	2769 => "00000000",
	2770 => "00000000",
	2771 => "00000000",
	2772 => "00000000",
	2773 => "00000000",
	2774 => "00000000",
	2775 => "00000000",
	2776 => "00000000",
	2777 => "00000000",
	2778 => "00000000",
	2779 => "00000000",
	2780 => "00000000",
	2781 => "00000000",
	2782 => "11111111",
	2783 => "11111111",
	2784 => "11111111",
	2785 => "11111111",
	2786 => "11111111",
	2787 => "11111111",
	2788 => "11111111",
	2789 => "11111111",
	2790 => "11111111",
	2791 => "11111111",
	2792 => "00000000",
	2793 => "00000000",
	2794 => "00000000",
	2795 => "00000000",
	2796 => "00000000",
	2797 => "00000000",
	2798 => "00000000",
	2799 => "00000000",
	2800 => "00000000",
	2801 => "00000000",
	2802 => "00000000",
	2803 => "00000000",
	2804 => "00000000",
	2805 => "00000000",
	2806 => "00000000",
	2807 => "00000000",
	2816 => "00000000",
	2817 => "00000000",
	2818 => "00000000",
	2819 => "00000000",
	2820 => "00000000",
	2821 => "00000000",
	2822 => "00000000",
	2823 => "00000000",
	2824 => "00000000",
	2825 => "00000000",
	2826 => "00000000",
	2827 => "00000000",
	2828 => "00000000",
	2829 => "00000000",
	2830 => "00000000",
	2831 => "00000000",
	2832 => "00000000",
	2833 => "11111111",
	2834 => "11111111",
	2835 => "11111111",
	2836 => "11111111",
	2837 => "11111111",
	2838 => "11111111",
	2839 => "11111111",
	2840 => "11111111",
	2841 => "11111111",
	2842 => "11111111",
	2843 => "11111111",
	2844 => "00000000",
	2845 => "00000000",
	2846 => "00000000",
	2847 => "00000000",
	2848 => "00000000",
	2849 => "00000000",
	2850 => "00000000",
	2851 => "00000000",
	2852 => "00000000",
	2853 => "00000000",
	2854 => "00000000",
	2855 => "00000000",
	2856 => "00000000",
	2857 => "00000000",
	2858 => "00000000",
	2859 => "00000000",
	2860 => "00000000",
	2861 => "00000000",
	2862 => "00000000",
	2863 => "00000000",
	2864 => "00000000",
	2865 => "00000000",
	2866 => "00000000",
	2867 => "00000000",
	2868 => "00000000",
	2869 => "00000000",
	2870 => "00000000",
	2871 => "00000000",
	2872 => "00000000",
	2873 => "00000000",
	2874 => "00000000",
	2875 => "00000000",
	2876 => "00000000",
	2877 => "00000000",
	2878 => "00000000",
	2879 => "00000000",
	2880 => "00000000",
	2881 => "00000000",
	2882 => "00000000",
	2883 => "00000000",
	2884 => "00000000",
	2885 => "00000000",
	2886 => "00000000",
	2887 => "00000000",
	2888 => "00000000",
	2889 => "00000000",
	2890 => "00000000",
	2891 => "00000000",
	2892 => "00000000",
	2893 => "00000000",
	2894 => "00000000",
	2895 => "00000000",
	2896 => "00000000",
	2897 => "00000000",
	2898 => "00000000",
	2899 => "00000000",
	2900 => "00000000",
	2901 => "00000000",
	2902 => "00000000",
	2903 => "00000000",
	2904 => "00000000",
	2905 => "00000000",
	2906 => "00000000",
	2907 => "00000000",
	2908 => "00000000",
	2909 => "11111111",
	2910 => "11111111",
	2911 => "11111111",
	2912 => "11111111",
	2913 => "11111111",
	2914 => "11111111",
	2915 => "11111111",
	2916 => "11111111",
	2917 => "11111111",
	2918 => "11111111",
	2919 => "11111111",
	2920 => "00000000",
	2921 => "00000000",
	2922 => "00000000",
	2923 => "00000000",
	2924 => "00000000",
	2925 => "00000000",
	2926 => "00000000",
	2927 => "00000000",
	2928 => "00000000",
	2929 => "00000000",
	2930 => "00000000",
	2931 => "00000000",
	2932 => "00000000",
	2933 => "00000000",
	2934 => "00000000",
	2935 => "00000000",
	2944 => "00000000",
	2945 => "00000000",
	2946 => "00000000",
	2947 => "00000000",
	2948 => "00000000",
	2949 => "00000000",
	2950 => "00000000",
	2951 => "00000000",
	2952 => "00000000",
	2953 => "00000000",
	2954 => "00000000",
	2955 => "00000000",
	2956 => "00000000",
	2957 => "00000000",
	2958 => "00000000",
	2959 => "00000000",
	2960 => "00000000",
	2961 => "00000000",
	2962 => "11111111",
	2963 => "11111111",
	2964 => "11111111",
	2965 => "11111111",
	2966 => "11111111",
	2967 => "11111111",
	2968 => "11111111",
	2969 => "11111111",
	2970 => "11111111",
	2971 => "11111111",
	2972 => "11111111",
	2973 => "00000000",
	2974 => "00000000",
	2975 => "00000000",
	2976 => "00000000",
	2977 => "00000000",
	2978 => "00000000",
	2979 => "00000000",
	2980 => "00000000",
	2981 => "00000000",
	2982 => "00000000",
	2983 => "00000000",
	2984 => "00000000",
	2985 => "00000000",
	2986 => "00000000",
	2987 => "00000000",
	2988 => "00000000",
	2989 => "00000000",
	2990 => "00000000",
	2991 => "00000000",
	2992 => "00000000",
	2993 => "00000000",
	2994 => "00000000",
	2995 => "00000000",
	2996 => "00000000",
	2997 => "00000000",
	2998 => "00000000",
	2999 => "00000000",
	3000 => "00000000",
	3001 => "00000000",
	3002 => "00000000",
	3003 => "00000000",
	3004 => "00000000",
	3005 => "00000000",
	3006 => "00000000",
	3007 => "00000000",
	3008 => "00000000",
	3009 => "00000000",
	3010 => "00000000",
	3011 => "00000000",
	3012 => "00000000",
	3013 => "00000000",
	3014 => "00000000",
	3015 => "00000000",
	3016 => "00000000",
	3017 => "00000000",
	3018 => "00000000",
	3019 => "00000000",
	3020 => "00000000",
	3021 => "00000000",
	3022 => "00000000",
	3023 => "00000000",
	3024 => "00000000",
	3025 => "00000000",
	3026 => "00000000",
	3027 => "00000000",
	3028 => "00000000",
	3029 => "00000000",
	3030 => "00000000",
	3031 => "00000000",
	3032 => "00000000",
	3033 => "00000000",
	3034 => "00000000",
	3035 => "00000000",
	3036 => "11111111",
	3037 => "11111111",
	3038 => "11111111",
	3039 => "11111111",
	3040 => "11111111",
	3041 => "11111111",
	3042 => "11111111",
	3043 => "11111111",
	3044 => "11111111",
	3045 => "11111111",
	3046 => "11111111",
	3047 => "00000000",
	3048 => "00000000",
	3049 => "00000000",
	3050 => "00000000",
	3051 => "00000000",
	3052 => "00000000",
	3053 => "00000000",
	3054 => "00000000",
	3055 => "00000000",
	3056 => "00000000",
	3057 => "00000000",
	3058 => "00000000",
	3059 => "00000000",
	3060 => "00000000",
	3061 => "00000000",
	3062 => "00000000",
	3063 => "00000000",
	3072 => "00000000",
	3073 => "00000000",
	3074 => "00000000",
	3075 => "00000000",
	3076 => "00000000",
	3077 => "00000000",
	3078 => "00000000",
	3079 => "00000000",
	3080 => "00000000",
	3081 => "00000000",
	3082 => "00000000",
	3083 => "00000000",
	3084 => "00000000",
	3085 => "00000000",
	3086 => "00000000",
	3087 => "00000000",
	3088 => "00000000",
	3089 => "00000000",
	3090 => "00000000",
	3091 => "11111111",
	3092 => "11111111",
	3093 => "11111111",
	3094 => "11111111",
	3095 => "11111111",
	3096 => "11111111",
	3097 => "11111111",
	3098 => "11111111",
	3099 => "11111111",
	3100 => "11111111",
	3101 => "11111111",
	3102 => "00000000",
	3103 => "00000000",
	3104 => "00000000",
	3105 => "00000000",
	3106 => "00000000",
	3107 => "00000000",
	3108 => "00000000",
	3109 => "00000000",
	3110 => "00000000",
	3111 => "00000000",
	3112 => "00000000",
	3113 => "00000000",
	3114 => "00000000",
	3115 => "00000000",
	3116 => "00000000",
	3117 => "00000000",
	3118 => "00000000",
	3119 => "00000000",
	3120 => "00000000",
	3121 => "00000000",
	3122 => "00000000",
	3123 => "00000000",
	3124 => "00000000",
	3125 => "00000000",
	3126 => "00000000",
	3127 => "00000000",
	3128 => "00000000",
	3129 => "00000000",
	3130 => "00000000",
	3131 => "00000000",
	3132 => "00000000",
	3133 => "00000000",
	3134 => "00000000",
	3135 => "00000000",
	3136 => "00000000",
	3137 => "00000000",
	3138 => "00000000",
	3139 => "00000000",
	3140 => "00000000",
	3141 => "00000000",
	3142 => "00000000",
	3143 => "00000000",
	3144 => "00000000",
	3145 => "00000000",
	3146 => "00000000",
	3147 => "00000000",
	3148 => "00000000",
	3149 => "00000000",
	3150 => "00000000",
	3151 => "00000000",
	3152 => "00000000",
	3153 => "00000000",
	3154 => "00000000",
	3155 => "00000000",
	3156 => "00000000",
	3157 => "00000000",
	3158 => "00000000",
	3159 => "00000000",
	3160 => "00000000",
	3161 => "00000000",
	3162 => "00000000",
	3163 => "11111111",
	3164 => "11111111",
	3165 => "11111111",
	3166 => "11111111",
	3167 => "11111111",
	3168 => "11111111",
	3169 => "11111111",
	3170 => "11111111",
	3171 => "11111111",
	3172 => "11111111",
	3173 => "11111111",
	3174 => "00000000",
	3175 => "00000000",
	3176 => "00000000",
	3177 => "00000000",
	3178 => "00000000",
	3179 => "00000000",
	3180 => "00000000",
	3181 => "00000000",
	3182 => "00000000",
	3183 => "00000000",
	3184 => "00000000",
	3185 => "00000000",
	3186 => "00000000",
	3187 => "00000000",
	3188 => "00000000",
	3189 => "00000000",
	3190 => "00000000",
	3191 => "00000000",
	3200 => "00000000",
	3201 => "00000000",
	3202 => "00000000",
	3203 => "00000000",
	3204 => "00000000",
	3205 => "00000000",
	3206 => "00000000",
	3207 => "00000000",
	3208 => "00000000",
	3209 => "00000000",
	3210 => "00000000",
	3211 => "00000000",
	3212 => "00000000",
	3213 => "00000000",
	3214 => "00000000",
	3215 => "00000000",
	3216 => "00000000",
	3217 => "00000000",
	3218 => "00000000",
	3219 => "00000000",
	3220 => "11111111",
	3221 => "11111111",
	3222 => "11111111",
	3223 => "11111111",
	3224 => "11111111",
	3225 => "11111111",
	3226 => "11111111",
	3227 => "11111111",
	3228 => "11111111",
	3229 => "11111111",
	3230 => "11111111",
	3231 => "00000000",
	3232 => "00000000",
	3233 => "00000000",
	3234 => "00000000",
	3235 => "00000000",
	3236 => "00000000",
	3237 => "00000000",
	3238 => "00000000",
	3239 => "00000000",
	3240 => "00000000",
	3241 => "00000000",
	3242 => "00000000",
	3243 => "00000000",
	3244 => "00000000",
	3245 => "00000000",
	3246 => "00000000",
	3247 => "00000000",
	3248 => "00000000",
	3249 => "00000000",
	3250 => "00000000",
	3251 => "00000000",
	3252 => "00000000",
	3253 => "00000000",
	3254 => "00000000",
	3255 => "00000000",
	3256 => "00000000",
	3257 => "00000000",
	3258 => "00000000",
	3259 => "00000000",
	3260 => "00000000",
	3261 => "00000000",
	3262 => "00000000",
	3263 => "00000000",
	3264 => "00000000",
	3265 => "00000000",
	3266 => "00000000",
	3267 => "00000000",
	3268 => "00000000",
	3269 => "00000000",
	3270 => "00000000",
	3271 => "00000000",
	3272 => "00000000",
	3273 => "00000000",
	3274 => "00000000",
	3275 => "00000000",
	3276 => "00000000",
	3277 => "00000000",
	3278 => "00000000",
	3279 => "00000000",
	3280 => "00000000",
	3281 => "00000000",
	3282 => "00000000",
	3283 => "00000000",
	3284 => "00000000",
	3285 => "00000000",
	3286 => "00000000",
	3287 => "00000000",
	3288 => "00000000",
	3289 => "00000000",
	3290 => "11111111",
	3291 => "11111111",
	3292 => "11111111",
	3293 => "11111111",
	3294 => "11111111",
	3295 => "11111111",
	3296 => "11111111",
	3297 => "11111111",
	3298 => "11111111",
	3299 => "11111111",
	3300 => "11111111",
	3301 => "00000000",
	3302 => "00000000",
	3303 => "00000000",
	3304 => "00000000",
	3305 => "00000000",
	3306 => "00000000",
	3307 => "00000000",
	3308 => "00000000",
	3309 => "00000000",
	3310 => "00000000",
	3311 => "00000000",
	3312 => "00000000",
	3313 => "00000000",
	3314 => "00000000",
	3315 => "00000000",
	3316 => "00000000",
	3317 => "00000000",
	3318 => "00000000",
	3319 => "00000000",
	3328 => "00000000",
	3329 => "00000000",
	3330 => "00000000",
	3331 => "00000000",
	3332 => "00000000",
	3333 => "00000000",
	3334 => "00000000",
	3335 => "00000000",
	3336 => "00000000",
	3337 => "00000000",
	3338 => "00000000",
	3339 => "00000000",
	3340 => "00000000",
	3341 => "00000000",
	3342 => "00000000",
	3343 => "00000000",
	3344 => "00000000",
	3345 => "00000000",
	3346 => "00000000",
	3347 => "00000000",
	3348 => "00000000",
	3349 => "11111111",
	3350 => "11111111",
	3351 => "11111111",
	3352 => "11111111",
	3353 => "11111111",
	3354 => "11111111",
	3355 => "11111111",
	3356 => "11111111",
	3357 => "11111111",
	3358 => "11111111",
	3359 => "11111111",
	3360 => "00000000",
	3361 => "00000000",
	3362 => "00000000",
	3363 => "00000000",
	3364 => "00000000",
	3365 => "00000000",
	3366 => "00000000",
	3367 => "00000000",
	3368 => "00000000",
	3369 => "00000000",
	3370 => "00000000",
	3371 => "00000000",
	3372 => "00000000",
	3373 => "00000000",
	3374 => "00000000",
	3375 => "00000000",
	3376 => "00000000",
	3377 => "00000000",
	3378 => "00000000",
	3379 => "00000000",
	3380 => "00000000",
	3381 => "00000000",
	3382 => "00000000",
	3383 => "00000000",
	3384 => "00000000",
	3385 => "00000000",
	3386 => "00000000",
	3387 => "00000000",
	3388 => "00000000",
	3389 => "00000000",
	3390 => "00000000",
	3391 => "00000000",
	3392 => "00000000",
	3393 => "00000000",
	3394 => "00000000",
	3395 => "00000000",
	3396 => "00000000",
	3397 => "00000000",
	3398 => "00000000",
	3399 => "00000000",
	3400 => "00000000",
	3401 => "00000000",
	3402 => "00000000",
	3403 => "00000000",
	3404 => "00000000",
	3405 => "00000000",
	3406 => "00000000",
	3407 => "00000000",
	3408 => "00000000",
	3409 => "00000000",
	3410 => "00000000",
	3411 => "00000000",
	3412 => "00000000",
	3413 => "00000000",
	3414 => "00000000",
	3415 => "00000000",
	3416 => "00000000",
	3417 => "11111111",
	3418 => "11111111",
	3419 => "11111111",
	3420 => "11111111",
	3421 => "11111111",
	3422 => "11111111",
	3423 => "11111111",
	3424 => "11111111",
	3425 => "11111111",
	3426 => "11111111",
	3427 => "11111111",
	3428 => "00000000",
	3429 => "00000000",
	3430 => "00000000",
	3431 => "00000000",
	3432 => "00000000",
	3433 => "00000000",
	3434 => "00000000",
	3435 => "00000000",
	3436 => "00000000",
	3437 => "00000000",
	3438 => "00000000",
	3439 => "00000000",
	3440 => "00000000",
	3441 => "00000000",
	3442 => "00000000",
	3443 => "00000000",
	3444 => "00000000",
	3445 => "00000000",
	3446 => "00000000",
	3447 => "00000000",
	3456 => "00000000",
	3457 => "00000000",
	3458 => "00000000",
	3459 => "00000000",
	3460 => "00000000",
	3461 => "00000000",
	3462 => "00000000",
	3463 => "00000000",
	3464 => "00000000",
	3465 => "00000000",
	3466 => "00000000",
	3467 => "00000000",
	3468 => "00000000",
	3469 => "00000000",
	3470 => "00000000",
	3471 => "00000000",
	3472 => "00000000",
	3473 => "00000000",
	3474 => "00000000",
	3475 => "00000000",
	3476 => "00000000",
	3477 => "00000000",
	3478 => "11111111",
	3479 => "11111111",
	3480 => "11111111",
	3481 => "11111111",
	3482 => "11111111",
	3483 => "11111111",
	3484 => "11111111",
	3485 => "11111111",
	3486 => "11111111",
	3487 => "11111111",
	3488 => "11111111",
	3489 => "00000000",
	3490 => "00000000",
	3491 => "00000000",
	3492 => "00000000",
	3493 => "00000000",
	3494 => "00000000",
	3495 => "00000000",
	3496 => "00000000",
	3497 => "00000000",
	3498 => "00000000",
	3499 => "00000000",
	3500 => "00000000",
	3501 => "00000000",
	3502 => "00000000",
	3503 => "00000000",
	3504 => "00000000",
	3505 => "00000000",
	3506 => "00000000",
	3507 => "00000000",
	3508 => "00000000",
	3509 => "00000000",
	3510 => "00000000",
	3511 => "00000000",
	3512 => "00000000",
	3513 => "00000000",
	3514 => "00000000",
	3515 => "00000000",
	3516 => "00000000",
	3517 => "00000000",
	3518 => "00000000",
	3519 => "00000000",
	3520 => "00000000",
	3521 => "00000000",
	3522 => "00000000",
	3523 => "00000000",
	3524 => "00000000",
	3525 => "00000000",
	3526 => "00000000",
	3527 => "00000000",
	3528 => "00000000",
	3529 => "00000000",
	3530 => "00000000",
	3531 => "00000000",
	3532 => "00000000",
	3533 => "00000000",
	3534 => "00000000",
	3535 => "00000000",
	3536 => "00000000",
	3537 => "00000000",
	3538 => "00000000",
	3539 => "00000000",
	3540 => "00000000",
	3541 => "00000000",
	3542 => "00000000",
	3543 => "00000000",
	3544 => "11111111",
	3545 => "11111111",
	3546 => "11111111",
	3547 => "11111111",
	3548 => "11111111",
	3549 => "11111111",
	3550 => "11111111",
	3551 => "11111111",
	3552 => "11111111",
	3553 => "11111111",
	3554 => "11111111",
	3555 => "00000000",
	3556 => "00000000",
	3557 => "00000000",
	3558 => "00000000",
	3559 => "00000000",
	3560 => "00000000",
	3561 => "00000000",
	3562 => "00000000",
	3563 => "00000000",
	3564 => "00000000",
	3565 => "00000000",
	3566 => "00000000",
	3567 => "00000000",
	3568 => "00000000",
	3569 => "00000000",
	3570 => "00000000",
	3571 => "00000000",
	3572 => "00000000",
	3573 => "00000000",
	3574 => "00000000",
	3575 => "00000000",
	3584 => "00000000",
	3585 => "00000000",
	3586 => "00000000",
	3587 => "00000000",
	3588 => "00000000",
	3589 => "00000000",
	3590 => "00000000",
	3591 => "00000000",
	3592 => "00000000",
	3593 => "00000000",
	3594 => "00000000",
	3595 => "00000000",
	3596 => "00000000",
	3597 => "00000000",
	3598 => "00000000",
	3599 => "00000000",
	3600 => "00000000",
	3601 => "00000000",
	3602 => "00000000",
	3603 => "00000000",
	3604 => "00000000",
	3605 => "00000000",
	3606 => "00000000",
	3607 => "11111111",
	3608 => "11111111",
	3609 => "11111111",
	3610 => "11111111",
	3611 => "11111111",
	3612 => "11111111",
	3613 => "11111111",
	3614 => "11111111",
	3615 => "11111111",
	3616 => "11111111",
	3617 => "11111111",
	3618 => "00000000",
	3619 => "00000000",
	3620 => "00000000",
	3621 => "00000000",
	3622 => "00000000",
	3623 => "00000000",
	3624 => "00000000",
	3625 => "00000000",
	3626 => "00000000",
	3627 => "00000000",
	3628 => "00000000",
	3629 => "00000000",
	3630 => "00000000",
	3631 => "00000000",
	3632 => "00000000",
	3633 => "00000000",
	3634 => "00000000",
	3635 => "00000000",
	3636 => "00000000",
	3637 => "00000000",
	3638 => "00000000",
	3639 => "00000000",
	3640 => "00000000",
	3641 => "00000000",
	3642 => "00000000",
	3643 => "00000000",
	3644 => "00000000",
	3645 => "00000000",
	3646 => "00000000",
	3647 => "00000000",
	3648 => "00000000",
	3649 => "00000000",
	3650 => "00000000",
	3651 => "00000000",
	3652 => "00000000",
	3653 => "00000000",
	3654 => "00000000",
	3655 => "00000000",
	3656 => "00000000",
	3657 => "00000000",
	3658 => "00000000",
	3659 => "00000000",
	3660 => "00000000",
	3661 => "00000000",
	3662 => "00000000",
	3663 => "00000000",
	3664 => "00000000",
	3665 => "00000000",
	3666 => "00000000",
	3667 => "00000000",
	3668 => "00000000",
	3669 => "00000000",
	3670 => "00000000",
	3671 => "11111111",
	3672 => "11111111",
	3673 => "11111111",
	3674 => "11111111",
	3675 => "11111111",
	3676 => "11111111",
	3677 => "11111111",
	3678 => "11111111",
	3679 => "11111111",
	3680 => "11111111",
	3681 => "11111111",
	3682 => "00000000",
	3683 => "00000000",
	3684 => "00000000",
	3685 => "00000000",
	3686 => "00000000",
	3687 => "00000000",
	3688 => "00000000",
	3689 => "00000000",
	3690 => "00000000",
	3691 => "00000000",
	3692 => "00000000",
	3693 => "00000000",
	3694 => "00000000",
	3695 => "00000000",
	3696 => "00000000",
	3697 => "00000000",
	3698 => "00000000",
	3699 => "00000000",
	3700 => "00000000",
	3701 => "00000000",
	3702 => "00000000",
	3703 => "00000000",
	3712 => "00000000",
	3713 => "00000000",
	3714 => "00000000",
	3715 => "00000000",
	3716 => "00000000",
	3717 => "00000000",
	3718 => "00000000",
	3719 => "00000000",
	3720 => "00000000",
	3721 => "00000000",
	3722 => "00000000",
	3723 => "00000000",
	3724 => "00000000",
	3725 => "00000000",
	3726 => "00000000",
	3727 => "00000000",
	3728 => "00000000",
	3729 => "00000000",
	3730 => "00000000",
	3731 => "00000000",
	3732 => "00000000",
	3733 => "00000000",
	3734 => "00000000",
	3735 => "00000000",
	3736 => "11111111",
	3737 => "11111111",
	3738 => "11111111",
	3739 => "11111111",
	3740 => "11111111",
	3741 => "11111111",
	3742 => "11111111",
	3743 => "11111111",
	3744 => "11111111",
	3745 => "11111111",
	3746 => "11111111",
	3747 => "00000000",
	3748 => "00000000",
	3749 => "00000000",
	3750 => "00000000",
	3751 => "00000000",
	3752 => "00000000",
	3753 => "00000000",
	3754 => "00000000",
	3755 => "00000000",
	3756 => "00000000",
	3757 => "00000000",
	3758 => "00000000",
	3759 => "00000000",
	3760 => "00000000",
	3761 => "00000000",
	3762 => "00000000",
	3763 => "00000000",
	3764 => "00000000",
	3765 => "00000000",
	3766 => "00000000",
	3767 => "00000000",
	3768 => "00000000",
	3769 => "00000000",
	3770 => "00000000",
	3771 => "00000000",
	3772 => "00000000",
	3773 => "00000000",
	3774 => "00000000",
	3775 => "00000000",
	3776 => "00000000",
	3777 => "00000000",
	3778 => "00000000",
	3779 => "00000000",
	3780 => "00000000",
	3781 => "00000000",
	3782 => "00000000",
	3783 => "00000000",
	3784 => "00000000",
	3785 => "00000000",
	3786 => "00000000",
	3787 => "00000000",
	3788 => "00000000",
	3789 => "00000000",
	3790 => "00000000",
	3791 => "00000000",
	3792 => "00000000",
	3793 => "00000000",
	3794 => "00000000",
	3795 => "00000000",
	3796 => "00000000",
	3797 => "00000000",
	3798 => "11111111",
	3799 => "11111111",
	3800 => "11111111",
	3801 => "11111111",
	3802 => "11111111",
	3803 => "11111111",
	3804 => "11111111",
	3805 => "11111111",
	3806 => "11111111",
	3807 => "11111111",
	3808 => "11111111",
	3809 => "00000000",
	3810 => "00000000",
	3811 => "00000000",
	3812 => "00000000",
	3813 => "00000000",
	3814 => "00000000",
	3815 => "00000000",
	3816 => "00000000",
	3817 => "00000000",
	3818 => "00000000",
	3819 => "00000000",
	3820 => "00000000",
	3821 => "00000000",
	3822 => "00000000",
	3823 => "00000000",
	3824 => "00000000",
	3825 => "00000000",
	3826 => "00000000",
	3827 => "00000000",
	3828 => "00000000",
	3829 => "00000000",
	3830 => "00000000",
	3831 => "00000000",
	3840 => "00000000",
	3841 => "00000000",
	3842 => "00000000",
	3843 => "00000000",
	3844 => "00000000",
	3845 => "00000000",
	3846 => "00000000",
	3847 => "00000000",
	3848 => "00000000",
	3849 => "00000000",
	3850 => "00000000",
	3851 => "00000000",
	3852 => "00000000",
	3853 => "00000000",
	3854 => "00000000",
	3855 => "00000000",
	3856 => "00000000",
	3857 => "00000000",
	3858 => "00000000",
	3859 => "00000000",
	3860 => "00000000",
	3861 => "00000000",
	3862 => "00000000",
	3863 => "00000000",
	3864 => "00000000",
	3865 => "11111111",
	3866 => "11111111",
	3867 => "11111111",
	3868 => "11111111",
	3869 => "11111111",
	3870 => "11111111",
	3871 => "11111111",
	3872 => "11111111",
	3873 => "11111111",
	3874 => "11111111",
	3875 => "11111111",
	3876 => "00000000",
	3877 => "00000000",
	3878 => "00000000",
	3879 => "00000000",
	3880 => "00000000",
	3881 => "00000000",
	3882 => "00000000",
	3883 => "00000000",
	3884 => "00000000",
	3885 => "00000000",
	3886 => "00000000",
	3887 => "00000000",
	3888 => "00000000",
	3889 => "00000000",
	3890 => "00000000",
	3891 => "00000000",
	3892 => "00000000",
	3893 => "00000000",
	3894 => "00000000",
	3895 => "00000000",
	3896 => "00000000",
	3897 => "00000000",
	3898 => "00000000",
	3899 => "00000000",
	3900 => "00000000",
	3901 => "00000000",
	3902 => "00000000",
	3903 => "00000000",
	3904 => "00000000",
	3905 => "00000000",
	3906 => "00000000",
	3907 => "00000000",
	3908 => "00000000",
	3909 => "00000000",
	3910 => "00000000",
	3911 => "00000000",
	3912 => "00000000",
	3913 => "00000000",
	3914 => "00000000",
	3915 => "00000000",
	3916 => "00000000",
	3917 => "00000000",
	3918 => "00000000",
	3919 => "00000000",
	3920 => "00000000",
	3921 => "00000000",
	3922 => "00000000",
	3923 => "00000000",
	3924 => "00000000",
	3925 => "11111111",
	3926 => "11111111",
	3927 => "11111111",
	3928 => "11111111",
	3929 => "11111111",
	3930 => "11111111",
	3931 => "11111111",
	3932 => "11111111",
	3933 => "11111111",
	3934 => "11111111",
	3935 => "11111111",
	3936 => "00000000",
	3937 => "00000000",
	3938 => "00000000",
	3939 => "00000000",
	3940 => "00000000",
	3941 => "00000000",
	3942 => "00000000",
	3943 => "00000000",
	3944 => "00000000",
	3945 => "00000000",
	3946 => "00000000",
	3947 => "00000000",
	3948 => "00000000",
	3949 => "00000000",
	3950 => "00000000",
	3951 => "00000000",
	3952 => "00000000",
	3953 => "00000000",
	3954 => "00000000",
	3955 => "00000000",
	3956 => "00000000",
	3957 => "00000000",
	3958 => "00000000",
	3959 => "00000000",
	3968 => "00000000",
	3969 => "00000000",
	3970 => "00000000",
	3971 => "00000000",
	3972 => "00000000",
	3973 => "00000000",
	3974 => "00000000",
	3975 => "00000000",
	3976 => "00000000",
	3977 => "00000000",
	3978 => "00000000",
	3979 => "00000000",
	3980 => "00000000",
	3981 => "00000000",
	3982 => "00000000",
	3983 => "00000000",
	3984 => "00000000",
	3985 => "00000000",
	3986 => "00000000",
	3987 => "00000000",
	3988 => "00000000",
	3989 => "00000000",
	3990 => "00000000",
	3991 => "00000000",
	3992 => "00000000",
	3993 => "00000000",
	3994 => "11111111",
	3995 => "11111111",
	3996 => "11111111",
	3997 => "11111111",
	3998 => "11111111",
	3999 => "11111111",
	4000 => "11111111",
	4001 => "11111111",
	4002 => "11111111",
	4003 => "11111111",
	4004 => "11111111",
	4005 => "00000000",
	4006 => "00000000",
	4007 => "00000000",
	4008 => "00000000",
	4009 => "00000000",
	4010 => "00000000",
	4011 => "00000000",
	4012 => "00000000",
	4013 => "00000000",
	4014 => "00000000",
	4015 => "00000000",
	4016 => "00000000",
	4017 => "00000000",
	4018 => "00000000",
	4019 => "00000000",
	4020 => "00000000",
	4021 => "00000000",
	4022 => "00000000",
	4023 => "00000000",
	4024 => "00000000",
	4025 => "00000000",
	4026 => "00000000",
	4027 => "00000000",
	4028 => "00000000",
	4029 => "00000000",
	4030 => "00000000",
	4031 => "00000000",
	4032 => "00000000",
	4033 => "00000000",
	4034 => "00000000",
	4035 => "00000000",
	4036 => "00000000",
	4037 => "00000000",
	4038 => "00000000",
	4039 => "00000000",
	4040 => "00000000",
	4041 => "00000000",
	4042 => "00000000",
	4043 => "00000000",
	4044 => "00000000",
	4045 => "00000000",
	4046 => "00000000",
	4047 => "00000000",
	4048 => "00000000",
	4049 => "00000000",
	4050 => "00000000",
	4051 => "00000000",
	4052 => "11111111",
	4053 => "11111111",
	4054 => "11111111",
	4055 => "11111111",
	4056 => "11111111",
	4057 => "11111111",
	4058 => "11111111",
	4059 => "11111111",
	4060 => "11111111",
	4061 => "11111111",
	4062 => "11111111",
	4063 => "00000000",
	4064 => "00000000",
	4065 => "00000000",
	4066 => "00000000",
	4067 => "00000000",
	4068 => "00000000",
	4069 => "00000000",
	4070 => "00000000",
	4071 => "00000000",
	4072 => "00000000",
	4073 => "00000000",
	4074 => "00000000",
	4075 => "00000000",
	4076 => "00000000",
	4077 => "00000000",
	4078 => "00000000",
	4079 => "00000000",
	4080 => "00000000",
	4081 => "00000000",
	4082 => "00000000",
	4083 => "00000000",
	4084 => "00000000",
	4085 => "00000000",
	4086 => "00000000",
	4087 => "00000000",
	4096 => "00000000",
	4097 => "00000000",
	4098 => "00000000",
	4099 => "00000000",
	4100 => "00000000",
	4101 => "00000000",
	4102 => "00000000",
	4103 => "00000000",
	4104 => "00000000",
	4105 => "00000000",
	4106 => "00000000",
	4107 => "00000000",
	4108 => "00000000",
	4109 => "00000000",
	4110 => "00000000",
	4111 => "00000000",
	4112 => "00000000",
	4113 => "00000000",
	4114 => "00000000",
	4115 => "00000000",
	4116 => "00000000",
	4117 => "00000000",
	4118 => "00000000",
	4119 => "00000000",
	4120 => "00000000",
	4121 => "00000000",
	4122 => "00000000",
	4123 => "11111111",
	4124 => "11111111",
	4125 => "11111111",
	4126 => "11111111",
	4127 => "11111111",
	4128 => "11111111",
	4129 => "11111111",
	4130 => "11111111",
	4131 => "11111111",
	4132 => "11111111",
	4133 => "11111111",
	4134 => "00000000",
	4135 => "00000000",
	4136 => "00000000",
	4137 => "00000000",
	4138 => "00000000",
	4139 => "00000000",
	4140 => "00000000",
	4141 => "00000000",
	4142 => "00000000",
	4143 => "00000000",
	4144 => "00000000",
	4145 => "00000000",
	4146 => "00000000",
	4147 => "00000000",
	4148 => "00000000",
	4149 => "00000000",
	4150 => "00000000",
	4151 => "00000000",
	4152 => "00000000",
	4153 => "00000000",
	4154 => "00000000",
	4155 => "00000000",
	4156 => "00000000",
	4157 => "00000000",
	4158 => "00000000",
	4159 => "00000000",
	4160 => "00000000",
	4161 => "00000000",
	4162 => "00000000",
	4163 => "00000000",
	4164 => "00000000",
	4165 => "00000000",
	4166 => "00000000",
	4167 => "00000000",
	4168 => "00000000",
	4169 => "00000000",
	4170 => "00000000",
	4171 => "00000000",
	4172 => "00000000",
	4173 => "00000000",
	4174 => "00000000",
	4175 => "00000000",
	4176 => "00000000",
	4177 => "00000000",
	4178 => "00000000",
	4179 => "11111111",
	4180 => "11111111",
	4181 => "11111111",
	4182 => "11111111",
	4183 => "11111111",
	4184 => "11111111",
	4185 => "11111111",
	4186 => "11111111",
	4187 => "11111111",
	4188 => "11111111",
	4189 => "11111111",
	4190 => "00000000",
	4191 => "00000000",
	4192 => "00000000",
	4193 => "00000000",
	4194 => "00000000",
	4195 => "00000000",
	4196 => "00000000",
	4197 => "00000000",
	4198 => "00000000",
	4199 => "00000000",
	4200 => "00000000",
	4201 => "00000000",
	4202 => "00000000",
	4203 => "00000000",
	4204 => "00000000",
	4205 => "00000000",
	4206 => "00000000",
	4207 => "00000000",
	4208 => "00000000",
	4209 => "00000000",
	4210 => "00000000",
	4211 => "00000000",
	4212 => "00000000",
	4213 => "00000000",
	4214 => "00000000",
	4215 => "00000000",
	4224 => "00000000",
	4225 => "00000000",
	4226 => "00000000",
	4227 => "00000000",
	4228 => "00000000",
	4229 => "00000000",
	4230 => "00000000",
	4231 => "00000000",
	4232 => "00000000",
	4233 => "00000000",
	4234 => "00000000",
	4235 => "00000000",
	4236 => "00000000",
	4237 => "00000000",
	4238 => "00000000",
	4239 => "00000000",
	4240 => "00000000",
	4241 => "00000000",
	4242 => "00000000",
	4243 => "00000000",
	4244 => "00000000",
	4245 => "00000000",
	4246 => "00000000",
	4247 => "00000000",
	4248 => "00000000",
	4249 => "00000000",
	4250 => "00000000",
	4251 => "00000000",
	4252 => "11111111",
	4253 => "11111111",
	4254 => "11111111",
	4255 => "11111111",
	4256 => "11111111",
	4257 => "11111111",
	4258 => "11111111",
	4259 => "11111111",
	4260 => "11111111",
	4261 => "11111111",
	4262 => "11111111",
	4263 => "00000000",
	4264 => "00000000",
	4265 => "00000000",
	4266 => "00000000",
	4267 => "00000000",
	4268 => "00000000",
	4269 => "00000000",
	4270 => "00000000",
	4271 => "00000000",
	4272 => "00000000",
	4273 => "00000000",
	4274 => "00000000",
	4275 => "00000000",
	4276 => "00000000",
	4277 => "00000000",
	4278 => "00000000",
	4279 => "00000000",
	4280 => "00000000",
	4281 => "00000000",
	4282 => "00000000",
	4283 => "00000000",
	4284 => "00000000",
	4285 => "00000000",
	4286 => "00000000",
	4287 => "00000000",
	4288 => "00000000",
	4289 => "00000000",
	4290 => "00000000",
	4291 => "00000000",
	4292 => "00000000",
	4293 => "00000000",
	4294 => "00000000",
	4295 => "00000000",
	4296 => "00000000",
	4297 => "00000000",
	4298 => "00000000",
	4299 => "00000000",
	4300 => "00000000",
	4301 => "00000000",
	4302 => "00000000",
	4303 => "00000000",
	4304 => "00000000",
	4305 => "00000000",
	4306 => "11111111",
	4307 => "11111111",
	4308 => "11111111",
	4309 => "11111111",
	4310 => "11111111",
	4311 => "11111111",
	4312 => "11111111",
	4313 => "11111111",
	4314 => "11111111",
	4315 => "11111111",
	4316 => "11111111",
	4317 => "00000000",
	4318 => "00000000",
	4319 => "00000000",
	4320 => "00000000",
	4321 => "00000000",
	4322 => "00000000",
	4323 => "00000000",
	4324 => "00000000",
	4325 => "00000000",
	4326 => "00000000",
	4327 => "00000000",
	4328 => "00000000",
	4329 => "00000000",
	4330 => "00000000",
	4331 => "00000000",
	4332 => "00000000",
	4333 => "00000000",
	4334 => "00000000",
	4335 => "00000000",
	4336 => "00000000",
	4337 => "00000000",
	4338 => "00000000",
	4339 => "00000000",
	4340 => "00000000",
	4341 => "00000000",
	4342 => "00000000",
	4343 => "00000000",
	4352 => "00000000",
	4353 => "00000000",
	4354 => "00000000",
	4355 => "00000000",
	4356 => "00000000",
	4357 => "00000000",
	4358 => "00000000",
	4359 => "00000000",
	4360 => "00000000",
	4361 => "00000000",
	4362 => "00000000",
	4363 => "00000000",
	4364 => "00000000",
	4365 => "00000000",
	4366 => "00000000",
	4367 => "00000000",
	4368 => "00000000",
	4369 => "00000000",
	4370 => "00000000",
	4371 => "00000000",
	4372 => "00000000",
	4373 => "00000000",
	4374 => "00000000",
	4375 => "00000000",
	4376 => "00000000",
	4377 => "00000000",
	4378 => "00000000",
	4379 => "00000000",
	4380 => "00000000",
	4381 => "11111111",
	4382 => "11111111",
	4383 => "11111111",
	4384 => "11111111",
	4385 => "11111111",
	4386 => "11111111",
	4387 => "11111111",
	4388 => "11111111",
	4389 => "11111111",
	4390 => "11111111",
	4391 => "11111111",
	4392 => "00000000",
	4393 => "00000000",
	4394 => "00000000",
	4395 => "00000000",
	4396 => "00000000",
	4397 => "00000000",
	4398 => "00000000",
	4399 => "00000000",
	4400 => "00000000",
	4401 => "00000000",
	4402 => "00000000",
	4403 => "00000000",
	4404 => "00000000",
	4405 => "00000000",
	4406 => "00000000",
	4407 => "00000000",
	4408 => "00000000",
	4409 => "00000000",
	4410 => "00000000",
	4411 => "00000000",
	4412 => "00000000",
	4413 => "00000000",
	4414 => "00000000",
	4415 => "00000000",
	4416 => "00000000",
	4417 => "00000000",
	4418 => "00000000",
	4419 => "00000000",
	4420 => "00000000",
	4421 => "00000000",
	4422 => "00000000",
	4423 => "00000000",
	4424 => "00000000",
	4425 => "00000000",
	4426 => "00000000",
	4427 => "00000000",
	4428 => "00000000",
	4429 => "00000000",
	4430 => "00000000",
	4431 => "00000000",
	4432 => "00000000",
	4433 => "11111111",
	4434 => "11111111",
	4435 => "11111111",
	4436 => "11111111",
	4437 => "11111111",
	4438 => "11111111",
	4439 => "11111111",
	4440 => "11111111",
	4441 => "11111111",
	4442 => "11111111",
	4443 => "11111111",
	4444 => "00000000",
	4445 => "00000000",
	4446 => "00000000",
	4447 => "00000000",
	4448 => "00000000",
	4449 => "00000000",
	4450 => "00000000",
	4451 => "00000000",
	4452 => "00000000",
	4453 => "00000000",
	4454 => "00000000",
	4455 => "00000000",
	4456 => "00000000",
	4457 => "00000000",
	4458 => "00000000",
	4459 => "00000000",
	4460 => "00000000",
	4461 => "00000000",
	4462 => "00000000",
	4463 => "00000000",
	4464 => "00000000",
	4465 => "00000000",
	4466 => "00000000",
	4467 => "00000000",
	4468 => "00000000",
	4469 => "00000000",
	4470 => "00000000",
	4471 => "00000000",
	4480 => "00000000",
	4481 => "00000000",
	4482 => "00000000",
	4483 => "00000000",
	4484 => "00000000",
	4485 => "00000000",
	4486 => "00000000",
	4487 => "00000000",
	4488 => "00000000",
	4489 => "00000000",
	4490 => "00000000",
	4491 => "00000000",
	4492 => "00000000",
	4493 => "00000000",
	4494 => "00000000",
	4495 => "00000000",
	4496 => "00000000",
	4497 => "00000000",
	4498 => "00000000",
	4499 => "00000000",
	4500 => "00000000",
	4501 => "00000000",
	4502 => "00000000",
	4503 => "00000000",
	4504 => "00000000",
	4505 => "00000000",
	4506 => "00000000",
	4507 => "00000000",
	4508 => "00000000",
	4509 => "00000000",
	4510 => "11111111",
	4511 => "11111111",
	4512 => "11111111",
	4513 => "11111111",
	4514 => "11111111",
	4515 => "11111111",
	4516 => "11111111",
	4517 => "11111111",
	4518 => "11111111",
	4519 => "11111111",
	4520 => "11111111",
	4521 => "00000000",
	4522 => "00000000",
	4523 => "00000000",
	4524 => "00000000",
	4525 => "00000000",
	4526 => "00000000",
	4527 => "00000000",
	4528 => "00000000",
	4529 => "00000000",
	4530 => "00000000",
	4531 => "00000000",
	4532 => "00000000",
	4533 => "00000000",
	4534 => "00000000",
	4535 => "00000000",
	4536 => "00000000",
	4537 => "00000000",
	4538 => "00000000",
	4539 => "00000000",
	4540 => "00000000",
	4541 => "00000000",
	4542 => "00000000",
	4543 => "00000000",
	4544 => "00000000",
	4545 => "00000000",
	4546 => "00000000",
	4547 => "00000000",
	4548 => "00000000",
	4549 => "00000000",
	4550 => "00000000",
	4551 => "00000000",
	4552 => "00000000",
	4553 => "00000000",
	4554 => "00000000",
	4555 => "00000000",
	4556 => "00000000",
	4557 => "00000000",
	4558 => "00000000",
	4559 => "00000000",
	4560 => "11111111",
	4561 => "11111111",
	4562 => "11111111",
	4563 => "11111111",
	4564 => "11111111",
	4565 => "11111111",
	4566 => "11111111",
	4567 => "11111111",
	4568 => "11111111",
	4569 => "11111111",
	4570 => "11111111",
	4571 => "00000000",
	4572 => "00000000",
	4573 => "00000000",
	4574 => "00000000",
	4575 => "00000000",
	4576 => "00000000",
	4577 => "00000000",
	4578 => "00000000",
	4579 => "00000000",
	4580 => "00000000",
	4581 => "00000000",
	4582 => "00000000",
	4583 => "00000000",
	4584 => "00000000",
	4585 => "00000000",
	4586 => "00000000",
	4587 => "00000000",
	4588 => "00000000",
	4589 => "00000000",
	4590 => "00000000",
	4591 => "00000000",
	4592 => "00000000",
	4593 => "00000000",
	4594 => "00000000",
	4595 => "00000000",
	4596 => "00000000",
	4597 => "00000000",
	4598 => "00000000",
	4599 => "00000000",
	4608 => "00000000",
	4609 => "00000000",
	4610 => "00000000",
	4611 => "00000000",
	4612 => "00000000",
	4613 => "00000000",
	4614 => "00000000",
	4615 => "00000000",
	4616 => "00000000",
	4617 => "00000000",
	4618 => "00000000",
	4619 => "00000000",
	4620 => "00000000",
	4621 => "00000000",
	4622 => "00000000",
	4623 => "00000000",
	4624 => "00000000",
	4625 => "00000000",
	4626 => "00000000",
	4627 => "00000000",
	4628 => "00000000",
	4629 => "00000000",
	4630 => "00000000",
	4631 => "00000000",
	4632 => "00000000",
	4633 => "00000000",
	4634 => "00000000",
	4635 => "00000000",
	4636 => "00000000",
	4637 => "00000000",
	4638 => "00000000",
	4639 => "11111111",
	4640 => "11111111",
	4641 => "11111111",
	4642 => "11111111",
	4643 => "11111111",
	4644 => "11111111",
	4645 => "11111111",
	4646 => "11111111",
	4647 => "11111111",
	4648 => "11111111",
	4649 => "11111111",
	4650 => "00000000",
	4651 => "00000000",
	4652 => "00000000",
	4653 => "00000000",
	4654 => "00000000",
	4655 => "00000000",
	4656 => "00000000",
	4657 => "00000000",
	4658 => "00000000",
	4659 => "00000000",
	4660 => "00000000",
	4661 => "00000000",
	4662 => "00000000",
	4663 => "00000000",
	4664 => "00000000",
	4665 => "00000000",
	4666 => "00000000",
	4667 => "00000000",
	4668 => "00000000",
	4669 => "00000000",
	4670 => "00000000",
	4671 => "00000000",
	4672 => "00000000",
	4673 => "00000000",
	4674 => "00000000",
	4675 => "00000000",
	4676 => "00000000",
	4677 => "00000000",
	4678 => "00000000",
	4679 => "00000000",
	4680 => "00000000",
	4681 => "00000000",
	4682 => "00000000",
	4683 => "00000000",
	4684 => "00000000",
	4685 => "00000000",
	4686 => "00000000",
	4687 => "11111111",
	4688 => "11111111",
	4689 => "11111111",
	4690 => "11111111",
	4691 => "11111111",
	4692 => "11111111",
	4693 => "11111111",
	4694 => "11111111",
	4695 => "11111111",
	4696 => "11111111",
	4697 => "11111111",
	4698 => "00000000",
	4699 => "00000000",
	4700 => "00000000",
	4701 => "00000000",
	4702 => "00000000",
	4703 => "00000000",
	4704 => "00000000",
	4705 => "00000000",
	4706 => "00000000",
	4707 => "00000000",
	4708 => "00000000",
	4709 => "00000000",
	4710 => "00000000",
	4711 => "00000000",
	4712 => "00000000",
	4713 => "00000000",
	4714 => "00000000",
	4715 => "00000000",
	4716 => "00000000",
	4717 => "00000000",
	4718 => "00000000",
	4719 => "00000000",
	4720 => "00000000",
	4721 => "00000000",
	4722 => "00000000",
	4723 => "00000000",
	4724 => "00000000",
	4725 => "00000000",
	4726 => "00000000",
	4727 => "00000000",
	4736 => "00000000",
	4737 => "00000000",
	4738 => "00000000",
	4739 => "00000000",
	4740 => "00000000",
	4741 => "00000000",
	4742 => "00000000",
	4743 => "00000000",
	4744 => "00000000",
	4745 => "00000000",
	4746 => "00000000",
	4747 => "00000000",
	4748 => "00000000",
	4749 => "00000000",
	4750 => "00000000",
	4751 => "00000000",
	4752 => "00000000",
	4753 => "00000000",
	4754 => "00000000",
	4755 => "00000000",
	4756 => "00000000",
	4757 => "00000000",
	4758 => "00000000",
	4759 => "00000000",
	4760 => "00000000",
	4761 => "00000000",
	4762 => "00000000",
	4763 => "00000000",
	4764 => "00000000",
	4765 => "00000000",
	4766 => "00000000",
	4767 => "00000000",
	4768 => "11111111",
	4769 => "11111111",
	4770 => "11111111",
	4771 => "11111111",
	4772 => "11111111",
	4773 => "11111111",
	4774 => "11111111",
	4775 => "11111111",
	4776 => "11111111",
	4777 => "11111111",
	4778 => "11111111",
	4779 => "00000000",
	4780 => "00000000",
	4781 => "00000000",
	4782 => "00000000",
	4783 => "00000000",
	4784 => "00000000",
	4785 => "00000000",
	4786 => "00000000",
	4787 => "00000000",
	4788 => "00000000",
	4789 => "00000000",
	4790 => "00000000",
	4791 => "00000000",
	4792 => "00000000",
	4793 => "00000000",
	4794 => "00000000",
	4795 => "00000000",
	4796 => "00000000",
	4797 => "00000000",
	4798 => "00000000",
	4799 => "00000000",
	4800 => "00000000",
	4801 => "00000000",
	4802 => "00000000",
	4803 => "00000000",
	4804 => "00000000",
	4805 => "00000000",
	4806 => "00000000",
	4807 => "00000000",
	4808 => "00000000",
	4809 => "00000000",
	4810 => "00000000",
	4811 => "00000000",
	4812 => "00000000",
	4813 => "00000000",
	4814 => "11111111",
	4815 => "11111111",
	4816 => "11111111",
	4817 => "11111111",
	4818 => "11111111",
	4819 => "11111111",
	4820 => "11111111",
	4821 => "11111111",
	4822 => "11111111",
	4823 => "11111111",
	4824 => "11111111",
	4825 => "00000000",
	4826 => "00000000",
	4827 => "00000000",
	4828 => "00000000",
	4829 => "00000000",
	4830 => "00000000",
	4831 => "00000000",
	4832 => "00000000",
	4833 => "00000000",
	4834 => "00000000",
	4835 => "00000000",
	4836 => "00000000",
	4837 => "00000000",
	4838 => "00000000",
	4839 => "00000000",
	4840 => "00000000",
	4841 => "00000000",
	4842 => "00000000",
	4843 => "00000000",
	4844 => "00000000",
	4845 => "00000000",
	4846 => "00000000",
	4847 => "00000000",
	4848 => "00000000",
	4849 => "00000000",
	4850 => "00000000",
	4851 => "00000000",
	4852 => "00000000",
	4853 => "00000000",
	4854 => "00000000",
	4855 => "00000000",
	4864 => "00000000",
	4865 => "00000000",
	4866 => "00000000",
	4867 => "00000000",
	4868 => "00000000",
	4869 => "00000000",
	4870 => "00000000",
	4871 => "00000000",
	4872 => "00000000",
	4873 => "00000000",
	4874 => "00000000",
	4875 => "00000000",
	4876 => "00000000",
	4877 => "00000000",
	4878 => "00000000",
	4879 => "00000000",
	4880 => "00000000",
	4881 => "00000000",
	4882 => "00000000",
	4883 => "00000000",
	4884 => "00000000",
	4885 => "00000000",
	4886 => "00000000",
	4887 => "00000000",
	4888 => "00000000",
	4889 => "00000000",
	4890 => "00000000",
	4891 => "00000000",
	4892 => "00000000",
	4893 => "00000000",
	4894 => "00000000",
	4895 => "00000000",
	4896 => "00000000",
	4897 => "11111111",
	4898 => "11111111",
	4899 => "11111111",
	4900 => "11111111",
	4901 => "11111111",
	4902 => "11111111",
	4903 => "11111111",
	4904 => "11111111",
	4905 => "11111111",
	4906 => "11111111",
	4907 => "11111111",
	4908 => "00000000",
	4909 => "00000000",
	4910 => "00000000",
	4911 => "00000000",
	4912 => "00000000",
	4913 => "00000000",
	4914 => "00000000",
	4915 => "00000000",
	4916 => "00000000",
	4917 => "00000000",
	4918 => "00000000",
	4919 => "00000000",
	4920 => "00000000",
	4921 => "00000000",
	4922 => "00000000",
	4923 => "00000000",
	4924 => "00000000",
	4925 => "00000000",
	4926 => "00000000",
	4927 => "00000000",
	4928 => "00000000",
	4929 => "00000000",
	4930 => "00000000",
	4931 => "00000000",
	4932 => "00000000",
	4933 => "00000000",
	4934 => "00000000",
	4935 => "00000000",
	4936 => "00000000",
	4937 => "00000000",
	4938 => "00000000",
	4939 => "00000000",
	4940 => "00000000",
	4941 => "11111111",
	4942 => "11111111",
	4943 => "11111111",
	4944 => "11111111",
	4945 => "11111111",
	4946 => "11111111",
	4947 => "11111111",
	4948 => "11111111",
	4949 => "11111111",
	4950 => "11111111",
	4951 => "11111111",
	4952 => "00000000",
	4953 => "00000000",
	4954 => "00000000",
	4955 => "00000000",
	4956 => "00000000",
	4957 => "00000000",
	4958 => "00000000",
	4959 => "00000000",
	4960 => "00000000",
	4961 => "00000000",
	4962 => "00000000",
	4963 => "00000000",
	4964 => "00000000",
	4965 => "00000000",
	4966 => "00000000",
	4967 => "00000000",
	4968 => "00000000",
	4969 => "00000000",
	4970 => "00000000",
	4971 => "00000000",
	4972 => "00000000",
	4973 => "00000000",
	4974 => "00000000",
	4975 => "00000000",
	4976 => "00000000",
	4977 => "00000000",
	4978 => "00000000",
	4979 => "00000000",
	4980 => "00000000",
	4981 => "00000000",
	4982 => "00000000",
	4983 => "00000000",
	4992 => "00000000",
	4993 => "00000000",
	4994 => "00000000",
	4995 => "00000000",
	4996 => "00000000",
	4997 => "00000000",
	4998 => "00000000",
	4999 => "00000000",
	5000 => "00000000",
	5001 => "00000000",
	5002 => "00000000",
	5003 => "00000000",
	5004 => "00000000",
	5005 => "00000000",
	5006 => "00000000",
	5007 => "00000000",
	5008 => "00000000",
	5009 => "00000000",
	5010 => "00000000",
	5011 => "00000000",
	5012 => "00000000",
	5013 => "00000000",
	5014 => "00000000",
	5015 => "00000000",
	5016 => "00000000",
	5017 => "00000000",
	5018 => "00000000",
	5019 => "00000000",
	5020 => "00000000",
	5021 => "00000000",
	5022 => "00000000",
	5023 => "00000000",
	5024 => "00000000",
	5025 => "00000000",
	5026 => "11111111",
	5027 => "11111111",
	5028 => "11111111",
	5029 => "11111111",
	5030 => "11111111",
	5031 => "11111111",
	5032 => "11111111",
	5033 => "11111111",
	5034 => "11111111",
	5035 => "11111111",
	5036 => "11111111",
	5037 => "00000000",
	5038 => "00000000",
	5039 => "00000000",
	5040 => "00000000",
	5041 => "00000000",
	5042 => "00000000",
	5043 => "00000000",
	5044 => "00000000",
	5045 => "00000000",
	5046 => "00000000",
	5047 => "00000000",
	5048 => "00000000",
	5049 => "00000000",
	5050 => "00000000",
	5051 => "00000000",
	5052 => "00000000",
	5053 => "00000000",
	5054 => "00000000",
	5055 => "00000000",
	5056 => "00000000",
	5057 => "00000000",
	5058 => "00000000",
	5059 => "00000000",
	5060 => "00000000",
	5061 => "00000000",
	5062 => "00000000",
	5063 => "00000000",
	5064 => "00000000",
	5065 => "00000000",
	5066 => "00000000",
	5067 => "00000000",
	5068 => "11111111",
	5069 => "11111111",
	5070 => "11111111",
	5071 => "11111111",
	5072 => "11111111",
	5073 => "11111111",
	5074 => "11111111",
	5075 => "11111111",
	5076 => "11111111",
	5077 => "11111111",
	5078 => "11111111",
	5079 => "00000000",
	5080 => "00000000",
	5081 => "00000000",
	5082 => "00000000",
	5083 => "00000000",
	5084 => "00000000",
	5085 => "00000000",
	5086 => "00000000",
	5087 => "00000000",
	5088 => "00000000",
	5089 => "00000000",
	5090 => "00000000",
	5091 => "00000000",
	5092 => "00000000",
	5093 => "00000000",
	5094 => "00000000",
	5095 => "00000000",
	5096 => "00000000",
	5097 => "00000000",
	5098 => "00000000",
	5099 => "00000000",
	5100 => "00000000",
	5101 => "00000000",
	5102 => "00000000",
	5103 => "00000000",
	5104 => "00000000",
	5105 => "00000000",
	5106 => "00000000",
	5107 => "00000000",
	5108 => "00000000",
	5109 => "00000000",
	5110 => "00000000",
	5111 => "00000000",
	5120 => "00000000",
	5121 => "00000000",
	5122 => "00000000",
	5123 => "00000000",
	5124 => "00000000",
	5125 => "00000000",
	5126 => "00000000",
	5127 => "00000000",
	5128 => "00000000",
	5129 => "00000000",
	5130 => "00000000",
	5131 => "00000000",
	5132 => "00000000",
	5133 => "00000000",
	5134 => "00000000",
	5135 => "00000000",
	5136 => "00000000",
	5137 => "00000000",
	5138 => "00000000",
	5139 => "00000000",
	5140 => "00000000",
	5141 => "00000000",
	5142 => "00000000",
	5143 => "00000000",
	5144 => "00000000",
	5145 => "00000000",
	5146 => "00000000",
	5147 => "00000000",
	5148 => "00000000",
	5149 => "00000000",
	5150 => "00000000",
	5151 => "00000000",
	5152 => "00000000",
	5153 => "00000000",
	5154 => "00000000",
	5155 => "11111111",
	5156 => "11111111",
	5157 => "11111111",
	5158 => "11111111",
	5159 => "11111111",
	5160 => "11111111",
	5161 => "11111111",
	5162 => "11111111",
	5163 => "11111111",
	5164 => "11111111",
	5165 => "11111111",
	5166 => "00000000",
	5167 => "00000000",
	5168 => "00000000",
	5169 => "00000000",
	5170 => "00000000",
	5171 => "00000000",
	5172 => "00000000",
	5173 => "00000000",
	5174 => "00000000",
	5175 => "00000000",
	5176 => "00000000",
	5177 => "00000000",
	5178 => "00000000",
	5179 => "00000000",
	5180 => "00000000",
	5181 => "00000000",
	5182 => "00000000",
	5183 => "00000000",
	5184 => "00000000",
	5185 => "00000000",
	5186 => "00000000",
	5187 => "00000000",
	5188 => "00000000",
	5189 => "00000000",
	5190 => "00000000",
	5191 => "00000000",
	5192 => "00000000",
	5193 => "00000000",
	5194 => "00000000",
	5195 => "11111111",
	5196 => "11111111",
	5197 => "11111111",
	5198 => "11111111",
	5199 => "11111111",
	5200 => "11111111",
	5201 => "11111111",
	5202 => "11111111",
	5203 => "11111111",
	5204 => "11111111",
	5205 => "11111111",
	5206 => "00000000",
	5207 => "00000000",
	5208 => "00000000",
	5209 => "00000000",
	5210 => "00000000",
	5211 => "00000000",
	5212 => "00000000",
	5213 => "00000000",
	5214 => "00000000",
	5215 => "00000000",
	5216 => "00000000",
	5217 => "00000000",
	5218 => "00000000",
	5219 => "00000000",
	5220 => "00000000",
	5221 => "00000000",
	5222 => "00000000",
	5223 => "00000000",
	5224 => "00000000",
	5225 => "00000000",
	5226 => "00000000",
	5227 => "00000000",
	5228 => "00000000",
	5229 => "00000000",
	5230 => "00000000",
	5231 => "00000000",
	5232 => "00000000",
	5233 => "00000000",
	5234 => "00000000",
	5235 => "00000000",
	5236 => "00000000",
	5237 => "00000000",
	5238 => "00000000",
	5239 => "00000000",
	5248 => "00000000",
	5249 => "00000000",
	5250 => "00000000",
	5251 => "00000000",
	5252 => "00000000",
	5253 => "00000000",
	5254 => "00000000",
	5255 => "00000000",
	5256 => "00000000",
	5257 => "00000000",
	5258 => "00000000",
	5259 => "00000000",
	5260 => "00000000",
	5261 => "00000000",
	5262 => "00000000",
	5263 => "00000000",
	5264 => "00000000",
	5265 => "00000000",
	5266 => "00000000",
	5267 => "00000000",
	5268 => "00000000",
	5269 => "00000000",
	5270 => "00000000",
	5271 => "00000000",
	5272 => "00000000",
	5273 => "00000000",
	5274 => "00000000",
	5275 => "00000000",
	5276 => "00000000",
	5277 => "00000000",
	5278 => "00000000",
	5279 => "00000000",
	5280 => "00000000",
	5281 => "00000000",
	5282 => "00000000",
	5283 => "00000000",
	5284 => "11111111",
	5285 => "11111111",
	5286 => "11111111",
	5287 => "11111111",
	5288 => "11111111",
	5289 => "11111111",
	5290 => "11111111",
	5291 => "11111111",
	5292 => "11111111",
	5293 => "11111111",
	5294 => "11111111",
	5295 => "00000000",
	5296 => "00000000",
	5297 => "00000000",
	5298 => "00000000",
	5299 => "00000000",
	5300 => "00000000",
	5301 => "00000000",
	5302 => "00000000",
	5303 => "00000000",
	5304 => "00000000",
	5305 => "00000000",
	5306 => "00000000",
	5307 => "00000000",
	5308 => "00000000",
	5309 => "00000000",
	5310 => "00000000",
	5311 => "00000000",
	5312 => "00000000",
	5313 => "00000000",
	5314 => "00000000",
	5315 => "00000000",
	5316 => "00000000",
	5317 => "00000000",
	5318 => "00000000",
	5319 => "00000000",
	5320 => "00000000",
	5321 => "00000000",
	5322 => "11111111",
	5323 => "11111111",
	5324 => "11111111",
	5325 => "11111111",
	5326 => "11111111",
	5327 => "11111111",
	5328 => "11111111",
	5329 => "11111111",
	5330 => "11111111",
	5331 => "11111111",
	5332 => "11111111",
	5333 => "00000000",
	5334 => "00000000",
	5335 => "00000000",
	5336 => "00000000",
	5337 => "00000000",
	5338 => "00000000",
	5339 => "00000000",
	5340 => "00000000",
	5341 => "00000000",
	5342 => "00000000",
	5343 => "00000000",
	5344 => "00000000",
	5345 => "00000000",
	5346 => "00000000",
	5347 => "00000000",
	5348 => "00000000",
	5349 => "00000000",
	5350 => "00000000",
	5351 => "00000000",
	5352 => "00000000",
	5353 => "00000000",
	5354 => "00000000",
	5355 => "00000000",
	5356 => "00000000",
	5357 => "00000000",
	5358 => "00000000",
	5359 => "00000000",
	5360 => "00000000",
	5361 => "00000000",
	5362 => "00000000",
	5363 => "00000000",
	5364 => "00000000",
	5365 => "00000000",
	5366 => "00000000",
	5367 => "00000000",
	5376 => "00000000",
	5377 => "00000000",
	5378 => "00000000",
	5379 => "00000000",
	5380 => "00000000",
	5381 => "00000000",
	5382 => "00000000",
	5383 => "00000000",
	5384 => "00000000",
	5385 => "00000000",
	5386 => "00000000",
	5387 => "00000000",
	5388 => "00000000",
	5389 => "00000000",
	5390 => "00000000",
	5391 => "00000000",
	5392 => "00000000",
	5393 => "00000000",
	5394 => "00000000",
	5395 => "00000000",
	5396 => "00000000",
	5397 => "00000000",
	5398 => "00000000",
	5399 => "00000000",
	5400 => "00000000",
	5401 => "00000000",
	5402 => "00000000",
	5403 => "00000000",
	5404 => "00000000",
	5405 => "00000000",
	5406 => "00000000",
	5407 => "00000000",
	5408 => "00000000",
	5409 => "00000000",
	5410 => "00000000",
	5411 => "00000000",
	5412 => "00000000",
	5413 => "11111111",
	5414 => "11111111",
	5415 => "11111111",
	5416 => "11111111",
	5417 => "11111111",
	5418 => "11111111",
	5419 => "11111111",
	5420 => "11111111",
	5421 => "11111111",
	5422 => "11111111",
	5423 => "11111111",
	5424 => "00000000",
	5425 => "00000000",
	5426 => "00000000",
	5427 => "00000000",
	5428 => "00000000",
	5429 => "00000000",
	5430 => "00000000",
	5431 => "00000000",
	5432 => "00000000",
	5433 => "00000000",
	5434 => "00000000",
	5435 => "00000000",
	5436 => "00000000",
	5437 => "00000000",
	5438 => "00000000",
	5439 => "00000000",
	5440 => "00000000",
	5441 => "00000000",
	5442 => "00000000",
	5443 => "00000000",
	5444 => "00000000",
	5445 => "00000000",
	5446 => "00000000",
	5447 => "00000000",
	5448 => "00000000",
	5449 => "11111111",
	5450 => "11111111",
	5451 => "11111111",
	5452 => "11111111",
	5453 => "11111111",
	5454 => "11111111",
	5455 => "11111111",
	5456 => "11111111",
	5457 => "11111111",
	5458 => "11111111",
	5459 => "11111111",
	5460 => "00000000",
	5461 => "00000000",
	5462 => "00000000",
	5463 => "00000000",
	5464 => "00000000",
	5465 => "00000000",
	5466 => "00000000",
	5467 => "00000000",
	5468 => "00000000",
	5469 => "00000000",
	5470 => "00000000",
	5471 => "00000000",
	5472 => "00000000",
	5473 => "00000000",
	5474 => "00000000",
	5475 => "00000000",
	5476 => "00000000",
	5477 => "00000000",
	5478 => "00000000",
	5479 => "00000000",
	5480 => "00000000",
	5481 => "00000000",
	5482 => "00000000",
	5483 => "00000000",
	5484 => "00000000",
	5485 => "00000000",
	5486 => "00000000",
	5487 => "00000000",
	5488 => "00000000",
	5489 => "00000000",
	5490 => "00000000",
	5491 => "00000000",
	5492 => "00000000",
	5493 => "00000000",
	5494 => "00000000",
	5495 => "00000000",
	5504 => "00000000",
	5505 => "00000000",
	5506 => "00000000",
	5507 => "00000000",
	5508 => "00000000",
	5509 => "00000000",
	5510 => "00000000",
	5511 => "00000000",
	5512 => "00000000",
	5513 => "00000000",
	5514 => "00000000",
	5515 => "00000000",
	5516 => "00000000",
	5517 => "00000000",
	5518 => "00000000",
	5519 => "00000000",
	5520 => "00000000",
	5521 => "00000000",
	5522 => "00000000",
	5523 => "00000000",
	5524 => "00000000",
	5525 => "00000000",
	5526 => "00000000",
	5527 => "00000000",
	5528 => "00000000",
	5529 => "00000000",
	5530 => "00000000",
	5531 => "00000000",
	5532 => "00000000",
	5533 => "00000000",
	5534 => "00000000",
	5535 => "00000000",
	5536 => "00000000",
	5537 => "00000000",
	5538 => "00000000",
	5539 => "00000000",
	5540 => "00000000",
	5541 => "00000000",
	5542 => "11111111",
	5543 => "11111111",
	5544 => "11111111",
	5545 => "11111111",
	5546 => "11111111",
	5547 => "11111111",
	5548 => "11111111",
	5549 => "11111111",
	5550 => "11111111",
	5551 => "11111111",
	5552 => "11111111",
	5553 => "00000000",
	5554 => "00000000",
	5555 => "00000000",
	5556 => "00000000",
	5557 => "00000000",
	5558 => "00000000",
	5559 => "00000000",
	5560 => "00000000",
	5561 => "00000000",
	5562 => "00000000",
	5563 => "00000000",
	5564 => "00000000",
	5565 => "00000000",
	5566 => "00000000",
	5567 => "00000000",
	5568 => "00000000",
	5569 => "00000000",
	5570 => "00000000",
	5571 => "00000000",
	5572 => "00000000",
	5573 => "00000000",
	5574 => "00000000",
	5575 => "00000000",
	5576 => "11111111",
	5577 => "11111111",
	5578 => "11111111",
	5579 => "11111111",
	5580 => "11111111",
	5581 => "11111111",
	5582 => "11111111",
	5583 => "11111111",
	5584 => "11111111",
	5585 => "11111111",
	5586 => "11111111",
	5587 => "00000000",
	5588 => "00000000",
	5589 => "00000000",
	5590 => "00000000",
	5591 => "00000000",
	5592 => "00000000",
	5593 => "00000000",
	5594 => "00000000",
	5595 => "00000000",
	5596 => "00000000",
	5597 => "00000000",
	5598 => "00000000",
	5599 => "00000000",
	5600 => "00000000",
	5601 => "00000000",
	5602 => "00000000",
	5603 => "00000000",
	5604 => "00000000",
	5605 => "00000000",
	5606 => "00000000",
	5607 => "00000000",
	5608 => "00000000",
	5609 => "00000000",
	5610 => "00000000",
	5611 => "00000000",
	5612 => "00000000",
	5613 => "00000000",
	5614 => "00000000",
	5615 => "00000000",
	5616 => "00000000",
	5617 => "00000000",
	5618 => "00000000",
	5619 => "00000000",
	5620 => "00000000",
	5621 => "00000000",
	5622 => "00000000",
	5623 => "00000000",
	5632 => "00000000",
	5633 => "00000000",
	5634 => "00000000",
	5635 => "00000000",
	5636 => "00000000",
	5637 => "00000000",
	5638 => "00000000",
	5639 => "00000000",
	5640 => "00000000",
	5641 => "00000000",
	5642 => "00000000",
	5643 => "00000000",
	5644 => "00000000",
	5645 => "00000000",
	5646 => "00000000",
	5647 => "00000000",
	5648 => "00000000",
	5649 => "00000000",
	5650 => "00000000",
	5651 => "00000000",
	5652 => "00000000",
	5653 => "00000000",
	5654 => "00000000",
	5655 => "00000000",
	5656 => "00000000",
	5657 => "00000000",
	5658 => "00000000",
	5659 => "00000000",
	5660 => "00000000",
	5661 => "00000000",
	5662 => "00000000",
	5663 => "00000000",
	5664 => "00000000",
	5665 => "00000000",
	5666 => "00000000",
	5667 => "00000000",
	5668 => "00000000",
	5669 => "00000000",
	5670 => "00000000",
	5671 => "11111111",
	5672 => "11111111",
	5673 => "11111111",
	5674 => "11111111",
	5675 => "11111111",
	5676 => "11111111",
	5677 => "11111111",
	5678 => "11111111",
	5679 => "11111111",
	5680 => "11111111",
	5681 => "11111111",
	5682 => "00000000",
	5683 => "00000000",
	5684 => "00000000",
	5685 => "00000000",
	5686 => "00000000",
	5687 => "00000000",
	5688 => "00000000",
	5689 => "00000000",
	5690 => "00000000",
	5691 => "00000000",
	5692 => "00000000",
	5693 => "00000000",
	5694 => "00000000",
	5695 => "00000000",
	5696 => "00000000",
	5697 => "00000000",
	5698 => "00000000",
	5699 => "00000000",
	5700 => "00000000",
	5701 => "00000000",
	5702 => "00000000",
	5703 => "11111111",
	5704 => "11111111",
	5705 => "11111111",
	5706 => "11111111",
	5707 => "11111111",
	5708 => "11111111",
	5709 => "11111111",
	5710 => "11111111",
	5711 => "11111111",
	5712 => "11111111",
	5713 => "11111111",
	5714 => "00000000",
	5715 => "00000000",
	5716 => "00000000",
	5717 => "00000000",
	5718 => "00000000",
	5719 => "00000000",
	5720 => "00000000",
	5721 => "00000000",
	5722 => "00000000",
	5723 => "00000000",
	5724 => "00000000",
	5725 => "00000000",
	5726 => "00000000",
	5727 => "00000000",
	5728 => "00000000",
	5729 => "00000000",
	5730 => "00000000",
	5731 => "00000000",
	5732 => "00000000",
	5733 => "00000000",
	5734 => "00000000",
	5735 => "00000000",
	5736 => "00000000",
	5737 => "00000000",
	5738 => "00000000",
	5739 => "00000000",
	5740 => "00000000",
	5741 => "00000000",
	5742 => "00000000",
	5743 => "00000000",
	5744 => "00000000",
	5745 => "00000000",
	5746 => "00000000",
	5747 => "00000000",
	5748 => "00000000",
	5749 => "00000000",
	5750 => "00000000",
	5751 => "00000000",
	5760 => "00000000",
	5761 => "00000000",
	5762 => "00000000",
	5763 => "00000000",
	5764 => "00000000",
	5765 => "00000000",
	5766 => "00000000",
	5767 => "00000000",
	5768 => "00000000",
	5769 => "00000000",
	5770 => "00000000",
	5771 => "00000000",
	5772 => "00000000",
	5773 => "00000000",
	5774 => "00000000",
	5775 => "00000000",
	5776 => "00000000",
	5777 => "00000000",
	5778 => "00000000",
	5779 => "00000000",
	5780 => "00000000",
	5781 => "00000000",
	5782 => "00000000",
	5783 => "00000000",
	5784 => "00000000",
	5785 => "00000000",
	5786 => "00000000",
	5787 => "00000000",
	5788 => "00000000",
	5789 => "00000000",
	5790 => "00000000",
	5791 => "00000000",
	5792 => "00000000",
	5793 => "00000000",
	5794 => "00000000",
	5795 => "00000000",
	5796 => "00000000",
	5797 => "00000000",
	5798 => "00000000",
	5799 => "00000000",
	5800 => "11111111",
	5801 => "11111111",
	5802 => "11111111",
	5803 => "11111111",
	5804 => "11111111",
	5805 => "11111111",
	5806 => "11111111",
	5807 => "11111111",
	5808 => "11111111",
	5809 => "11111111",
	5810 => "11111111",
	5811 => "00000000",
	5812 => "00000000",
	5813 => "00000000",
	5814 => "00000000",
	5815 => "00000000",
	5816 => "00000000",
	5817 => "00000000",
	5818 => "00000000",
	5819 => "00000000",
	5820 => "00000000",
	5821 => "00000000",
	5822 => "00000000",
	5823 => "00000000",
	5824 => "00000000",
	5825 => "00000000",
	5826 => "00000000",
	5827 => "00000000",
	5828 => "00000000",
	5829 => "00000000",
	5830 => "11111111",
	5831 => "11111111",
	5832 => "11111111",
	5833 => "11111111",
	5834 => "11111111",
	5835 => "11111111",
	5836 => "11111111",
	5837 => "11111111",
	5838 => "11111111",
	5839 => "11111111",
	5840 => "11111111",
	5841 => "00000000",
	5842 => "00000000",
	5843 => "00000000",
	5844 => "00000000",
	5845 => "00000000",
	5846 => "00000000",
	5847 => "00000000",
	5848 => "00000000",
	5849 => "00000000",
	5850 => "00000000",
	5851 => "00000000",
	5852 => "00000000",
	5853 => "00000000",
	5854 => "00000000",
	5855 => "00000000",
	5856 => "00000000",
	5857 => "00000000",
	5858 => "00000000",
	5859 => "00000000",
	5860 => "00000000",
	5861 => "00000000",
	5862 => "00000000",
	5863 => "00000000",
	5864 => "00000000",
	5865 => "00000000",
	5866 => "00000000",
	5867 => "00000000",
	5868 => "00000000",
	5869 => "00000000",
	5870 => "00000000",
	5871 => "00000000",
	5872 => "00000000",
	5873 => "00000000",
	5874 => "00000000",
	5875 => "00000000",
	5876 => "00000000",
	5877 => "00000000",
	5878 => "00000000",
	5879 => "00000000",
	5888 => "00000000",
	5889 => "00000000",
	5890 => "00000000",
	5891 => "00000000",
	5892 => "00000000",
	5893 => "00000000",
	5894 => "00000000",
	5895 => "00000000",
	5896 => "00000000",
	5897 => "00000000",
	5898 => "00000000",
	5899 => "00000000",
	5900 => "00000000",
	5901 => "00000000",
	5902 => "00000000",
	5903 => "00000000",
	5904 => "00000000",
	5905 => "00000000",
	5906 => "00000000",
	5907 => "00000000",
	5908 => "00000000",
	5909 => "00000000",
	5910 => "00000000",
	5911 => "00000000",
	5912 => "00000000",
	5913 => "00000000",
	5914 => "00000000",
	5915 => "00000000",
	5916 => "00000000",
	5917 => "00000000",
	5918 => "00000000",
	5919 => "00000000",
	5920 => "00000000",
	5921 => "00000000",
	5922 => "00000000",
	5923 => "00000000",
	5924 => "00000000",
	5925 => "00000000",
	5926 => "00000000",
	5927 => "00000000",
	5928 => "00000000",
	5929 => "11111111",
	5930 => "11111111",
	5931 => "11111111",
	5932 => "11111111",
	5933 => "11111111",
	5934 => "11111111",
	5935 => "11111111",
	5936 => "11111111",
	5937 => "11111111",
	5938 => "11111111",
	5939 => "11111111",
	5940 => "00000000",
	5941 => "00000000",
	5942 => "00000000",
	5943 => "00000000",
	5944 => "00000000",
	5945 => "00000000",
	5946 => "00000000",
	5947 => "00000000",
	5948 => "00000000",
	5949 => "00000000",
	5950 => "00000000",
	5951 => "00000000",
	5952 => "00000000",
	5953 => "00000000",
	5954 => "00000000",
	5955 => "00000000",
	5956 => "00000000",
	5957 => "11111111",
	5958 => "11111111",
	5959 => "11111111",
	5960 => "11111111",
	5961 => "11111111",
	5962 => "11111111",
	5963 => "11111111",
	5964 => "11111111",
	5965 => "11111111",
	5966 => "11111111",
	5967 => "11111111",
	5968 => "00000000",
	5969 => "00000000",
	5970 => "00000000",
	5971 => "00000000",
	5972 => "00000000",
	5973 => "00000000",
	5974 => "00000000",
	5975 => "00000000",
	5976 => "00000000",
	5977 => "00000000",
	5978 => "00000000",
	5979 => "00000000",
	5980 => "00000000",
	5981 => "00000000",
	5982 => "00000000",
	5983 => "00000000",
	5984 => "00000000",
	5985 => "00000000",
	5986 => "00000000",
	5987 => "00000000",
	5988 => "00000000",
	5989 => "00000000",
	5990 => "00000000",
	5991 => "00000000",
	5992 => "00000000",
	5993 => "00000000",
	5994 => "00000000",
	5995 => "00000000",
	5996 => "00000000",
	5997 => "00000000",
	5998 => "00000000",
	5999 => "00000000",
	6000 => "00000000",
	6001 => "00000000",
	6002 => "00000000",
	6003 => "00000000",
	6004 => "00000000",
	6005 => "00000000",
	6006 => "00000000",
	6007 => "00000000",
	6016 => "00000000",
	6017 => "00000000",
	6018 => "00000000",
	6019 => "00000000",
	6020 => "00000000",
	6021 => "00000000",
	6022 => "00000000",
	6023 => "00000000",
	6024 => "00000000",
	6025 => "00000000",
	6026 => "00000000",
	6027 => "00000000",
	6028 => "00000000",
	6029 => "00000000",
	6030 => "00000000",
	6031 => "00000000",
	6032 => "00000000",
	6033 => "00000000",
	6034 => "00000000",
	6035 => "00000000",
	6036 => "00000000",
	6037 => "00000000",
	6038 => "00000000",
	6039 => "00000000",
	6040 => "00000000",
	6041 => "00000000",
	6042 => "00000000",
	6043 => "00000000",
	6044 => "00000000",
	6045 => "00000000",
	6046 => "00000000",
	6047 => "00000000",
	6048 => "00000000",
	6049 => "00000000",
	6050 => "00000000",
	6051 => "00000000",
	6052 => "00000000",
	6053 => "00000000",
	6054 => "00000000",
	6055 => "00000000",
	6056 => "00000000",
	6057 => "00000000",
	6058 => "11111111",
	6059 => "11111111",
	6060 => "11111111",
	6061 => "11111111",
	6062 => "11111111",
	6063 => "11111111",
	6064 => "11111111",
	6065 => "11111111",
	6066 => "11111111",
	6067 => "11111111",
	6068 => "11111111",
	6069 => "00000000",
	6070 => "00000000",
	6071 => "00000000",
	6072 => "00000000",
	6073 => "00000000",
	6074 => "00000000",
	6075 => "00000000",
	6076 => "00000000",
	6077 => "00000000",
	6078 => "00000000",
	6079 => "00000000",
	6080 => "00000000",
	6081 => "00000000",
	6082 => "00000000",
	6083 => "00000000",
	6084 => "11111111",
	6085 => "11111111",
	6086 => "11111111",
	6087 => "11111111",
	6088 => "11111111",
	6089 => "11111111",
	6090 => "11111111",
	6091 => "11111111",
	6092 => "11111111",
	6093 => "11111111",
	6094 => "11111111",
	6095 => "00000000",
	6096 => "00000000",
	6097 => "00000000",
	6098 => "00000000",
	6099 => "00000000",
	6100 => "00000000",
	6101 => "00000000",
	6102 => "00000000",
	6103 => "00000000",
	6104 => "00000000",
	6105 => "00000000",
	6106 => "00000000",
	6107 => "00000000",
	6108 => "00000000",
	6109 => "00000000",
	6110 => "00000000",
	6111 => "00000000",
	6112 => "00000000",
	6113 => "00000000",
	6114 => "00000000",
	6115 => "00000000",
	6116 => "00000000",
	6117 => "00000000",
	6118 => "00000000",
	6119 => "00000000",
	6120 => "00000000",
	6121 => "00000000",
	6122 => "00000000",
	6123 => "00000000",
	6124 => "00000000",
	6125 => "00000000",
	6126 => "00000000",
	6127 => "00000000",
	6128 => "00000000",
	6129 => "00000000",
	6130 => "00000000",
	6131 => "00000000",
	6132 => "00000000",
	6133 => "00000000",
	6134 => "00000000",
	6135 => "00000000",
	6144 => "00000000",
	6145 => "00000000",
	6146 => "00000000",
	6147 => "00000000",
	6148 => "00000000",
	6149 => "00000000",
	6150 => "00000000",
	6151 => "00000000",
	6152 => "00000000",
	6153 => "00000000",
	6154 => "00000000",
	6155 => "00000000",
	6156 => "00000000",
	6157 => "00000000",
	6158 => "00000000",
	6159 => "00000000",
	6160 => "00000000",
	6161 => "00000000",
	6162 => "00000000",
	6163 => "00000000",
	6164 => "00000000",
	6165 => "00000000",
	6166 => "00000000",
	6167 => "00000000",
	6168 => "00000000",
	6169 => "00000000",
	6170 => "00000000",
	6171 => "00000000",
	6172 => "00000000",
	6173 => "00000000",
	6174 => "00000000",
	6175 => "00000000",
	6176 => "00000000",
	6177 => "00000000",
	6178 => "00000000",
	6179 => "00000000",
	6180 => "00000000",
	6181 => "00000000",
	6182 => "00000000",
	6183 => "00000000",
	6184 => "00000000",
	6185 => "00000000",
	6186 => "00000000",
	6187 => "11111111",
	6188 => "11111111",
	6189 => "11111111",
	6190 => "11111111",
	6191 => "11111111",
	6192 => "11111111",
	6193 => "11111111",
	6194 => "11111111",
	6195 => "11111111",
	6196 => "11111111",
	6197 => "11111111",
	6198 => "00000000",
	6199 => "00000000",
	6200 => "00000000",
	6201 => "00000000",
	6202 => "00000000",
	6203 => "00000000",
	6204 => "00000000",
	6205 => "00000000",
	6206 => "00000000",
	6207 => "00000000",
	6208 => "00000000",
	6209 => "00000000",
	6210 => "00000000",
	6211 => "11111111",
	6212 => "11111111",
	6213 => "11111111",
	6214 => "11111111",
	6215 => "11111111",
	6216 => "11111111",
	6217 => "11111111",
	6218 => "11111111",
	6219 => "11111111",
	6220 => "11111111",
	6221 => "11111111",
	6222 => "00000000",
	6223 => "00000000",
	6224 => "00000000",
	6225 => "00000000",
	6226 => "00000000",
	6227 => "00000000",
	6228 => "00000000",
	6229 => "00000000",
	6230 => "00000000",
	6231 => "00000000",
	6232 => "00000000",
	6233 => "00000000",
	6234 => "00000000",
	6235 => "00000000",
	6236 => "00000000",
	6237 => "00000000",
	6238 => "00000000",
	6239 => "00000000",
	6240 => "00000000",
	6241 => "00000000",
	6242 => "00000000",
	6243 => "00000000",
	6244 => "00000000",
	6245 => "00000000",
	6246 => "00000000",
	6247 => "00000000",
	6248 => "00000000",
	6249 => "00000000",
	6250 => "00000000",
	6251 => "00000000",
	6252 => "00000000",
	6253 => "00000000",
	6254 => "00000000",
	6255 => "00000000",
	6256 => "00000000",
	6257 => "00000000",
	6258 => "00000000",
	6259 => "00000000",
	6260 => "00000000",
	6261 => "00000000",
	6262 => "00000000",
	6263 => "00000000",
	6272 => "00000000",
	6273 => "00000000",
	6274 => "00000000",
	6275 => "00000000",
	6276 => "00000000",
	6277 => "00000000",
	6278 => "00000000",
	6279 => "00000000",
	6280 => "00000000",
	6281 => "00000000",
	6282 => "00000000",
	6283 => "00000000",
	6284 => "00000000",
	6285 => "00000000",
	6286 => "00000000",
	6287 => "00000000",
	6288 => "00000000",
	6289 => "00000000",
	6290 => "00000000",
	6291 => "00000000",
	6292 => "00000000",
	6293 => "00000000",
	6294 => "00000000",
	6295 => "00000000",
	6296 => "00000000",
	6297 => "00000000",
	6298 => "00000000",
	6299 => "00000000",
	6300 => "00000000",
	6301 => "00000000",
	6302 => "00000000",
	6303 => "00000000",
	6304 => "00000000",
	6305 => "00000000",
	6306 => "00000000",
	6307 => "00000000",
	6308 => "00000000",
	6309 => "00000000",
	6310 => "00000000",
	6311 => "00000000",
	6312 => "00000000",
	6313 => "00000000",
	6314 => "00000000",
	6315 => "00000000",
	6316 => "11111111",
	6317 => "11111111",
	6318 => "11111111",
	6319 => "11111111",
	6320 => "11111111",
	6321 => "11111111",
	6322 => "11111111",
	6323 => "11111111",
	6324 => "11111111",
	6325 => "11111111",
	6326 => "11111111",
	6327 => "00000000",
	6328 => "00000000",
	6329 => "00000000",
	6330 => "00000000",
	6331 => "00000000",
	6332 => "00000000",
	6333 => "00000000",
	6334 => "00000000",
	6335 => "00000000",
	6336 => "00000000",
	6337 => "00000000",
	6338 => "11111111",
	6339 => "11111111",
	6340 => "11111111",
	6341 => "11111111",
	6342 => "11111111",
	6343 => "11111111",
	6344 => "11111111",
	6345 => "11111111",
	6346 => "11111111",
	6347 => "11111111",
	6348 => "11111111",
	6349 => "00000000",
	6350 => "00000000",
	6351 => "00000000",
	6352 => "00000000",
	6353 => "00000000",
	6354 => "00000000",
	6355 => "00000000",
	6356 => "00000000",
	6357 => "00000000",
	6358 => "00000000",
	6359 => "00000000",
	6360 => "00000000",
	6361 => "00000000",
	6362 => "00000000",
	6363 => "00000000",
	6364 => "00000000",
	6365 => "00000000",
	6366 => "00000000",
	6367 => "00000000",
	6368 => "00000000",
	6369 => "00000000",
	6370 => "00000000",
	6371 => "00000000",
	6372 => "00000000",
	6373 => "00000000",
	6374 => "00000000",
	6375 => "00000000",
	6376 => "00000000",
	6377 => "00000000",
	6378 => "00000000",
	6379 => "00000000",
	6380 => "00000000",
	6381 => "00000000",
	6382 => "00000000",
	6383 => "00000000",
	6384 => "00000000",
	6385 => "00000000",
	6386 => "00000000",
	6387 => "00000000",
	6388 => "00000000",
	6389 => "00000000",
	6390 => "00000000",
	6391 => "00000000",
	6400 => "00000000",
	6401 => "00000000",
	6402 => "00000000",
	6403 => "00000000",
	6404 => "00000000",
	6405 => "00000000",
	6406 => "00000000",
	6407 => "00000000",
	6408 => "00000000",
	6409 => "00000000",
	6410 => "00000000",
	6411 => "00000000",
	6412 => "00000000",
	6413 => "00000000",
	6414 => "00000000",
	6415 => "00000000",
	6416 => "00000000",
	6417 => "00000000",
	6418 => "00000000",
	6419 => "00000000",
	6420 => "00000000",
	6421 => "00000000",
	6422 => "00000000",
	6423 => "00000000",
	6424 => "00000000",
	6425 => "00000000",
	6426 => "00000000",
	6427 => "00000000",
	6428 => "00000000",
	6429 => "00000000",
	6430 => "00000000",
	6431 => "00000000",
	6432 => "00000000",
	6433 => "00000000",
	6434 => "00000000",
	6435 => "00000000",
	6436 => "00000000",
	6437 => "00000000",
	6438 => "00000000",
	6439 => "00000000",
	6440 => "00000000",
	6441 => "00000000",
	6442 => "00000000",
	6443 => "00000000",
	6444 => "00000000",
	6445 => "11111111",
	6446 => "11111111",
	6447 => "11111111",
	6448 => "11111111",
	6449 => "11111111",
	6450 => "11111111",
	6451 => "11111111",
	6452 => "11111111",
	6453 => "11111111",
	6454 => "11111111",
	6455 => "11111111",
	6456 => "00000000",
	6457 => "00000000",
	6458 => "00000000",
	6459 => "00000000",
	6460 => "00000000",
	6461 => "00000000",
	6462 => "00000000",
	6463 => "00000000",
	6464 => "00000000",
	6465 => "11111111",
	6466 => "11111111",
	6467 => "11111111",
	6468 => "11111111",
	6469 => "11111111",
	6470 => "11111111",
	6471 => "11111111",
	6472 => "11111111",
	6473 => "11111111",
	6474 => "11111111",
	6475 => "11111111",
	6476 => "00000000",
	6477 => "00000000",
	6478 => "00000000",
	6479 => "00000000",
	6480 => "00000000",
	6481 => "00000000",
	6482 => "00000000",
	6483 => "00000000",
	6484 => "00000000",
	6485 => "00000000",
	6486 => "00000000",
	6487 => "00000000",
	6488 => "00000000",
	6489 => "00000000",
	6490 => "00000000",
	6491 => "00000000",
	6492 => "00000000",
	6493 => "00000000",
	6494 => "00000000",
	6495 => "00000000",
	6496 => "00000000",
	6497 => "00000000",
	6498 => "00000000",
	6499 => "00000000",
	6500 => "00000000",
	6501 => "00000000",
	6502 => "00000000",
	6503 => "00000000",
	6504 => "00000000",
	6505 => "00000000",
	6506 => "00000000",
	6507 => "00000000",
	6508 => "00000000",
	6509 => "00000000",
	6510 => "00000000",
	6511 => "00000000",
	6512 => "00000000",
	6513 => "00000000",
	6514 => "00000000",
	6515 => "00000000",
	6516 => "00000000",
	6517 => "00000000",
	6518 => "00000000",
	6519 => "00000000",
	6528 => "00000000",
	6529 => "00000000",
	6530 => "00000000",
	6531 => "00000000",
	6532 => "00000000",
	6533 => "00000000",
	6534 => "00000000",
	6535 => "00000000",
	6536 => "00000000",
	6537 => "00000000",
	6538 => "00000000",
	6539 => "00000000",
	6540 => "00000000",
	6541 => "00000000",
	6542 => "00000000",
	6543 => "00000000",
	6544 => "00000000",
	6545 => "00000000",
	6546 => "00000000",
	6547 => "00000000",
	6548 => "00000000",
	6549 => "00000000",
	6550 => "00000000",
	6551 => "00000000",
	6552 => "00000000",
	6553 => "00000000",
	6554 => "00000000",
	6555 => "00000000",
	6556 => "00000000",
	6557 => "00000000",
	6558 => "00000000",
	6559 => "00000000",
	6560 => "00000000",
	6561 => "00000000",
	6562 => "00000000",
	6563 => "00000000",
	6564 => "00000000",
	6565 => "00000000",
	6566 => "00000000",
	6567 => "00000000",
	6568 => "00000000",
	6569 => "00000000",
	6570 => "00000000",
	6571 => "00000000",
	6572 => "00000000",
	6573 => "00000000",
	6574 => "11111111",
	6575 => "11111111",
	6576 => "11111111",
	6577 => "11111111",
	6578 => "11111111",
	6579 => "11111111",
	6580 => "11111111",
	6581 => "11111111",
	6582 => "11111111",
	6583 => "11111111",
	6584 => "11111111",
	6585 => "00000000",
	6586 => "00000000",
	6587 => "00000000",
	6588 => "00000000",
	6589 => "00000000",
	6590 => "00000000",
	6591 => "00000000",
	6592 => "11111111",
	6593 => "11111111",
	6594 => "11111111",
	6595 => "11111111",
	6596 => "11111111",
	6597 => "11111111",
	6598 => "11111111",
	6599 => "11111111",
	6600 => "11111111",
	6601 => "11111111",
	6602 => "11111111",
	6603 => "00000000",
	6604 => "00000000",
	6605 => "00000000",
	6606 => "00000000",
	6607 => "00000000",
	6608 => "00000000",
	6609 => "00000000",
	6610 => "00000000",
	6611 => "00000000",
	6612 => "00000000",
	6613 => "00000000",
	6614 => "00000000",
	6615 => "00000000",
	6616 => "00000000",
	6617 => "00000000",
	6618 => "00000000",
	6619 => "00000000",
	6620 => "00000000",
	6621 => "00000000",
	6622 => "00000000",
	6623 => "00000000",
	6624 => "00000000",
	6625 => "00000000",
	6626 => "00000000",
	6627 => "00000000",
	6628 => "00000000",
	6629 => "00000000",
	6630 => "00000000",
	6631 => "00000000",
	6632 => "00000000",
	6633 => "00000000",
	6634 => "00000000",
	6635 => "00000000",
	6636 => "00000000",
	6637 => "00000000",
	6638 => "00000000",
	6639 => "00000000",
	6640 => "00000000",
	6641 => "00000000",
	6642 => "00000000",
	6643 => "00000000",
	6644 => "00000000",
	6645 => "00000000",
	6646 => "00000000",
	6647 => "00000000",
	6656 => "00000000",
	6657 => "00000000",
	6658 => "00000000",
	6659 => "00000000",
	6660 => "00000000",
	6661 => "00000000",
	6662 => "00000000",
	6663 => "00000000",
	6664 => "00000000",
	6665 => "00000000",
	6666 => "00000000",
	6667 => "00000000",
	6668 => "00000000",
	6669 => "00000000",
	6670 => "00000000",
	6671 => "00000000",
	6672 => "00000000",
	6673 => "00000000",
	6674 => "00000000",
	6675 => "00000000",
	6676 => "00000000",
	6677 => "00000000",
	6678 => "00000000",
	6679 => "00000000",
	6680 => "00000000",
	6681 => "00000000",
	6682 => "00000000",
	6683 => "00000000",
	6684 => "00000000",
	6685 => "00000000",
	6686 => "00000000",
	6687 => "00000000",
	6688 => "00000000",
	6689 => "00000000",
	6690 => "00000000",
	6691 => "00000000",
	6692 => "00000000",
	6693 => "00000000",
	6694 => "00000000",
	6695 => "00000000",
	6696 => "00000000",
	6697 => "00000000",
	6698 => "00000000",
	6699 => "00000000",
	6700 => "00000000",
	6701 => "00000000",
	6702 => "00000000",
	6703 => "11111111",
	6704 => "11111111",
	6705 => "11111111",
	6706 => "11111111",
	6707 => "11111111",
	6708 => "11111111",
	6709 => "11111111",
	6710 => "11111111",
	6711 => "11111111",
	6712 => "11111111",
	6713 => "11111111",
	6714 => "00000000",
	6715 => "00000000",
	6716 => "00000000",
	6717 => "00000000",
	6718 => "00000000",
	6719 => "11111111",
	6720 => "11111111",
	6721 => "11111111",
	6722 => "11111111",
	6723 => "11111111",
	6724 => "11111111",
	6725 => "11111111",
	6726 => "11111111",
	6727 => "11111111",
	6728 => "11111111",
	6729 => "11111111",
	6730 => "00000000",
	6731 => "00000000",
	6732 => "00000000",
	6733 => "00000000",
	6734 => "00000000",
	6735 => "00000000",
	6736 => "00000000",
	6737 => "00000000",
	6738 => "00000000",
	6739 => "00000000",
	6740 => "00000000",
	6741 => "00000000",
	6742 => "00000000",
	6743 => "00000000",
	6744 => "00000000",
	6745 => "00000000",
	6746 => "00000000",
	6747 => "00000000",
	6748 => "00000000",
	6749 => "00000000",
	6750 => "00000000",
	6751 => "00000000",
	6752 => "00000000",
	6753 => "00000000",
	6754 => "00000000",
	6755 => "00000000",
	6756 => "00000000",
	6757 => "00000000",
	6758 => "00000000",
	6759 => "00000000",
	6760 => "00000000",
	6761 => "00000000",
	6762 => "00000000",
	6763 => "00000000",
	6764 => "00000000",
	6765 => "00000000",
	6766 => "00000000",
	6767 => "00000000",
	6768 => "00000000",
	6769 => "00000000",
	6770 => "00000000",
	6771 => "00000000",
	6772 => "00000000",
	6773 => "00000000",
	6774 => "00000000",
	6775 => "00000000",
	6784 => "00000000",
	6785 => "00000000",
	6786 => "00000000",
	6787 => "00000000",
	6788 => "00000000",
	6789 => "00000000",
	6790 => "00000000",
	6791 => "00000000",
	6792 => "00000000",
	6793 => "00000000",
	6794 => "00000000",
	6795 => "00000000",
	6796 => "00000000",
	6797 => "00000000",
	6798 => "00000000",
	6799 => "00000000",
	6800 => "00000000",
	6801 => "00000000",
	6802 => "00000000",
	6803 => "00000000",
	6804 => "00000000",
	6805 => "00000000",
	6806 => "00000000",
	6807 => "00000000",
	6808 => "00000000",
	6809 => "00000000",
	6810 => "00000000",
	6811 => "00000000",
	6812 => "00000000",
	6813 => "00000000",
	6814 => "00000000",
	6815 => "00000000",
	6816 => "00000000",
	6817 => "00000000",
	6818 => "00000000",
	6819 => "00000000",
	6820 => "00000000",
	6821 => "00000000",
	6822 => "00000000",
	6823 => "00000000",
	6824 => "00000000",
	6825 => "00000000",
	6826 => "00000000",
	6827 => "00000000",
	6828 => "00000000",
	6829 => "00000000",
	6830 => "00000000",
	6831 => "00000000",
	6832 => "11111111",
	6833 => "11111111",
	6834 => "11111111",
	6835 => "11111111",
	6836 => "11111111",
	6837 => "11111111",
	6838 => "11111111",
	6839 => "11111111",
	6840 => "11111111",
	6841 => "11111111",
	6842 => "11111111",
	6843 => "00000000",
	6844 => "00000000",
	6845 => "00000000",
	6846 => "11111111",
	6847 => "11111111",
	6848 => "11111111",
	6849 => "11111111",
	6850 => "11111111",
	6851 => "11111111",
	6852 => "11111111",
	6853 => "11111111",
	6854 => "11111111",
	6855 => "11111111",
	6856 => "11111111",
	6857 => "00000000",
	6858 => "00000000",
	6859 => "00000000",
	6860 => "00000000",
	6861 => "00000000",
	6862 => "00000000",
	6863 => "00000000",
	6864 => "00000000",
	6865 => "00000000",
	6866 => "00000000",
	6867 => "00000000",
	6868 => "00000000",
	6869 => "00000000",
	6870 => "00000000",
	6871 => "00000000",
	6872 => "00000000",
	6873 => "00000000",
	6874 => "00000000",
	6875 => "00000000",
	6876 => "00000000",
	6877 => "00000000",
	6878 => "00000000",
	6879 => "00000000",
	6880 => "00000000",
	6881 => "00000000",
	6882 => "00000000",
	6883 => "00000000",
	6884 => "00000000",
	6885 => "00000000",
	6886 => "00000000",
	6887 => "00000000",
	6888 => "00000000",
	6889 => "00000000",
	6890 => "00000000",
	6891 => "00000000",
	6892 => "00000000",
	6893 => "00000000",
	6894 => "00000000",
	6895 => "00000000",
	6896 => "00000000",
	6897 => "00000000",
	6898 => "00000000",
	6899 => "00000000",
	6900 => "00000000",
	6901 => "00000000",
	6902 => "00000000",
	6903 => "00000000",
	6912 => "00000000",
	6913 => "00000000",
	6914 => "00000000",
	6915 => "00000000",
	6916 => "00000000",
	6917 => "00000000",
	6918 => "00000000",
	6919 => "00000000",
	6920 => "00000000",
	6921 => "00000000",
	6922 => "00000000",
	6923 => "00000000",
	6924 => "00000000",
	6925 => "00000000",
	6926 => "00000000",
	6927 => "00000000",
	6928 => "00000000",
	6929 => "00000000",
	6930 => "00000000",
	6931 => "00000000",
	6932 => "00000000",
	6933 => "00000000",
	6934 => "00000000",
	6935 => "00000000",
	6936 => "00000000",
	6937 => "00000000",
	6938 => "00000000",
	6939 => "00000000",
	6940 => "00000000",
	6941 => "00000000",
	6942 => "00000000",
	6943 => "00000000",
	6944 => "00000000",
	6945 => "00000000",
	6946 => "00000000",
	6947 => "00000000",
	6948 => "00000000",
	6949 => "00000000",
	6950 => "00000000",
	6951 => "00000000",
	6952 => "00000000",
	6953 => "00000000",
	6954 => "00000000",
	6955 => "00000000",
	6956 => "00000000",
	6957 => "00000000",
	6958 => "00000000",
	6959 => "00000000",
	6960 => "00000000",
	6961 => "11111111",
	6962 => "11111111",
	6963 => "11111111",
	6964 => "11111111",
	6965 => "11111111",
	6966 => "11111111",
	6967 => "11111111",
	6968 => "11111111",
	6969 => "11111111",
	6970 => "11111111",
	6971 => "11111111",
	6972 => "00000000",
	6973 => "11111111",
	6974 => "11111111",
	6975 => "11111111",
	6976 => "11111111",
	6977 => "11111111",
	6978 => "11111111",
	6979 => "11111111",
	6980 => "11111111",
	6981 => "11111111",
	6982 => "11111111",
	6983 => "11111111",
	6984 => "00000000",
	6985 => "00000000",
	6986 => "00000000",
	6987 => "00000000",
	6988 => "00000000",
	6989 => "00000000",
	6990 => "00000000",
	6991 => "00000000",
	6992 => "00000000",
	6993 => "00000000",
	6994 => "00000000",
	6995 => "00000000",
	6996 => "00000000",
	6997 => "00000000",
	6998 => "00000000",
	6999 => "00000000",
	7000 => "00000000",
	7001 => "00000000",
	7002 => "00000000",
	7003 => "00000000",
	7004 => "00000000",
	7005 => "00000000",
	7006 => "00000000",
	7007 => "00000000",
	7008 => "00000000",
	7009 => "00000000",
	7010 => "00000000",
	7011 => "00000000",
	7012 => "00000000",
	7013 => "00000000",
	7014 => "00000000",
	7015 => "00000000",
	7016 => "00000000",
	7017 => "00000000",
	7018 => "00000000",
	7019 => "00000000",
	7020 => "00000000",
	7021 => "00000000",
	7022 => "00000000",
	7023 => "00000000",
	7024 => "00000000",
	7025 => "00000000",
	7026 => "00000000",
	7027 => "00000000",
	7028 => "00000000",
	7029 => "00000000",
	7030 => "00000000",
	7031 => "00000000",
	7040 => "00000000",
	7041 => "00000000",
	7042 => "00000000",
	7043 => "00000000",
	7044 => "00000000",
	7045 => "00000000",
	7046 => "00000000",
	7047 => "00000000",
	7048 => "00000000",
	7049 => "00000000",
	7050 => "00000000",
	7051 => "00000000",
	7052 => "00000000",
	7053 => "00000000",
	7054 => "00000000",
	7055 => "00000000",
	7056 => "00000000",
	7057 => "00000000",
	7058 => "00000000",
	7059 => "00000000",
	7060 => "00000000",
	7061 => "00000000",
	7062 => "00000000",
	7063 => "00000000",
	7064 => "00000000",
	7065 => "00000000",
	7066 => "00000000",
	7067 => "00000000",
	7068 => "00000000",
	7069 => "00000000",
	7070 => "00000000",
	7071 => "00000000",
	7072 => "00000000",
	7073 => "00000000",
	7074 => "00000000",
	7075 => "00000000",
	7076 => "00000000",
	7077 => "00000000",
	7078 => "00000000",
	7079 => "00000000",
	7080 => "00000000",
	7081 => "00000000",
	7082 => "00000000",
	7083 => "00000000",
	7084 => "00000000",
	7085 => "00000000",
	7086 => "00000000",
	7087 => "00000000",
	7088 => "00000000",
	7089 => "00000000",
	7090 => "11111111",
	7091 => "11111111",
	7092 => "11111111",
	7093 => "11111111",
	7094 => "11111111",
	7095 => "11111111",
	7096 => "11111111",
	7097 => "11111111",
	7098 => "11111111",
	7099 => "11111111",
	7100 => "11111111",
	7101 => "11111111",
	7102 => "11111111",
	7103 => "11111111",
	7104 => "11111111",
	7105 => "11111111",
	7106 => "11111111",
	7107 => "11111111",
	7108 => "11111111",
	7109 => "11111111",
	7110 => "11111111",
	7111 => "00000000",
	7112 => "00000000",
	7113 => "00000000",
	7114 => "00000000",
	7115 => "00000000",
	7116 => "00000000",
	7117 => "00000000",
	7118 => "00000000",
	7119 => "00000000",
	7120 => "00000000",
	7121 => "00000000",
	7122 => "00000000",
	7123 => "00000000",
	7124 => "00000000",
	7125 => "00000000",
	7126 => "00000000",
	7127 => "00000000",
	7128 => "00000000",
	7129 => "00000000",
	7130 => "00000000",
	7131 => "00000000",
	7132 => "00000000",
	7133 => "00000000",
	7134 => "00000000",
	7135 => "00000000",
	7136 => "00000000",
	7137 => "00000000",
	7138 => "00000000",
	7139 => "00000000",
	7140 => "00000000",
	7141 => "00000000",
	7142 => "00000000",
	7143 => "00000000",
	7144 => "00000000",
	7145 => "00000000",
	7146 => "00000000",
	7147 => "00000000",
	7148 => "00000000",
	7149 => "00000000",
	7150 => "00000000",
	7151 => "00000000",
	7152 => "00000000",
	7153 => "00000000",
	7154 => "00000000",
	7155 => "00000000",
	7156 => "00000000",
	7157 => "00000000",
	7158 => "00000000",
	7159 => "00000000",
	7168 => "00000000",
	7169 => "00000000",
	7170 => "00000000",
	7171 => "00000000",
	7172 => "00000000",
	7173 => "00000000",
	7174 => "00000000",
	7175 => "00000000",
	7176 => "00000000",
	7177 => "00000000",
	7178 => "00000000",
	7179 => "00000000",
	7180 => "00000000",
	7181 => "00000000",
	7182 => "00000000",
	7183 => "00000000",
	7184 => "00000000",
	7185 => "00000000",
	7186 => "00000000",
	7187 => "00000000",
	7188 => "00000000",
	7189 => "00000000",
	7190 => "00000000",
	7191 => "00000000",
	7192 => "00000000",
	7193 => "00000000",
	7194 => "00000000",
	7195 => "00000000",
	7196 => "00000000",
	7197 => "00000000",
	7198 => "00000000",
	7199 => "00000000",
	7200 => "00000000",
	7201 => "00000000",
	7202 => "00000000",
	7203 => "00000000",
	7204 => "00000000",
	7205 => "00000000",
	7206 => "00000000",
	7207 => "00000000",
	7208 => "00000000",
	7209 => "00000000",
	7210 => "00000000",
	7211 => "00000000",
	7212 => "00000000",
	7213 => "00000000",
	7214 => "00000000",
	7215 => "00000000",
	7216 => "00000000",
	7217 => "00000000",
	7218 => "00000000",
	7219 => "11111111",
	7220 => "11111111",
	7221 => "11111111",
	7222 => "11111111",
	7223 => "11111111",
	7224 => "11111111",
	7225 => "11111111",
	7226 => "11111111",
	7227 => "11111111",
	7228 => "11111111",
	7229 => "11111111",
	7230 => "11111111",
	7231 => "11111111",
	7232 => "11111111",
	7233 => "11111111",
	7234 => "11111111",
	7235 => "11111111",
	7236 => "11111111",
	7237 => "11111111",
	7238 => "00000000",
	7239 => "00000000",
	7240 => "00000000",
	7241 => "00000000",
	7242 => "00000000",
	7243 => "00000000",
	7244 => "00000000",
	7245 => "00000000",
	7246 => "00000000",
	7247 => "00000000",
	7248 => "00000000",
	7249 => "00000000",
	7250 => "00000000",
	7251 => "00000000",
	7252 => "00000000",
	7253 => "00000000",
	7254 => "00000000",
	7255 => "00000000",
	7256 => "00000000",
	7257 => "00000000",
	7258 => "00000000",
	7259 => "00000000",
	7260 => "00000000",
	7261 => "00000000",
	7262 => "00000000",
	7263 => "00000000",
	7264 => "00000000",
	7265 => "00000000",
	7266 => "00000000",
	7267 => "00000000",
	7268 => "00000000",
	7269 => "00000000",
	7270 => "00000000",
	7271 => "00000000",
	7272 => "00000000",
	7273 => "00000000",
	7274 => "00000000",
	7275 => "00000000",
	7276 => "00000000",
	7277 => "00000000",
	7278 => "00000000",
	7279 => "00000000",
	7280 => "00000000",
	7281 => "00000000",
	7282 => "00000000",
	7283 => "00000000",
	7284 => "00000000",
	7285 => "00000000",
	7286 => "00000000",
	7287 => "00000000",
	7296 => "00000000",
	7297 => "00000000",
	7298 => "00000000",
	7299 => "00000000",
	7300 => "00000000",
	7301 => "00000000",
	7302 => "00000000",
	7303 => "00000000",
	7304 => "00000000",
	7305 => "00000000",
	7306 => "00000000",
	7307 => "00000000",
	7308 => "00000000",
	7309 => "00000000",
	7310 => "00000000",
	7311 => "00000000",
	7312 => "00000000",
	7313 => "00000000",
	7314 => "00000000",
	7315 => "00000000",
	7316 => "00000000",
	7317 => "00000000",
	7318 => "00000000",
	7319 => "00000000",
	7320 => "00000000",
	7321 => "00000000",
	7322 => "00000000",
	7323 => "00000000",
	7324 => "00000000",
	7325 => "00000000",
	7326 => "00000000",
	7327 => "00000000",
	7328 => "00000000",
	7329 => "00000000",
	7330 => "00000000",
	7331 => "00000000",
	7332 => "00000000",
	7333 => "00000000",
	7334 => "00000000",
	7335 => "00000000",
	7336 => "00000000",
	7337 => "00000000",
	7338 => "00000000",
	7339 => "00000000",
	7340 => "00000000",
	7341 => "00000000",
	7342 => "00000000",
	7343 => "00000000",
	7344 => "00000000",
	7345 => "00000000",
	7346 => "00000000",
	7347 => "00000000",
	7348 => "11111111",
	7349 => "11111111",
	7350 => "11111111",
	7351 => "11111111",
	7352 => "11111111",
	7353 => "11111111",
	7354 => "11111111",
	7355 => "11111111",
	7356 => "11111111",
	7357 => "11111111",
	7358 => "11111111",
	7359 => "11111111",
	7360 => "11111111",
	7361 => "11111111",
	7362 => "11111111",
	7363 => "11111111",
	7364 => "11111111",
	7365 => "00000000",
	7366 => "00000000",
	7367 => "00000000",
	7368 => "00000000",
	7369 => "00000000",
	7370 => "00000000",
	7371 => "00000000",
	7372 => "00000000",
	7373 => "00000000",
	7374 => "00000000",
	7375 => "00000000",
	7376 => "00000000",
	7377 => "00000000",
	7378 => "00000000",
	7379 => "00000000",
	7380 => "00000000",
	7381 => "00000000",
	7382 => "00000000",
	7383 => "00000000",
	7384 => "00000000",
	7385 => "00000000",
	7386 => "00000000",
	7387 => "00000000",
	7388 => "00000000",
	7389 => "00000000",
	7390 => "00000000",
	7391 => "00000000",
	7392 => "00000000",
	7393 => "00000000",
	7394 => "00000000",
	7395 => "00000000",
	7396 => "00000000",
	7397 => "00000000",
	7398 => "00000000",
	7399 => "00000000",
	7400 => "00000000",
	7401 => "00000000",
	7402 => "00000000",
	7403 => "00000000",
	7404 => "00000000",
	7405 => "00000000",
	7406 => "00000000",
	7407 => "00000000",
	7408 => "00000000",
	7409 => "00000000",
	7410 => "00000000",
	7411 => "00000000",
	7412 => "00000000",
	7413 => "00000000",
	7414 => "00000000",
	7415 => "00000000",
	7424 => "00000000",
	7425 => "00000000",
	7426 => "00000000",
	7427 => "00000000",
	7428 => "00000000",
	7429 => "00000000",
	7430 => "00000000",
	7431 => "00000000",
	7432 => "00000000",
	7433 => "00000000",
	7434 => "00000000",
	7435 => "00000000",
	7436 => "00000000",
	7437 => "00000000",
	7438 => "00000000",
	7439 => "00000000",
	7440 => "00000000",
	7441 => "00000000",
	7442 => "00000000",
	7443 => "00000000",
	7444 => "00000000",
	7445 => "00000000",
	7446 => "00000000",
	7447 => "00000000",
	7448 => "00000000",
	7449 => "00000000",
	7450 => "00000000",
	7451 => "00000000",
	7452 => "00000000",
	7453 => "00000000",
	7454 => "00000000",
	7455 => "00000000",
	7456 => "00000000",
	7457 => "00000000",
	7458 => "00000000",
	7459 => "00000000",
	7460 => "00000000",
	7461 => "00000000",
	7462 => "00000000",
	7463 => "00000000",
	7464 => "00000000",
	7465 => "00000000",
	7466 => "00000000",
	7467 => "00000000",
	7468 => "00000000",
	7469 => "00000000",
	7470 => "00000000",
	7471 => "00000000",
	7472 => "00000000",
	7473 => "00000000",
	7474 => "00000000",
	7475 => "00000000",
	7476 => "00000000",
	7477 => "11111111",
	7478 => "11111111",
	7479 => "11111111",
	7480 => "11111111",
	7481 => "11111111",
	7482 => "11111111",
	7483 => "11111111",
	7484 => "11111111",
	7485 => "11111111",
	7486 => "11111111",
	7487 => "11111111",
	7488 => "11111111",
	7489 => "11111111",
	7490 => "11111111",
	7491 => "11111111",
	7492 => "00000000",
	7493 => "00000000",
	7494 => "00000000",
	7495 => "00000000",
	7496 => "00000000",
	7497 => "00000000",
	7498 => "00000000",
	7499 => "00000000",
	7500 => "00000000",
	7501 => "00000000",
	7502 => "00000000",
	7503 => "00000000",
	7504 => "00000000",
	7505 => "00000000",
	7506 => "00000000",
	7507 => "00000000",
	7508 => "00000000",
	7509 => "00000000",
	7510 => "00000000",
	7511 => "00000000",
	7512 => "00000000",
	7513 => "00000000",
	7514 => "00000000",
	7515 => "00000000",
	7516 => "00000000",
	7517 => "00000000",
	7518 => "00000000",
	7519 => "00000000",
	7520 => "00000000",
	7521 => "00000000",
	7522 => "00000000",
	7523 => "00000000",
	7524 => "00000000",
	7525 => "00000000",
	7526 => "00000000",
	7527 => "00000000",
	7528 => "00000000",
	7529 => "00000000",
	7530 => "00000000",
	7531 => "00000000",
	7532 => "00000000",
	7533 => "00000000",
	7534 => "00000000",
	7535 => "00000000",
	7536 => "00000000",
	7537 => "00000000",
	7538 => "00000000",
	7539 => "00000000",
	7540 => "00000000",
	7541 => "00000000",
	7542 => "00000000",
	7543 => "00000000",
	7552 => "00000000",
	7553 => "00000000",
	7554 => "00000000",
	7555 => "00000000",
	7556 => "00000000",
	7557 => "00000000",
	7558 => "00000000",
	7559 => "00000000",
	7560 => "00000000",
	7561 => "00000000",
	7562 => "00000000",
	7563 => "00000000",
	7564 => "00000000",
	7565 => "00000000",
	7566 => "00000000",
	7567 => "00000000",
	7568 => "00000000",
	7569 => "00000000",
	7570 => "00000000",
	7571 => "00000000",
	7572 => "00000000",
	7573 => "00000000",
	7574 => "00000000",
	7575 => "00000000",
	7576 => "00000000",
	7577 => "00000000",
	7578 => "00000000",
	7579 => "00000000",
	7580 => "00000000",
	7581 => "00000000",
	7582 => "00000000",
	7583 => "00000000",
	7584 => "00000000",
	7585 => "00000000",
	7586 => "00000000",
	7587 => "00000000",
	7588 => "00000000",
	7589 => "00000000",
	7590 => "00000000",
	7591 => "00000000",
	7592 => "00000000",
	7593 => "00000000",
	7594 => "00000000",
	7595 => "00000000",
	7596 => "00000000",
	7597 => "00000000",
	7598 => "00000000",
	7599 => "00000000",
	7600 => "00000000",
	7601 => "00000000",
	7602 => "00000000",
	7603 => "00000000",
	7604 => "00000000",
	7605 => "00000000",
	7606 => "11111111",
	7607 => "11111111",
	7608 => "11111111",
	7609 => "11111111",
	7610 => "11111111",
	7611 => "11111111",
	7612 => "11111111",
	7613 => "11111111",
	7614 => "11111111",
	7615 => "11111111",
	7616 => "11111111",
	7617 => "11111111",
	7618 => "11111111",
	7619 => "00000000",
	7620 => "00000000",
	7621 => "00000000",
	7622 => "00000000",
	7623 => "00000000",
	7624 => "00000000",
	7625 => "00000000",
	7626 => "00000000",
	7627 => "00000000",
	7628 => "00000000",
	7629 => "00000000",
	7630 => "00000000",
	7631 => "00000000",
	7632 => "00000000",
	7633 => "00000000",
	7634 => "00000000",
	7635 => "00000000",
	7636 => "00000000",
	7637 => "00000000",
	7638 => "00000000",
	7639 => "00000000",
	7640 => "00000000",
	7641 => "00000000",
	7642 => "00000000",
	7643 => "00000000",
	7644 => "00000000",
	7645 => "00000000",
	7646 => "00000000",
	7647 => "00000000",
	7648 => "00000000",
	7649 => "00000000",
	7650 => "00000000",
	7651 => "00000000",
	7652 => "00000000",
	7653 => "00000000",
	7654 => "00000000",
	7655 => "00000000",
	7656 => "00000000",
	7657 => "00000000",
	7658 => "00000000",
	7659 => "00000000",
	7660 => "00000000",
	7661 => "00000000",
	7662 => "00000000",
	7663 => "00000000",
	7664 => "00000000",
	7665 => "00000000",
	7666 => "00000000",
	7667 => "00000000",
	7668 => "00000000",
	7669 => "00000000",
	7670 => "00000000",
	7671 => "00000000",
	7680 => "00000000",
	7681 => "00000000",
	7682 => "00000000",
	7683 => "00000000",
	7684 => "00000000",
	7685 => "00000000",
	7686 => "00000000",
	7687 => "00000000",
	7688 => "00000000",
	7689 => "00000000",
	7690 => "00000000",
	7691 => "00000000",
	7692 => "00000000",
	7693 => "00000000",
	7694 => "00000000",
	7695 => "00000000",
	7696 => "00000000",
	7697 => "00000000",
	7698 => "00000000",
	7699 => "00000000",
	7700 => "00000000",
	7701 => "00000000",
	7702 => "00000000",
	7703 => "00000000",
	7704 => "00000000",
	7705 => "00000000",
	7706 => "00000000",
	7707 => "00000000",
	7708 => "00000000",
	7709 => "00000000",
	7710 => "00000000",
	7711 => "00000000",
	7712 => "00000000",
	7713 => "00000000",
	7714 => "00000000",
	7715 => "00000000",
	7716 => "00000000",
	7717 => "00000000",
	7718 => "00000000",
	7719 => "00000000",
	7720 => "00000000",
	7721 => "00000000",
	7722 => "00000000",
	7723 => "00000000",
	7724 => "00000000",
	7725 => "00000000",
	7726 => "00000000",
	7727 => "00000000",
	7728 => "00000000",
	7729 => "00000000",
	7730 => "00000000",
	7731 => "00000000",
	7732 => "00000000",
	7733 => "00000000",
	7734 => "00000000",
	7735 => "11111111",
	7736 => "11111111",
	7737 => "11111111",
	7738 => "11111111",
	7739 => "11111111",
	7740 => "11111111",
	7741 => "11111111",
	7742 => "11111111",
	7743 => "11111111",
	7744 => "11111111",
	7745 => "11111111",
	7746 => "00000000",
	7747 => "00000000",
	7748 => "00000000",
	7749 => "00000000",
	7750 => "00000000",
	7751 => "00000000",
	7752 => "00000000",
	7753 => "00000000",
	7754 => "00000000",
	7755 => "00000000",
	7756 => "00000000",
	7757 => "00000000",
	7758 => "00000000",
	7759 => "00000000",
	7760 => "00000000",
	7761 => "00000000",
	7762 => "00000000",
	7763 => "00000000",
	7764 => "00000000",
	7765 => "00000000",
	7766 => "00000000",
	7767 => "00000000",
	7768 => "00000000",
	7769 => "00000000",
	7770 => "00000000",
	7771 => "00000000",
	7772 => "00000000",
	7773 => "00000000",
	7774 => "00000000",
	7775 => "00000000",
	7776 => "00000000",
	7777 => "00000000",
	7778 => "00000000",
	7779 => "00000000",
	7780 => "00000000",
	7781 => "00000000",
	7782 => "00000000",
	7783 => "00000000",
	7784 => "00000000",
	7785 => "00000000",
	7786 => "00000000",
	7787 => "00000000",
	7788 => "00000000",
	7789 => "00000000",
	7790 => "00000000",
	7791 => "00000000",
	7792 => "00000000",
	7793 => "00000000",
	7794 => "00000000",
	7795 => "00000000",
	7796 => "00000000",
	7797 => "00000000",
	7798 => "00000000",
	7799 => "00000000",
	7808 => "00000000",
	7809 => "00000000",
	7810 => "00000000",
	7811 => "00000000",
	7812 => "00000000",
	7813 => "00000000",
	7814 => "00000000",
	7815 => "00000000",
	7816 => "00000000",
	7817 => "00000000",
	7818 => "00000000",
	7819 => "00000000",
	7820 => "00000000",
	7821 => "00000000",
	7822 => "00000000",
	7823 => "00000000",
	7824 => "00000000",
	7825 => "00000000",
	7826 => "00000000",
	7827 => "00000000",
	7828 => "00000000",
	7829 => "00000000",
	7830 => "00000000",
	7831 => "00000000",
	7832 => "00000000",
	7833 => "00000000",
	7834 => "00000000",
	7835 => "00000000",
	7836 => "00000000",
	7837 => "00000000",
	7838 => "00000000",
	7839 => "00000000",
	7840 => "00000000",
	7841 => "00000000",
	7842 => "00000000",
	7843 => "00000000",
	7844 => "00000000",
	7845 => "00000000",
	7846 => "00000000",
	7847 => "00000000",
	7848 => "00000000",
	7849 => "00000000",
	7850 => "00000000",
	7851 => "00000000",
	7852 => "00000000",
	7853 => "00000000",
	7854 => "00000000",
	7855 => "00000000",
	7856 => "00000000",
	7857 => "00000000",
	7858 => "00000000",
	7859 => "00000000",
	7860 => "00000000",
	7861 => "00000000",
	7862 => "11111111",
	7863 => "11111111",
	7864 => "11111111",
	7865 => "11111111",
	7866 => "11111111",
	7867 => "11111111",
	7868 => "11111111",
	7869 => "11111111",
	7870 => "11111111",
	7871 => "11111111",
	7872 => "11111111",
	7873 => "11111111",
	7874 => "11111111",
	7875 => "00000000",
	7876 => "00000000",
	7877 => "00000000",
	7878 => "00000000",
	7879 => "00000000",
	7880 => "00000000",
	7881 => "00000000",
	7882 => "00000000",
	7883 => "00000000",
	7884 => "00000000",
	7885 => "00000000",
	7886 => "00000000",
	7887 => "00000000",
	7888 => "00000000",
	7889 => "00000000",
	7890 => "00000000",
	7891 => "00000000",
	7892 => "00000000",
	7893 => "00000000",
	7894 => "00000000",
	7895 => "00000000",
	7896 => "00000000",
	7897 => "00000000",
	7898 => "00000000",
	7899 => "00000000",
	7900 => "00000000",
	7901 => "00000000",
	7902 => "00000000",
	7903 => "00000000",
	7904 => "00000000",
	7905 => "00000000",
	7906 => "00000000",
	7907 => "00000000",
	7908 => "00000000",
	7909 => "00000000",
	7910 => "00000000",
	7911 => "00000000",
	7912 => "00000000",
	7913 => "00000000",
	7914 => "00000000",
	7915 => "00000000",
	7916 => "00000000",
	7917 => "00000000",
	7918 => "00000000",
	7919 => "00000000",
	7920 => "00000000",
	7921 => "00000000",
	7922 => "00000000",
	7923 => "00000000",
	7924 => "00000000",
	7925 => "00000000",
	7926 => "00000000",
	7927 => "00000000",
	7936 => "00000000",
	7937 => "00000000",
	7938 => "00000000",
	7939 => "00000000",
	7940 => "00000000",
	7941 => "00000000",
	7942 => "00000000",
	7943 => "00000000",
	7944 => "00000000",
	7945 => "00000000",
	7946 => "00000000",
	7947 => "00000000",
	7948 => "00000000",
	7949 => "00000000",
	7950 => "00000000",
	7951 => "00000000",
	7952 => "00000000",
	7953 => "00000000",
	7954 => "00000000",
	7955 => "00000000",
	7956 => "00000000",
	7957 => "00000000",
	7958 => "00000000",
	7959 => "00000000",
	7960 => "00000000",
	7961 => "00000000",
	7962 => "00000000",
	7963 => "00000000",
	7964 => "00000000",
	7965 => "00000000",
	7966 => "00000000",
	7967 => "00000000",
	7968 => "00000000",
	7969 => "00000000",
	7970 => "00000000",
	7971 => "00000000",
	7972 => "00000000",
	7973 => "00000000",
	7974 => "00000000",
	7975 => "00000000",
	7976 => "00000000",
	7977 => "00000000",
	7978 => "00000000",
	7979 => "00000000",
	7980 => "00000000",
	7981 => "00000000",
	7982 => "00000000",
	7983 => "00000000",
	7984 => "00000000",
	7985 => "00000000",
	7986 => "00000000",
	7987 => "00000000",
	7988 => "00000000",
	7989 => "11111111",
	7990 => "11111111",
	7991 => "11111111",
	7992 => "11111111",
	7993 => "11111111",
	7994 => "11111111",
	7995 => "11111111",
	7996 => "11111111",
	7997 => "11111111",
	7998 => "11111111",
	7999 => "11111111",
	8000 => "11111111",
	8001 => "11111111",
	8002 => "11111111",
	8003 => "11111111",
	8004 => "00000000",
	8005 => "00000000",
	8006 => "00000000",
	8007 => "00000000",
	8008 => "00000000",
	8009 => "00000000",
	8010 => "00000000",
	8011 => "00000000",
	8012 => "00000000",
	8013 => "00000000",
	8014 => "00000000",
	8015 => "00000000",
	8016 => "00000000",
	8017 => "00000000",
	8018 => "00000000",
	8019 => "00000000",
	8020 => "00000000",
	8021 => "00000000",
	8022 => "00000000",
	8023 => "00000000",
	8024 => "00000000",
	8025 => "00000000",
	8026 => "00000000",
	8027 => "00000000",
	8028 => "00000000",
	8029 => "00000000",
	8030 => "00000000",
	8031 => "00000000",
	8032 => "00000000",
	8033 => "00000000",
	8034 => "00000000",
	8035 => "00000000",
	8036 => "00000000",
	8037 => "00000000",
	8038 => "00000000",
	8039 => "00000000",
	8040 => "00000000",
	8041 => "00000000",
	8042 => "00000000",
	8043 => "00000000",
	8044 => "00000000",
	8045 => "00000000",
	8046 => "00000000",
	8047 => "00000000",
	8048 => "00000000",
	8049 => "00000000",
	8050 => "00000000",
	8051 => "00000000",
	8052 => "00000000",
	8053 => "00000000",
	8054 => "00000000",
	8055 => "00000000",
	8064 => "00000000",
	8065 => "00000000",
	8066 => "00000000",
	8067 => "00000000",
	8068 => "00000000",
	8069 => "00000000",
	8070 => "00000000",
	8071 => "00000000",
	8072 => "00000000",
	8073 => "00000000",
	8074 => "00000000",
	8075 => "00000000",
	8076 => "00000000",
	8077 => "00000000",
	8078 => "00000000",
	8079 => "00000000",
	8080 => "00000000",
	8081 => "00000000",
	8082 => "00000000",
	8083 => "00000000",
	8084 => "00000000",
	8085 => "00000000",
	8086 => "00000000",
	8087 => "00000000",
	8088 => "00000000",
	8089 => "00000000",
	8090 => "00000000",
	8091 => "00000000",
	8092 => "00000000",
	8093 => "00000000",
	8094 => "00000000",
	8095 => "00000000",
	8096 => "00000000",
	8097 => "00000000",
	8098 => "00000000",
	8099 => "00000000",
	8100 => "00000000",
	8101 => "00000000",
	8102 => "00000000",
	8103 => "00000000",
	8104 => "00000000",
	8105 => "00000000",
	8106 => "00000000",
	8107 => "00000000",
	8108 => "00000000",
	8109 => "00000000",
	8110 => "00000000",
	8111 => "00000000",
	8112 => "00000000",
	8113 => "00000000",
	8114 => "00000000",
	8115 => "00000000",
	8116 => "11111111",
	8117 => "11111111",
	8118 => "11111111",
	8119 => "11111111",
	8120 => "11111111",
	8121 => "11111111",
	8122 => "11111111",
	8123 => "11111111",
	8124 => "11111111",
	8125 => "11111111",
	8126 => "11111111",
	8127 => "11111111",
	8128 => "11111111",
	8129 => "11111111",
	8130 => "11111111",
	8131 => "11111111",
	8132 => "11111111",
	8133 => "00000000",
	8134 => "00000000",
	8135 => "00000000",
	8136 => "00000000",
	8137 => "00000000",
	8138 => "00000000",
	8139 => "00000000",
	8140 => "00000000",
	8141 => "00000000",
	8142 => "00000000",
	8143 => "00000000",
	8144 => "00000000",
	8145 => "00000000",
	8146 => "00000000",
	8147 => "00000000",
	8148 => "00000000",
	8149 => "00000000",
	8150 => "00000000",
	8151 => "00000000",
	8152 => "00000000",
	8153 => "00000000",
	8154 => "00000000",
	8155 => "00000000",
	8156 => "00000000",
	8157 => "00000000",
	8158 => "00000000",
	8159 => "00000000",
	8160 => "00000000",
	8161 => "00000000",
	8162 => "00000000",
	8163 => "00000000",
	8164 => "00000000",
	8165 => "00000000",
	8166 => "00000000",
	8167 => "00000000",
	8168 => "00000000",
	8169 => "00000000",
	8170 => "00000000",
	8171 => "00000000",
	8172 => "00000000",
	8173 => "00000000",
	8174 => "00000000",
	8175 => "00000000",
	8176 => "00000000",
	8177 => "00000000",
	8178 => "00000000",
	8179 => "00000000",
	8180 => "00000000",
	8181 => "00000000",
	8182 => "00000000",
	8183 => "00000000",
	8192 => "00000000",
	8193 => "00000000",
	8194 => "00000000",
	8195 => "00000000",
	8196 => "00000000",
	8197 => "00000000",
	8198 => "00000000",
	8199 => "00000000",
	8200 => "00000000",
	8201 => "00000000",
	8202 => "00000000",
	8203 => "00000000",
	8204 => "00000000",
	8205 => "00000000",
	8206 => "00000000",
	8207 => "00000000",
	8208 => "00000000",
	8209 => "00000000",
	8210 => "00000000",
	8211 => "00000000",
	8212 => "00000000",
	8213 => "00000000",
	8214 => "00000000",
	8215 => "00000000",
	8216 => "00000000",
	8217 => "00000000",
	8218 => "00000000",
	8219 => "00000000",
	8220 => "00000000",
	8221 => "00000000",
	8222 => "00000000",
	8223 => "00000000",
	8224 => "00000000",
	8225 => "00000000",
	8226 => "00000000",
	8227 => "00000000",
	8228 => "00000000",
	8229 => "00000000",
	8230 => "00000000",
	8231 => "00000000",
	8232 => "00000000",
	8233 => "00000000",
	8234 => "00000000",
	8235 => "00000000",
	8236 => "00000000",
	8237 => "00000000",
	8238 => "00000000",
	8239 => "00000000",
	8240 => "00000000",
	8241 => "00000000",
	8242 => "00000000",
	8243 => "11111111",
	8244 => "11111111",
	8245 => "11111111",
	8246 => "11111111",
	8247 => "11111111",
	8248 => "11111111",
	8249 => "11111111",
	8250 => "11111111",
	8251 => "11111111",
	8252 => "11111111",
	8253 => "11111111",
	8254 => "11111111",
	8255 => "11111111",
	8256 => "11111111",
	8257 => "11111111",
	8258 => "11111111",
	8259 => "11111111",
	8260 => "11111111",
	8261 => "11111111",
	8262 => "00000000",
	8263 => "00000000",
	8264 => "00000000",
	8265 => "00000000",
	8266 => "00000000",
	8267 => "00000000",
	8268 => "00000000",
	8269 => "00000000",
	8270 => "00000000",
	8271 => "00000000",
	8272 => "00000000",
	8273 => "00000000",
	8274 => "00000000",
	8275 => "00000000",
	8276 => "00000000",
	8277 => "00000000",
	8278 => "00000000",
	8279 => "00000000",
	8280 => "00000000",
	8281 => "00000000",
	8282 => "00000000",
	8283 => "00000000",
	8284 => "00000000",
	8285 => "00000000",
	8286 => "00000000",
	8287 => "00000000",
	8288 => "00000000",
	8289 => "00000000",
	8290 => "00000000",
	8291 => "00000000",
	8292 => "00000000",
	8293 => "00000000",
	8294 => "00000000",
	8295 => "00000000",
	8296 => "00000000",
	8297 => "00000000",
	8298 => "00000000",
	8299 => "00000000",
	8300 => "00000000",
	8301 => "00000000",
	8302 => "00000000",
	8303 => "00000000",
	8304 => "00000000",
	8305 => "00000000",
	8306 => "00000000",
	8307 => "00000000",
	8308 => "00000000",
	8309 => "00000000",
	8310 => "00000000",
	8311 => "00000000",
	8320 => "00000000",
	8321 => "00000000",
	8322 => "00000000",
	8323 => "00000000",
	8324 => "00000000",
	8325 => "00000000",
	8326 => "00000000",
	8327 => "00000000",
	8328 => "00000000",
	8329 => "00000000",
	8330 => "00000000",
	8331 => "00000000",
	8332 => "00000000",
	8333 => "00000000",
	8334 => "00000000",
	8335 => "00000000",
	8336 => "00000000",
	8337 => "00000000",
	8338 => "00000000",
	8339 => "00000000",
	8340 => "00000000",
	8341 => "00000000",
	8342 => "00000000",
	8343 => "00000000",
	8344 => "00000000",
	8345 => "00000000",
	8346 => "00000000",
	8347 => "00000000",
	8348 => "00000000",
	8349 => "00000000",
	8350 => "00000000",
	8351 => "00000000",
	8352 => "00000000",
	8353 => "00000000",
	8354 => "00000000",
	8355 => "00000000",
	8356 => "00000000",
	8357 => "00000000",
	8358 => "00000000",
	8359 => "00000000",
	8360 => "00000000",
	8361 => "00000000",
	8362 => "00000000",
	8363 => "00000000",
	8364 => "00000000",
	8365 => "00000000",
	8366 => "00000000",
	8367 => "00000000",
	8368 => "00000000",
	8369 => "00000000",
	8370 => "11111111",
	8371 => "11111111",
	8372 => "11111111",
	8373 => "11111111",
	8374 => "11111111",
	8375 => "11111111",
	8376 => "11111111",
	8377 => "11111111",
	8378 => "11111111",
	8379 => "11111111",
	8380 => "11111111",
	8381 => "11111111",
	8382 => "11111111",
	8383 => "11111111",
	8384 => "11111111",
	8385 => "11111111",
	8386 => "11111111",
	8387 => "11111111",
	8388 => "11111111",
	8389 => "11111111",
	8390 => "11111111",
	8391 => "00000000",
	8392 => "00000000",
	8393 => "00000000",
	8394 => "00000000",
	8395 => "00000000",
	8396 => "00000000",
	8397 => "00000000",
	8398 => "00000000",
	8399 => "00000000",
	8400 => "00000000",
	8401 => "00000000",
	8402 => "00000000",
	8403 => "00000000",
	8404 => "00000000",
	8405 => "00000000",
	8406 => "00000000",
	8407 => "00000000",
	8408 => "00000000",
	8409 => "00000000",
	8410 => "00000000",
	8411 => "00000000",
	8412 => "00000000",
	8413 => "00000000",
	8414 => "00000000",
	8415 => "00000000",
	8416 => "00000000",
	8417 => "00000000",
	8418 => "00000000",
	8419 => "00000000",
	8420 => "00000000",
	8421 => "00000000",
	8422 => "00000000",
	8423 => "00000000",
	8424 => "00000000",
	8425 => "00000000",
	8426 => "00000000",
	8427 => "00000000",
	8428 => "00000000",
	8429 => "00000000",
	8430 => "00000000",
	8431 => "00000000",
	8432 => "00000000",
	8433 => "00000000",
	8434 => "00000000",
	8435 => "00000000",
	8436 => "00000000",
	8437 => "00000000",
	8438 => "00000000",
	8439 => "00000000",
	8448 => "00000000",
	8449 => "00000000",
	8450 => "00000000",
	8451 => "00000000",
	8452 => "00000000",
	8453 => "00000000",
	8454 => "00000000",
	8455 => "00000000",
	8456 => "00000000",
	8457 => "00000000",
	8458 => "00000000",
	8459 => "00000000",
	8460 => "00000000",
	8461 => "00000000",
	8462 => "00000000",
	8463 => "00000000",
	8464 => "00000000",
	8465 => "00000000",
	8466 => "00000000",
	8467 => "00000000",
	8468 => "00000000",
	8469 => "00000000",
	8470 => "00000000",
	8471 => "00000000",
	8472 => "00000000",
	8473 => "00000000",
	8474 => "00000000",
	8475 => "00000000",
	8476 => "00000000",
	8477 => "00000000",
	8478 => "00000000",
	8479 => "00000000",
	8480 => "00000000",
	8481 => "00000000",
	8482 => "00000000",
	8483 => "00000000",
	8484 => "00000000",
	8485 => "00000000",
	8486 => "00000000",
	8487 => "00000000",
	8488 => "00000000",
	8489 => "00000000",
	8490 => "00000000",
	8491 => "00000000",
	8492 => "00000000",
	8493 => "00000000",
	8494 => "00000000",
	8495 => "00000000",
	8496 => "00000000",
	8497 => "11111111",
	8498 => "11111111",
	8499 => "11111111",
	8500 => "11111111",
	8501 => "11111111",
	8502 => "11111111",
	8503 => "11111111",
	8504 => "11111111",
	8505 => "11111111",
	8506 => "11111111",
	8507 => "11111111",
	8508 => "00000000",
	8509 => "11111111",
	8510 => "11111111",
	8511 => "11111111",
	8512 => "11111111",
	8513 => "11111111",
	8514 => "11111111",
	8515 => "11111111",
	8516 => "11111111",
	8517 => "11111111",
	8518 => "11111111",
	8519 => "11111111",
	8520 => "00000000",
	8521 => "00000000",
	8522 => "00000000",
	8523 => "00000000",
	8524 => "00000000",
	8525 => "00000000",
	8526 => "00000000",
	8527 => "00000000",
	8528 => "00000000",
	8529 => "00000000",
	8530 => "00000000",
	8531 => "00000000",
	8532 => "00000000",
	8533 => "00000000",
	8534 => "00000000",
	8535 => "00000000",
	8536 => "00000000",
	8537 => "00000000",
	8538 => "00000000",
	8539 => "00000000",
	8540 => "00000000",
	8541 => "00000000",
	8542 => "00000000",
	8543 => "00000000",
	8544 => "00000000",
	8545 => "00000000",
	8546 => "00000000",
	8547 => "00000000",
	8548 => "00000000",
	8549 => "00000000",
	8550 => "00000000",
	8551 => "00000000",
	8552 => "00000000",
	8553 => "00000000",
	8554 => "00000000",
	8555 => "00000000",
	8556 => "00000000",
	8557 => "00000000",
	8558 => "00000000",
	8559 => "00000000",
	8560 => "00000000",
	8561 => "00000000",
	8562 => "00000000",
	8563 => "00000000",
	8564 => "00000000",
	8565 => "00000000",
	8566 => "00000000",
	8567 => "00000000",
	8576 => "00000000",
	8577 => "00000000",
	8578 => "00000000",
	8579 => "00000000",
	8580 => "00000000",
	8581 => "00000000",
	8582 => "00000000",
	8583 => "00000000",
	8584 => "00000000",
	8585 => "00000000",
	8586 => "00000000",
	8587 => "00000000",
	8588 => "00000000",
	8589 => "00000000",
	8590 => "00000000",
	8591 => "00000000",
	8592 => "00000000",
	8593 => "00000000",
	8594 => "00000000",
	8595 => "00000000",
	8596 => "00000000",
	8597 => "00000000",
	8598 => "00000000",
	8599 => "00000000",
	8600 => "00000000",
	8601 => "00000000",
	8602 => "00000000",
	8603 => "00000000",
	8604 => "00000000",
	8605 => "00000000",
	8606 => "00000000",
	8607 => "00000000",
	8608 => "00000000",
	8609 => "00000000",
	8610 => "00000000",
	8611 => "00000000",
	8612 => "00000000",
	8613 => "00000000",
	8614 => "00000000",
	8615 => "00000000",
	8616 => "00000000",
	8617 => "00000000",
	8618 => "00000000",
	8619 => "00000000",
	8620 => "00000000",
	8621 => "00000000",
	8622 => "00000000",
	8623 => "00000000",
	8624 => "11111111",
	8625 => "11111111",
	8626 => "11111111",
	8627 => "11111111",
	8628 => "11111111",
	8629 => "11111111",
	8630 => "11111111",
	8631 => "11111111",
	8632 => "11111111",
	8633 => "11111111",
	8634 => "11111111",
	8635 => "00000000",
	8636 => "00000000",
	8637 => "00000000",
	8638 => "11111111",
	8639 => "11111111",
	8640 => "11111111",
	8641 => "11111111",
	8642 => "11111111",
	8643 => "11111111",
	8644 => "11111111",
	8645 => "11111111",
	8646 => "11111111",
	8647 => "11111111",
	8648 => "11111111",
	8649 => "00000000",
	8650 => "00000000",
	8651 => "00000000",
	8652 => "00000000",
	8653 => "00000000",
	8654 => "00000000",
	8655 => "00000000",
	8656 => "00000000",
	8657 => "00000000",
	8658 => "00000000",
	8659 => "00000000",
	8660 => "00000000",
	8661 => "00000000",
	8662 => "00000000",
	8663 => "00000000",
	8664 => "00000000",
	8665 => "00000000",
	8666 => "00000000",
	8667 => "00000000",
	8668 => "00000000",
	8669 => "00000000",
	8670 => "00000000",
	8671 => "00000000",
	8672 => "00000000",
	8673 => "00000000",
	8674 => "00000000",
	8675 => "00000000",
	8676 => "00000000",
	8677 => "00000000",
	8678 => "00000000",
	8679 => "00000000",
	8680 => "00000000",
	8681 => "00000000",
	8682 => "00000000",
	8683 => "00000000",
	8684 => "00000000",
	8685 => "00000000",
	8686 => "00000000",
	8687 => "00000000",
	8688 => "00000000",
	8689 => "00000000",
	8690 => "00000000",
	8691 => "00000000",
	8692 => "00000000",
	8693 => "00000000",
	8694 => "00000000",
	8695 => "00000000",
	8704 => "00000000",
	8705 => "00000000",
	8706 => "00000000",
	8707 => "00000000",
	8708 => "00000000",
	8709 => "00000000",
	8710 => "00000000",
	8711 => "00000000",
	8712 => "00000000",
	8713 => "00000000",
	8714 => "00000000",
	8715 => "00000000",
	8716 => "00000000",
	8717 => "00000000",
	8718 => "00000000",
	8719 => "00000000",
	8720 => "00000000",
	8721 => "00000000",
	8722 => "00000000",
	8723 => "00000000",
	8724 => "00000000",
	8725 => "00000000",
	8726 => "00000000",
	8727 => "00000000",
	8728 => "00000000",
	8729 => "00000000",
	8730 => "00000000",
	8731 => "00000000",
	8732 => "00000000",
	8733 => "00000000",
	8734 => "00000000",
	8735 => "00000000",
	8736 => "00000000",
	8737 => "00000000",
	8738 => "00000000",
	8739 => "00000000",
	8740 => "00000000",
	8741 => "00000000",
	8742 => "00000000",
	8743 => "00000000",
	8744 => "00000000",
	8745 => "00000000",
	8746 => "00000000",
	8747 => "00000000",
	8748 => "00000000",
	8749 => "00000000",
	8750 => "00000000",
	8751 => "11111111",
	8752 => "11111111",
	8753 => "11111111",
	8754 => "11111111",
	8755 => "11111111",
	8756 => "11111111",
	8757 => "11111111",
	8758 => "11111111",
	8759 => "11111111",
	8760 => "11111111",
	8761 => "11111111",
	8762 => "00000000",
	8763 => "00000000",
	8764 => "00000000",
	8765 => "00000000",
	8766 => "00000000",
	8767 => "11111111",
	8768 => "11111111",
	8769 => "11111111",
	8770 => "11111111",
	8771 => "11111111",
	8772 => "11111111",
	8773 => "11111111",
	8774 => "11111111",
	8775 => "11111111",
	8776 => "11111111",
	8777 => "11111111",
	8778 => "00000000",
	8779 => "00000000",
	8780 => "00000000",
	8781 => "00000000",
	8782 => "00000000",
	8783 => "00000000",
	8784 => "00000000",
	8785 => "00000000",
	8786 => "00000000",
	8787 => "00000000",
	8788 => "00000000",
	8789 => "00000000",
	8790 => "00000000",
	8791 => "00000000",
	8792 => "00000000",
	8793 => "00000000",
	8794 => "00000000",
	8795 => "00000000",
	8796 => "00000000",
	8797 => "00000000",
	8798 => "00000000",
	8799 => "00000000",
	8800 => "00000000",
	8801 => "00000000",
	8802 => "00000000",
	8803 => "00000000",
	8804 => "00000000",
	8805 => "00000000",
	8806 => "00000000",
	8807 => "00000000",
	8808 => "00000000",
	8809 => "00000000",
	8810 => "00000000",
	8811 => "00000000",
	8812 => "00000000",
	8813 => "00000000",
	8814 => "00000000",
	8815 => "00000000",
	8816 => "00000000",
	8817 => "00000000",
	8818 => "00000000",
	8819 => "00000000",
	8820 => "00000000",
	8821 => "00000000",
	8822 => "00000000",
	8823 => "00000000",
	8832 => "00000000",
	8833 => "00000000",
	8834 => "00000000",
	8835 => "00000000",
	8836 => "00000000",
	8837 => "00000000",
	8838 => "00000000",
	8839 => "00000000",
	8840 => "00000000",
	8841 => "00000000",
	8842 => "00000000",
	8843 => "00000000",
	8844 => "00000000",
	8845 => "00000000",
	8846 => "00000000",
	8847 => "00000000",
	8848 => "00000000",
	8849 => "00000000",
	8850 => "00000000",
	8851 => "00000000",
	8852 => "00000000",
	8853 => "00000000",
	8854 => "00000000",
	8855 => "00000000",
	8856 => "00000000",
	8857 => "00000000",
	8858 => "00000000",
	8859 => "00000000",
	8860 => "00000000",
	8861 => "00000000",
	8862 => "00000000",
	8863 => "00000000",
	8864 => "00000000",
	8865 => "00000000",
	8866 => "00000000",
	8867 => "00000000",
	8868 => "00000000",
	8869 => "00000000",
	8870 => "00000000",
	8871 => "00000000",
	8872 => "00000000",
	8873 => "00000000",
	8874 => "00000000",
	8875 => "00000000",
	8876 => "00000000",
	8877 => "00000000",
	8878 => "11111111",
	8879 => "11111111",
	8880 => "11111111",
	8881 => "11111111",
	8882 => "11111111",
	8883 => "11111111",
	8884 => "11111111",
	8885 => "11111111",
	8886 => "11111111",
	8887 => "11111111",
	8888 => "11111111",
	8889 => "00000000",
	8890 => "00000000",
	8891 => "00000000",
	8892 => "00000000",
	8893 => "00000000",
	8894 => "00000000",
	8895 => "00000000",
	8896 => "11111111",
	8897 => "11111111",
	8898 => "11111111",
	8899 => "11111111",
	8900 => "11111111",
	8901 => "11111111",
	8902 => "11111111",
	8903 => "11111111",
	8904 => "11111111",
	8905 => "11111111",
	8906 => "11111111",
	8907 => "00000000",
	8908 => "00000000",
	8909 => "00000000",
	8910 => "00000000",
	8911 => "00000000",
	8912 => "00000000",
	8913 => "00000000",
	8914 => "00000000",
	8915 => "00000000",
	8916 => "00000000",
	8917 => "00000000",
	8918 => "00000000",
	8919 => "00000000",
	8920 => "00000000",
	8921 => "00000000",
	8922 => "00000000",
	8923 => "00000000",
	8924 => "00000000",
	8925 => "00000000",
	8926 => "00000000",
	8927 => "00000000",
	8928 => "00000000",
	8929 => "00000000",
	8930 => "00000000",
	8931 => "00000000",
	8932 => "00000000",
	8933 => "00000000",
	8934 => "00000000",
	8935 => "00000000",
	8936 => "00000000",
	8937 => "00000000",
	8938 => "00000000",
	8939 => "00000000",
	8940 => "00000000",
	8941 => "00000000",
	8942 => "00000000",
	8943 => "00000000",
	8944 => "00000000",
	8945 => "00000000",
	8946 => "00000000",
	8947 => "00000000",
	8948 => "00000000",
	8949 => "00000000",
	8950 => "00000000",
	8951 => "00000000",
	8960 => "00000000",
	8961 => "00000000",
	8962 => "00000000",
	8963 => "00000000",
	8964 => "00000000",
	8965 => "00000000",
	8966 => "00000000",
	8967 => "00000000",
	8968 => "00000000",
	8969 => "00000000",
	8970 => "00000000",
	8971 => "00000000",
	8972 => "00000000",
	8973 => "00000000",
	8974 => "00000000",
	8975 => "00000000",
	8976 => "00000000",
	8977 => "00000000",
	8978 => "00000000",
	8979 => "00000000",
	8980 => "00000000",
	8981 => "00000000",
	8982 => "00000000",
	8983 => "00000000",
	8984 => "00000000",
	8985 => "00000000",
	8986 => "00000000",
	8987 => "00000000",
	8988 => "00000000",
	8989 => "00000000",
	8990 => "00000000",
	8991 => "00000000",
	8992 => "00000000",
	8993 => "00000000",
	8994 => "00000000",
	8995 => "00000000",
	8996 => "00000000",
	8997 => "00000000",
	8998 => "00000000",
	8999 => "00000000",
	9000 => "00000000",
	9001 => "00000000",
	9002 => "00000000",
	9003 => "00000000",
	9004 => "00000000",
	9005 => "11111111",
	9006 => "11111111",
	9007 => "11111111",
	9008 => "11111111",
	9009 => "11111111",
	9010 => "11111111",
	9011 => "11111111",
	9012 => "11111111",
	9013 => "11111111",
	9014 => "11111111",
	9015 => "11111111",
	9016 => "00000000",
	9017 => "00000000",
	9018 => "00000000",
	9019 => "00000000",
	9020 => "00000000",
	9021 => "00000000",
	9022 => "00000000",
	9023 => "00000000",
	9024 => "00000000",
	9025 => "11111111",
	9026 => "11111111",
	9027 => "11111111",
	9028 => "11111111",
	9029 => "11111111",
	9030 => "11111111",
	9031 => "11111111",
	9032 => "11111111",
	9033 => "11111111",
	9034 => "11111111",
	9035 => "11111111",
	9036 => "00000000",
	9037 => "00000000",
	9038 => "00000000",
	9039 => "00000000",
	9040 => "00000000",
	9041 => "00000000",
	9042 => "00000000",
	9043 => "00000000",
	9044 => "00000000",
	9045 => "00000000",
	9046 => "00000000",
	9047 => "00000000",
	9048 => "00000000",
	9049 => "00000000",
	9050 => "00000000",
	9051 => "00000000",
	9052 => "00000000",
	9053 => "00000000",
	9054 => "00000000",
	9055 => "00000000",
	9056 => "00000000",
	9057 => "00000000",
	9058 => "00000000",
	9059 => "00000000",
	9060 => "00000000",
	9061 => "00000000",
	9062 => "00000000",
	9063 => "00000000",
	9064 => "00000000",
	9065 => "00000000",
	9066 => "00000000",
	9067 => "00000000",
	9068 => "00000000",
	9069 => "00000000",
	9070 => "00000000",
	9071 => "00000000",
	9072 => "00000000",
	9073 => "00000000",
	9074 => "00000000",
	9075 => "00000000",
	9076 => "00000000",
	9077 => "00000000",
	9078 => "00000000",
	9079 => "00000000",
	9088 => "00000000",
	9089 => "00000000",
	9090 => "00000000",
	9091 => "00000000",
	9092 => "00000000",
	9093 => "00000000",
	9094 => "00000000",
	9095 => "00000000",
	9096 => "00000000",
	9097 => "00000000",
	9098 => "00000000",
	9099 => "00000000",
	9100 => "00000000",
	9101 => "00000000",
	9102 => "00000000",
	9103 => "00000000",
	9104 => "00000000",
	9105 => "00000000",
	9106 => "00000000",
	9107 => "00000000",
	9108 => "00000000",
	9109 => "00000000",
	9110 => "00000000",
	9111 => "00000000",
	9112 => "00000000",
	9113 => "00000000",
	9114 => "00000000",
	9115 => "00000000",
	9116 => "00000000",
	9117 => "00000000",
	9118 => "00000000",
	9119 => "00000000",
	9120 => "00000000",
	9121 => "00000000",
	9122 => "00000000",
	9123 => "00000000",
	9124 => "00000000",
	9125 => "00000000",
	9126 => "00000000",
	9127 => "00000000",
	9128 => "00000000",
	9129 => "00000000",
	9130 => "00000000",
	9131 => "00000000",
	9132 => "11111111",
	9133 => "11111111",
	9134 => "11111111",
	9135 => "11111111",
	9136 => "11111111",
	9137 => "11111111",
	9138 => "11111111",
	9139 => "11111111",
	9140 => "11111111",
	9141 => "11111111",
	9142 => "11111111",
	9143 => "00000000",
	9144 => "00000000",
	9145 => "00000000",
	9146 => "00000000",
	9147 => "00000000",
	9148 => "00000000",
	9149 => "00000000",
	9150 => "00000000",
	9151 => "00000000",
	9152 => "00000000",
	9153 => "00000000",
	9154 => "11111111",
	9155 => "11111111",
	9156 => "11111111",
	9157 => "11111111",
	9158 => "11111111",
	9159 => "11111111",
	9160 => "11111111",
	9161 => "11111111",
	9162 => "11111111",
	9163 => "11111111",
	9164 => "11111111",
	9165 => "00000000",
	9166 => "00000000",
	9167 => "00000000",
	9168 => "00000000",
	9169 => "00000000",
	9170 => "00000000",
	9171 => "00000000",
	9172 => "00000000",
	9173 => "00000000",
	9174 => "00000000",
	9175 => "00000000",
	9176 => "00000000",
	9177 => "00000000",
	9178 => "00000000",
	9179 => "00000000",
	9180 => "00000000",
	9181 => "00000000",
	9182 => "00000000",
	9183 => "00000000",
	9184 => "00000000",
	9185 => "00000000",
	9186 => "00000000",
	9187 => "00000000",
	9188 => "00000000",
	9189 => "00000000",
	9190 => "00000000",
	9191 => "00000000",
	9192 => "00000000",
	9193 => "00000000",
	9194 => "00000000",
	9195 => "00000000",
	9196 => "00000000",
	9197 => "00000000",
	9198 => "00000000",
	9199 => "00000000",
	9200 => "00000000",
	9201 => "00000000",
	9202 => "00000000",
	9203 => "00000000",
	9204 => "00000000",
	9205 => "00000000",
	9206 => "00000000",
	9207 => "00000000",
	9216 => "00000000",
	9217 => "00000000",
	9218 => "00000000",
	9219 => "00000000",
	9220 => "00000000",
	9221 => "00000000",
	9222 => "00000000",
	9223 => "00000000",
	9224 => "00000000",
	9225 => "00000000",
	9226 => "00000000",
	9227 => "00000000",
	9228 => "00000000",
	9229 => "00000000",
	9230 => "00000000",
	9231 => "00000000",
	9232 => "00000000",
	9233 => "00000000",
	9234 => "00000000",
	9235 => "00000000",
	9236 => "00000000",
	9237 => "00000000",
	9238 => "00000000",
	9239 => "00000000",
	9240 => "00000000",
	9241 => "00000000",
	9242 => "00000000",
	9243 => "00000000",
	9244 => "00000000",
	9245 => "00000000",
	9246 => "00000000",
	9247 => "00000000",
	9248 => "00000000",
	9249 => "00000000",
	9250 => "00000000",
	9251 => "00000000",
	9252 => "00000000",
	9253 => "00000000",
	9254 => "00000000",
	9255 => "00000000",
	9256 => "00000000",
	9257 => "00000000",
	9258 => "00000000",
	9259 => "11111111",
	9260 => "11111111",
	9261 => "11111111",
	9262 => "11111111",
	9263 => "11111111",
	9264 => "11111111",
	9265 => "11111111",
	9266 => "11111111",
	9267 => "11111111",
	9268 => "11111111",
	9269 => "11111111",
	9270 => "00000000",
	9271 => "00000000",
	9272 => "00000000",
	9273 => "00000000",
	9274 => "00000000",
	9275 => "00000000",
	9276 => "00000000",
	9277 => "00000000",
	9278 => "00000000",
	9279 => "00000000",
	9280 => "00000000",
	9281 => "00000000",
	9282 => "00000000",
	9283 => "11111111",
	9284 => "11111111",
	9285 => "11111111",
	9286 => "11111111",
	9287 => "11111111",
	9288 => "11111111",
	9289 => "11111111",
	9290 => "11111111",
	9291 => "11111111",
	9292 => "11111111",
	9293 => "11111111",
	9294 => "00000000",
	9295 => "00000000",
	9296 => "00000000",
	9297 => "00000000",
	9298 => "00000000",
	9299 => "00000000",
	9300 => "00000000",
	9301 => "00000000",
	9302 => "00000000",
	9303 => "00000000",
	9304 => "00000000",
	9305 => "00000000",
	9306 => "00000000",
	9307 => "00000000",
	9308 => "00000000",
	9309 => "00000000",
	9310 => "00000000",
	9311 => "00000000",
	9312 => "00000000",
	9313 => "00000000",
	9314 => "00000000",
	9315 => "00000000",
	9316 => "00000000",
	9317 => "00000000",
	9318 => "00000000",
	9319 => "00000000",
	9320 => "00000000",
	9321 => "00000000",
	9322 => "00000000",
	9323 => "00000000",
	9324 => "00000000",
	9325 => "00000000",
	9326 => "00000000",
	9327 => "00000000",
	9328 => "00000000",
	9329 => "00000000",
	9330 => "00000000",
	9331 => "00000000",
	9332 => "00000000",
	9333 => "00000000",
	9334 => "00000000",
	9335 => "00000000",
	9344 => "00000000",
	9345 => "00000000",
	9346 => "00000000",
	9347 => "00000000",
	9348 => "00000000",
	9349 => "00000000",
	9350 => "00000000",
	9351 => "00000000",
	9352 => "00000000",
	9353 => "00000000",
	9354 => "00000000",
	9355 => "00000000",
	9356 => "00000000",
	9357 => "00000000",
	9358 => "00000000",
	9359 => "00000000",
	9360 => "00000000",
	9361 => "00000000",
	9362 => "00000000",
	9363 => "00000000",
	9364 => "00000000",
	9365 => "00000000",
	9366 => "00000000",
	9367 => "00000000",
	9368 => "00000000",
	9369 => "00000000",
	9370 => "00000000",
	9371 => "00000000",
	9372 => "00000000",
	9373 => "00000000",
	9374 => "00000000",
	9375 => "00000000",
	9376 => "00000000",
	9377 => "00000000",
	9378 => "00000000",
	9379 => "00000000",
	9380 => "00000000",
	9381 => "00000000",
	9382 => "00000000",
	9383 => "00000000",
	9384 => "00000000",
	9385 => "00000000",
	9386 => "11111111",
	9387 => "11111111",
	9388 => "11111111",
	9389 => "11111111",
	9390 => "11111111",
	9391 => "11111111",
	9392 => "11111111",
	9393 => "11111111",
	9394 => "11111111",
	9395 => "11111111",
	9396 => "11111111",
	9397 => "00000000",
	9398 => "00000000",
	9399 => "00000000",
	9400 => "00000000",
	9401 => "00000000",
	9402 => "00000000",
	9403 => "00000000",
	9404 => "00000000",
	9405 => "00000000",
	9406 => "00000000",
	9407 => "00000000",
	9408 => "00000000",
	9409 => "00000000",
	9410 => "00000000",
	9411 => "00000000",
	9412 => "11111111",
	9413 => "11111111",
	9414 => "11111111",
	9415 => "11111111",
	9416 => "11111111",
	9417 => "11111111",
	9418 => "11111111",
	9419 => "11111111",
	9420 => "11111111",
	9421 => "11111111",
	9422 => "11111111",
	9423 => "00000000",
	9424 => "00000000",
	9425 => "00000000",
	9426 => "00000000",
	9427 => "00000000",
	9428 => "00000000",
	9429 => "00000000",
	9430 => "00000000",
	9431 => "00000000",
	9432 => "00000000",
	9433 => "00000000",
	9434 => "00000000",
	9435 => "00000000",
	9436 => "00000000",
	9437 => "00000000",
	9438 => "00000000",
	9439 => "00000000",
	9440 => "00000000",
	9441 => "00000000",
	9442 => "00000000",
	9443 => "00000000",
	9444 => "00000000",
	9445 => "00000000",
	9446 => "00000000",
	9447 => "00000000",
	9448 => "00000000",
	9449 => "00000000",
	9450 => "00000000",
	9451 => "00000000",
	9452 => "00000000",
	9453 => "00000000",
	9454 => "00000000",
	9455 => "00000000",
	9456 => "00000000",
	9457 => "00000000",
	9458 => "00000000",
	9459 => "00000000",
	9460 => "00000000",
	9461 => "00000000",
	9462 => "00000000",
	9463 => "00000000",
	9472 => "00000000",
	9473 => "00000000",
	9474 => "00000000",
	9475 => "00000000",
	9476 => "00000000",
	9477 => "00000000",
	9478 => "00000000",
	9479 => "00000000",
	9480 => "00000000",
	9481 => "00000000",
	9482 => "00000000",
	9483 => "00000000",
	9484 => "00000000",
	9485 => "00000000",
	9486 => "00000000",
	9487 => "00000000",
	9488 => "00000000",
	9489 => "00000000",
	9490 => "00000000",
	9491 => "00000000",
	9492 => "00000000",
	9493 => "00000000",
	9494 => "00000000",
	9495 => "00000000",
	9496 => "00000000",
	9497 => "00000000",
	9498 => "00000000",
	9499 => "00000000",
	9500 => "00000000",
	9501 => "00000000",
	9502 => "00000000",
	9503 => "00000000",
	9504 => "00000000",
	9505 => "00000000",
	9506 => "00000000",
	9507 => "00000000",
	9508 => "00000000",
	9509 => "00000000",
	9510 => "00000000",
	9511 => "00000000",
	9512 => "00000000",
	9513 => "11111111",
	9514 => "11111111",
	9515 => "11111111",
	9516 => "11111111",
	9517 => "11111111",
	9518 => "11111111",
	9519 => "11111111",
	9520 => "11111111",
	9521 => "11111111",
	9522 => "11111111",
	9523 => "11111111",
	9524 => "00000000",
	9525 => "00000000",
	9526 => "00000000",
	9527 => "00000000",
	9528 => "00000000",
	9529 => "00000000",
	9530 => "00000000",
	9531 => "00000000",
	9532 => "00000000",
	9533 => "00000000",
	9534 => "00000000",
	9535 => "00000000",
	9536 => "00000000",
	9537 => "00000000",
	9538 => "00000000",
	9539 => "00000000",
	9540 => "00000000",
	9541 => "11111111",
	9542 => "11111111",
	9543 => "11111111",
	9544 => "11111111",
	9545 => "11111111",
	9546 => "11111111",
	9547 => "11111111",
	9548 => "11111111",
	9549 => "11111111",
	9550 => "11111111",
	9551 => "11111111",
	9552 => "00000000",
	9553 => "00000000",
	9554 => "00000000",
	9555 => "00000000",
	9556 => "00000000",
	9557 => "00000000",
	9558 => "00000000",
	9559 => "00000000",
	9560 => "00000000",
	9561 => "00000000",
	9562 => "00000000",
	9563 => "00000000",
	9564 => "00000000",
	9565 => "00000000",
	9566 => "00000000",
	9567 => "00000000",
	9568 => "00000000",
	9569 => "00000000",
	9570 => "00000000",
	9571 => "00000000",
	9572 => "00000000",
	9573 => "00000000",
	9574 => "00000000",
	9575 => "00000000",
	9576 => "00000000",
	9577 => "00000000",
	9578 => "00000000",
	9579 => "00000000",
	9580 => "00000000",
	9581 => "00000000",
	9582 => "00000000",
	9583 => "00000000",
	9584 => "00000000",
	9585 => "00000000",
	9586 => "00000000",
	9587 => "00000000",
	9588 => "00000000",
	9589 => "00000000",
	9590 => "00000000",
	9591 => "00000000",
	9600 => "00000000",
	9601 => "00000000",
	9602 => "00000000",
	9603 => "00000000",
	9604 => "00000000",
	9605 => "00000000",
	9606 => "00000000",
	9607 => "00000000",
	9608 => "00000000",
	9609 => "00000000",
	9610 => "00000000",
	9611 => "00000000",
	9612 => "00000000",
	9613 => "00000000",
	9614 => "00000000",
	9615 => "00000000",
	9616 => "00000000",
	9617 => "00000000",
	9618 => "00000000",
	9619 => "00000000",
	9620 => "00000000",
	9621 => "00000000",
	9622 => "00000000",
	9623 => "00000000",
	9624 => "00000000",
	9625 => "00000000",
	9626 => "00000000",
	9627 => "00000000",
	9628 => "00000000",
	9629 => "00000000",
	9630 => "00000000",
	9631 => "00000000",
	9632 => "00000000",
	9633 => "00000000",
	9634 => "00000000",
	9635 => "00000000",
	9636 => "00000000",
	9637 => "00000000",
	9638 => "00000000",
	9639 => "00000000",
	9640 => "11111111",
	9641 => "11111111",
	9642 => "11111111",
	9643 => "11111111",
	9644 => "11111111",
	9645 => "11111111",
	9646 => "11111111",
	9647 => "11111111",
	9648 => "11111111",
	9649 => "11111111",
	9650 => "11111111",
	9651 => "00000000",
	9652 => "00000000",
	9653 => "00000000",
	9654 => "00000000",
	9655 => "00000000",
	9656 => "00000000",
	9657 => "00000000",
	9658 => "00000000",
	9659 => "00000000",
	9660 => "00000000",
	9661 => "00000000",
	9662 => "00000000",
	9663 => "00000000",
	9664 => "00000000",
	9665 => "00000000",
	9666 => "00000000",
	9667 => "00000000",
	9668 => "00000000",
	9669 => "00000000",
	9670 => "11111111",
	9671 => "11111111",
	9672 => "11111111",
	9673 => "11111111",
	9674 => "11111111",
	9675 => "11111111",
	9676 => "11111111",
	9677 => "11111111",
	9678 => "11111111",
	9679 => "11111111",
	9680 => "11111111",
	9681 => "00000000",
	9682 => "00000000",
	9683 => "00000000",
	9684 => "00000000",
	9685 => "00000000",
	9686 => "00000000",
	9687 => "00000000",
	9688 => "00000000",
	9689 => "00000000",
	9690 => "00000000",
	9691 => "00000000",
	9692 => "00000000",
	9693 => "00000000",
	9694 => "00000000",
	9695 => "00000000",
	9696 => "00000000",
	9697 => "00000000",
	9698 => "00000000",
	9699 => "00000000",
	9700 => "00000000",
	9701 => "00000000",
	9702 => "00000000",
	9703 => "00000000",
	9704 => "00000000",
	9705 => "00000000",
	9706 => "00000000",
	9707 => "00000000",
	9708 => "00000000",
	9709 => "00000000",
	9710 => "00000000",
	9711 => "00000000",
	9712 => "00000000",
	9713 => "00000000",
	9714 => "00000000",
	9715 => "00000000",
	9716 => "00000000",
	9717 => "00000000",
	9718 => "00000000",
	9719 => "00000000",
	9728 => "00000000",
	9729 => "00000000",
	9730 => "00000000",
	9731 => "00000000",
	9732 => "00000000",
	9733 => "00000000",
	9734 => "00000000",
	9735 => "00000000",
	9736 => "00000000",
	9737 => "00000000",
	9738 => "00000000",
	9739 => "00000000",
	9740 => "00000000",
	9741 => "00000000",
	9742 => "00000000",
	9743 => "00000000",
	9744 => "00000000",
	9745 => "00000000",
	9746 => "00000000",
	9747 => "00000000",
	9748 => "00000000",
	9749 => "00000000",
	9750 => "00000000",
	9751 => "00000000",
	9752 => "00000000",
	9753 => "00000000",
	9754 => "00000000",
	9755 => "00000000",
	9756 => "00000000",
	9757 => "00000000",
	9758 => "00000000",
	9759 => "00000000",
	9760 => "00000000",
	9761 => "00000000",
	9762 => "00000000",
	9763 => "00000000",
	9764 => "00000000",
	9765 => "00000000",
	9766 => "00000000",
	9767 => "11111111",
	9768 => "11111111",
	9769 => "11111111",
	9770 => "11111111",
	9771 => "11111111",
	9772 => "11111111",
	9773 => "11111111",
	9774 => "11111111",
	9775 => "11111111",
	9776 => "11111111",
	9777 => "11111111",
	9778 => "00000000",
	9779 => "00000000",
	9780 => "00000000",
	9781 => "00000000",
	9782 => "00000000",
	9783 => "00000000",
	9784 => "00000000",
	9785 => "00000000",
	9786 => "00000000",
	9787 => "00000000",
	9788 => "00000000",
	9789 => "00000000",
	9790 => "00000000",
	9791 => "00000000",
	9792 => "00000000",
	9793 => "00000000",
	9794 => "00000000",
	9795 => "00000000",
	9796 => "00000000",
	9797 => "00000000",
	9798 => "00000000",
	9799 => "11111111",
	9800 => "11111111",
	9801 => "11111111",
	9802 => "11111111",
	9803 => "11111111",
	9804 => "11111111",
	9805 => "11111111",
	9806 => "11111111",
	9807 => "11111111",
	9808 => "11111111",
	9809 => "11111111",
	9810 => "00000000",
	9811 => "00000000",
	9812 => "00000000",
	9813 => "00000000",
	9814 => "00000000",
	9815 => "00000000",
	9816 => "00000000",
	9817 => "00000000",
	9818 => "00000000",
	9819 => "00000000",
	9820 => "00000000",
	9821 => "00000000",
	9822 => "00000000",
	9823 => "00000000",
	9824 => "00000000",
	9825 => "00000000",
	9826 => "00000000",
	9827 => "00000000",
	9828 => "00000000",
	9829 => "00000000",
	9830 => "00000000",
	9831 => "00000000",
	9832 => "00000000",
	9833 => "00000000",
	9834 => "00000000",
	9835 => "00000000",
	9836 => "00000000",
	9837 => "00000000",
	9838 => "00000000",
	9839 => "00000000",
	9840 => "00000000",
	9841 => "00000000",
	9842 => "00000000",
	9843 => "00000000",
	9844 => "00000000",
	9845 => "00000000",
	9846 => "00000000",
	9847 => "00000000",
	9856 => "00000000",
	9857 => "00000000",
	9858 => "00000000",
	9859 => "00000000",
	9860 => "00000000",
	9861 => "00000000",
	9862 => "00000000",
	9863 => "00000000",
	9864 => "00000000",
	9865 => "00000000",
	9866 => "00000000",
	9867 => "00000000",
	9868 => "00000000",
	9869 => "00000000",
	9870 => "00000000",
	9871 => "00000000",
	9872 => "00000000",
	9873 => "00000000",
	9874 => "00000000",
	9875 => "00000000",
	9876 => "00000000",
	9877 => "00000000",
	9878 => "00000000",
	9879 => "00000000",
	9880 => "00000000",
	9881 => "00000000",
	9882 => "00000000",
	9883 => "00000000",
	9884 => "00000000",
	9885 => "00000000",
	9886 => "00000000",
	9887 => "00000000",
	9888 => "00000000",
	9889 => "00000000",
	9890 => "00000000",
	9891 => "00000000",
	9892 => "00000000",
	9893 => "00000000",
	9894 => "11111111",
	9895 => "11111111",
	9896 => "11111111",
	9897 => "11111111",
	9898 => "11111111",
	9899 => "11111111",
	9900 => "11111111",
	9901 => "11111111",
	9902 => "11111111",
	9903 => "11111111",
	9904 => "11111111",
	9905 => "00000000",
	9906 => "00000000",
	9907 => "00000000",
	9908 => "00000000",
	9909 => "00000000",
	9910 => "00000000",
	9911 => "00000000",
	9912 => "00000000",
	9913 => "00000000",
	9914 => "00000000",
	9915 => "00000000",
	9916 => "00000000",
	9917 => "00000000",
	9918 => "00000000",
	9919 => "00000000",
	9920 => "00000000",
	9921 => "00000000",
	9922 => "00000000",
	9923 => "00000000",
	9924 => "00000000",
	9925 => "00000000",
	9926 => "00000000",
	9927 => "00000000",
	9928 => "11111111",
	9929 => "11111111",
	9930 => "11111111",
	9931 => "11111111",
	9932 => "11111111",
	9933 => "11111111",
	9934 => "11111111",
	9935 => "11111111",
	9936 => "11111111",
	9937 => "11111111",
	9938 => "11111111",
	9939 => "00000000",
	9940 => "00000000",
	9941 => "00000000",
	9942 => "00000000",
	9943 => "00000000",
	9944 => "00000000",
	9945 => "00000000",
	9946 => "00000000",
	9947 => "00000000",
	9948 => "00000000",
	9949 => "00000000",
	9950 => "00000000",
	9951 => "00000000",
	9952 => "00000000",
	9953 => "00000000",
	9954 => "00000000",
	9955 => "00000000",
	9956 => "00000000",
	9957 => "00000000",
	9958 => "00000000",
	9959 => "00000000",
	9960 => "00000000",
	9961 => "00000000",
	9962 => "00000000",
	9963 => "00000000",
	9964 => "00000000",
	9965 => "00000000",
	9966 => "00000000",
	9967 => "00000000",
	9968 => "00000000",
	9969 => "00000000",
	9970 => "00000000",
	9971 => "00000000",
	9972 => "00000000",
	9973 => "00000000",
	9974 => "00000000",
	9975 => "00000000",
	9984 => "00000000",
	9985 => "00000000",
	9986 => "00000000",
	9987 => "00000000",
	9988 => "00000000",
	9989 => "00000000",
	9990 => "00000000",
	9991 => "00000000",
	9992 => "00000000",
	9993 => "00000000",
	9994 => "00000000",
	9995 => "00000000",
	9996 => "00000000",
	9997 => "00000000",
	9998 => "00000000",
	9999 => "00000000",
	10000 => "00000000",
	10001 => "00000000",
	10002 => "00000000",
	10003 => "00000000",
	10004 => "00000000",
	10005 => "00000000",
	10006 => "00000000",
	10007 => "00000000",
	10008 => "00000000",
	10009 => "00000000",
	10010 => "00000000",
	10011 => "00000000",
	10012 => "00000000",
	10013 => "00000000",
	10014 => "00000000",
	10015 => "00000000",
	10016 => "00000000",
	10017 => "00000000",
	10018 => "00000000",
	10019 => "00000000",
	10020 => "00000000",
	10021 => "11111111",
	10022 => "11111111",
	10023 => "11111111",
	10024 => "11111111",
	10025 => "11111111",
	10026 => "11111111",
	10027 => "11111111",
	10028 => "11111111",
	10029 => "11111111",
	10030 => "11111111",
	10031 => "11111111",
	10032 => "00000000",
	10033 => "00000000",
	10034 => "00000000",
	10035 => "00000000",
	10036 => "00000000",
	10037 => "00000000",
	10038 => "00000000",
	10039 => "00000000",
	10040 => "00000000",
	10041 => "00000000",
	10042 => "00000000",
	10043 => "00000000",
	10044 => "00000000",
	10045 => "00000000",
	10046 => "00000000",
	10047 => "00000000",
	10048 => "00000000",
	10049 => "00000000",
	10050 => "00000000",
	10051 => "00000000",
	10052 => "00000000",
	10053 => "00000000",
	10054 => "00000000",
	10055 => "00000000",
	10056 => "00000000",
	10057 => "11111111",
	10058 => "11111111",
	10059 => "11111111",
	10060 => "11111111",
	10061 => "11111111",
	10062 => "11111111",
	10063 => "11111111",
	10064 => "11111111",
	10065 => "11111111",
	10066 => "11111111",
	10067 => "11111111",
	10068 => "00000000",
	10069 => "00000000",
	10070 => "00000000",
	10071 => "00000000",
	10072 => "00000000",
	10073 => "00000000",
	10074 => "00000000",
	10075 => "00000000",
	10076 => "00000000",
	10077 => "00000000",
	10078 => "00000000",
	10079 => "00000000",
	10080 => "00000000",
	10081 => "00000000",
	10082 => "00000000",
	10083 => "00000000",
	10084 => "00000000",
	10085 => "00000000",
	10086 => "00000000",
	10087 => "00000000",
	10088 => "00000000",
	10089 => "00000000",
	10090 => "00000000",
	10091 => "00000000",
	10092 => "00000000",
	10093 => "00000000",
	10094 => "00000000",
	10095 => "00000000",
	10096 => "00000000",
	10097 => "00000000",
	10098 => "00000000",
	10099 => "00000000",
	10100 => "00000000",
	10101 => "00000000",
	10102 => "00000000",
	10103 => "00000000",
	10112 => "00000000",
	10113 => "00000000",
	10114 => "00000000",
	10115 => "00000000",
	10116 => "00000000",
	10117 => "00000000",
	10118 => "00000000",
	10119 => "00000000",
	10120 => "00000000",
	10121 => "00000000",
	10122 => "00000000",
	10123 => "00000000",
	10124 => "00000000",
	10125 => "00000000",
	10126 => "00000000",
	10127 => "00000000",
	10128 => "00000000",
	10129 => "00000000",
	10130 => "00000000",
	10131 => "00000000",
	10132 => "00000000",
	10133 => "00000000",
	10134 => "00000000",
	10135 => "00000000",
	10136 => "00000000",
	10137 => "00000000",
	10138 => "00000000",
	10139 => "00000000",
	10140 => "00000000",
	10141 => "00000000",
	10142 => "00000000",
	10143 => "00000000",
	10144 => "00000000",
	10145 => "00000000",
	10146 => "00000000",
	10147 => "00000000",
	10148 => "11111111",
	10149 => "11111111",
	10150 => "11111111",
	10151 => "11111111",
	10152 => "11111111",
	10153 => "11111111",
	10154 => "11111111",
	10155 => "11111111",
	10156 => "11111111",
	10157 => "11111111",
	10158 => "11111111",
	10159 => "00000000",
	10160 => "00000000",
	10161 => "00000000",
	10162 => "00000000",
	10163 => "00000000",
	10164 => "00000000",
	10165 => "00000000",
	10166 => "00000000",
	10167 => "00000000",
	10168 => "00000000",
	10169 => "00000000",
	10170 => "00000000",
	10171 => "00000000",
	10172 => "00000000",
	10173 => "00000000",
	10174 => "00000000",
	10175 => "00000000",
	10176 => "00000000",
	10177 => "00000000",
	10178 => "00000000",
	10179 => "00000000",
	10180 => "00000000",
	10181 => "00000000",
	10182 => "00000000",
	10183 => "00000000",
	10184 => "00000000",
	10185 => "00000000",
	10186 => "11111111",
	10187 => "11111111",
	10188 => "11111111",
	10189 => "11111111",
	10190 => "11111111",
	10191 => "11111111",
	10192 => "11111111",
	10193 => "11111111",
	10194 => "11111111",
	10195 => "11111111",
	10196 => "11111111",
	10197 => "00000000",
	10198 => "00000000",
	10199 => "00000000",
	10200 => "00000000",
	10201 => "00000000",
	10202 => "00000000",
	10203 => "00000000",
	10204 => "00000000",
	10205 => "00000000",
	10206 => "00000000",
	10207 => "00000000",
	10208 => "00000000",
	10209 => "00000000",
	10210 => "00000000",
	10211 => "00000000",
	10212 => "00000000",
	10213 => "00000000",
	10214 => "00000000",
	10215 => "00000000",
	10216 => "00000000",
	10217 => "00000000",
	10218 => "00000000",
	10219 => "00000000",
	10220 => "00000000",
	10221 => "00000000",
	10222 => "00000000",
	10223 => "00000000",
	10224 => "00000000",
	10225 => "00000000",
	10226 => "00000000",
	10227 => "00000000",
	10228 => "00000000",
	10229 => "00000000",
	10230 => "00000000",
	10231 => "00000000",
	10240 => "00000000",
	10241 => "00000000",
	10242 => "00000000",
	10243 => "00000000",
	10244 => "00000000",
	10245 => "00000000",
	10246 => "00000000",
	10247 => "00000000",
	10248 => "00000000",
	10249 => "00000000",
	10250 => "00000000",
	10251 => "00000000",
	10252 => "00000000",
	10253 => "00000000",
	10254 => "00000000",
	10255 => "00000000",
	10256 => "00000000",
	10257 => "00000000",
	10258 => "00000000",
	10259 => "00000000",
	10260 => "00000000",
	10261 => "00000000",
	10262 => "00000000",
	10263 => "00000000",
	10264 => "00000000",
	10265 => "00000000",
	10266 => "00000000",
	10267 => "00000000",
	10268 => "00000000",
	10269 => "00000000",
	10270 => "00000000",
	10271 => "00000000",
	10272 => "00000000",
	10273 => "00000000",
	10274 => "00000000",
	10275 => "11111111",
	10276 => "11111111",
	10277 => "11111111",
	10278 => "11111111",
	10279 => "11111111",
	10280 => "11111111",
	10281 => "11111111",
	10282 => "11111111",
	10283 => "11111111",
	10284 => "11111111",
	10285 => "11111111",
	10286 => "00000000",
	10287 => "00000000",
	10288 => "00000000",
	10289 => "00000000",
	10290 => "00000000",
	10291 => "00000000",
	10292 => "00000000",
	10293 => "00000000",
	10294 => "00000000",
	10295 => "00000000",
	10296 => "00000000",
	10297 => "00000000",
	10298 => "00000000",
	10299 => "00000000",
	10300 => "00000000",
	10301 => "00000000",
	10302 => "00000000",
	10303 => "00000000",
	10304 => "00000000",
	10305 => "00000000",
	10306 => "00000000",
	10307 => "00000000",
	10308 => "00000000",
	10309 => "00000000",
	10310 => "00000000",
	10311 => "00000000",
	10312 => "00000000",
	10313 => "00000000",
	10314 => "00000000",
	10315 => "11111111",
	10316 => "11111111",
	10317 => "11111111",
	10318 => "11111111",
	10319 => "11111111",
	10320 => "11111111",
	10321 => "11111111",
	10322 => "11111111",
	10323 => "11111111",
	10324 => "11111111",
	10325 => "11111111",
	10326 => "00000000",
	10327 => "00000000",
	10328 => "00000000",
	10329 => "00000000",
	10330 => "00000000",
	10331 => "00000000",
	10332 => "00000000",
	10333 => "00000000",
	10334 => "00000000",
	10335 => "00000000",
	10336 => "00000000",
	10337 => "00000000",
	10338 => "00000000",
	10339 => "00000000",
	10340 => "00000000",
	10341 => "00000000",
	10342 => "00000000",
	10343 => "00000000",
	10344 => "00000000",
	10345 => "00000000",
	10346 => "00000000",
	10347 => "00000000",
	10348 => "00000000",
	10349 => "00000000",
	10350 => "00000000",
	10351 => "00000000",
	10352 => "00000000",
	10353 => "00000000",
	10354 => "00000000",
	10355 => "00000000",
	10356 => "00000000",
	10357 => "00000000",
	10358 => "00000000",
	10359 => "00000000",
	10368 => "00000000",
	10369 => "00000000",
	10370 => "00000000",
	10371 => "00000000",
	10372 => "00000000",
	10373 => "00000000",
	10374 => "00000000",
	10375 => "00000000",
	10376 => "00000000",
	10377 => "00000000",
	10378 => "00000000",
	10379 => "00000000",
	10380 => "00000000",
	10381 => "00000000",
	10382 => "00000000",
	10383 => "00000000",
	10384 => "00000000",
	10385 => "00000000",
	10386 => "00000000",
	10387 => "00000000",
	10388 => "00000000",
	10389 => "00000000",
	10390 => "00000000",
	10391 => "00000000",
	10392 => "00000000",
	10393 => "00000000",
	10394 => "00000000",
	10395 => "00000000",
	10396 => "00000000",
	10397 => "00000000",
	10398 => "00000000",
	10399 => "00000000",
	10400 => "00000000",
	10401 => "00000000",
	10402 => "11111111",
	10403 => "11111111",
	10404 => "11111111",
	10405 => "11111111",
	10406 => "11111111",
	10407 => "11111111",
	10408 => "11111111",
	10409 => "11111111",
	10410 => "11111111",
	10411 => "11111111",
	10412 => "11111111",
	10413 => "00000000",
	10414 => "00000000",
	10415 => "00000000",
	10416 => "00000000",
	10417 => "00000000",
	10418 => "00000000",
	10419 => "00000000",
	10420 => "00000000",
	10421 => "00000000",
	10422 => "00000000",
	10423 => "00000000",
	10424 => "00000000",
	10425 => "00000000",
	10426 => "00000000",
	10427 => "00000000",
	10428 => "00000000",
	10429 => "00000000",
	10430 => "00000000",
	10431 => "00000000",
	10432 => "00000000",
	10433 => "00000000",
	10434 => "00000000",
	10435 => "00000000",
	10436 => "00000000",
	10437 => "00000000",
	10438 => "00000000",
	10439 => "00000000",
	10440 => "00000000",
	10441 => "00000000",
	10442 => "00000000",
	10443 => "00000000",
	10444 => "11111111",
	10445 => "11111111",
	10446 => "11111111",
	10447 => "11111111",
	10448 => "11111111",
	10449 => "11111111",
	10450 => "11111111",
	10451 => "11111111",
	10452 => "11111111",
	10453 => "11111111",
	10454 => "11111111",
	10455 => "00000000",
	10456 => "00000000",
	10457 => "00000000",
	10458 => "00000000",
	10459 => "00000000",
	10460 => "00000000",
	10461 => "00000000",
	10462 => "00000000",
	10463 => "00000000",
	10464 => "00000000",
	10465 => "00000000",
	10466 => "00000000",
	10467 => "00000000",
	10468 => "00000000",
	10469 => "00000000",
	10470 => "00000000",
	10471 => "00000000",
	10472 => "00000000",
	10473 => "00000000",
	10474 => "00000000",
	10475 => "00000000",
	10476 => "00000000",
	10477 => "00000000",
	10478 => "00000000",
	10479 => "00000000",
	10480 => "00000000",
	10481 => "00000000",
	10482 => "00000000",
	10483 => "00000000",
	10484 => "00000000",
	10485 => "00000000",
	10486 => "00000000",
	10487 => "00000000",
	10496 => "00000000",
	10497 => "00000000",
	10498 => "00000000",
	10499 => "00000000",
	10500 => "00000000",
	10501 => "00000000",
	10502 => "00000000",
	10503 => "00000000",
	10504 => "00000000",
	10505 => "00000000",
	10506 => "00000000",
	10507 => "00000000",
	10508 => "00000000",
	10509 => "00000000",
	10510 => "00000000",
	10511 => "00000000",
	10512 => "00000000",
	10513 => "00000000",
	10514 => "00000000",
	10515 => "00000000",
	10516 => "00000000",
	10517 => "00000000",
	10518 => "00000000",
	10519 => "00000000",
	10520 => "00000000",
	10521 => "00000000",
	10522 => "00000000",
	10523 => "00000000",
	10524 => "00000000",
	10525 => "00000000",
	10526 => "00000000",
	10527 => "00000000",
	10528 => "00000000",
	10529 => "11111111",
	10530 => "11111111",
	10531 => "11111111",
	10532 => "11111111",
	10533 => "11111111",
	10534 => "11111111",
	10535 => "11111111",
	10536 => "11111111",
	10537 => "11111111",
	10538 => "11111111",
	10539 => "11111111",
	10540 => "00000000",
	10541 => "00000000",
	10542 => "00000000",
	10543 => "00000000",
	10544 => "00000000",
	10545 => "00000000",
	10546 => "00000000",
	10547 => "00000000",
	10548 => "00000000",
	10549 => "00000000",
	10550 => "00000000",
	10551 => "00000000",
	10552 => "00000000",
	10553 => "00000000",
	10554 => "00000000",
	10555 => "00000000",
	10556 => "00000000",
	10557 => "00000000",
	10558 => "00000000",
	10559 => "00000000",
	10560 => "00000000",
	10561 => "00000000",
	10562 => "00000000",
	10563 => "00000000",
	10564 => "00000000",
	10565 => "00000000",
	10566 => "00000000",
	10567 => "00000000",
	10568 => "00000000",
	10569 => "00000000",
	10570 => "00000000",
	10571 => "00000000",
	10572 => "00000000",
	10573 => "11111111",
	10574 => "11111111",
	10575 => "11111111",
	10576 => "11111111",
	10577 => "11111111",
	10578 => "11111111",
	10579 => "11111111",
	10580 => "11111111",
	10581 => "11111111",
	10582 => "11111111",
	10583 => "11111111",
	10584 => "00000000",
	10585 => "00000000",
	10586 => "00000000",
	10587 => "00000000",
	10588 => "00000000",
	10589 => "00000000",
	10590 => "00000000",
	10591 => "00000000",
	10592 => "00000000",
	10593 => "00000000",
	10594 => "00000000",
	10595 => "00000000",
	10596 => "00000000",
	10597 => "00000000",
	10598 => "00000000",
	10599 => "00000000",
	10600 => "00000000",
	10601 => "00000000",
	10602 => "00000000",
	10603 => "00000000",
	10604 => "00000000",
	10605 => "00000000",
	10606 => "00000000",
	10607 => "00000000",
	10608 => "00000000",
	10609 => "00000000",
	10610 => "00000000",
	10611 => "00000000",
	10612 => "00000000",
	10613 => "00000000",
	10614 => "00000000",
	10615 => "00000000",
	10624 => "00000000",
	10625 => "00000000",
	10626 => "00000000",
	10627 => "00000000",
	10628 => "00000000",
	10629 => "00000000",
	10630 => "00000000",
	10631 => "00000000",
	10632 => "00000000",
	10633 => "00000000",
	10634 => "00000000",
	10635 => "00000000",
	10636 => "00000000",
	10637 => "00000000",
	10638 => "00000000",
	10639 => "00000000",
	10640 => "00000000",
	10641 => "00000000",
	10642 => "00000000",
	10643 => "00000000",
	10644 => "00000000",
	10645 => "00000000",
	10646 => "00000000",
	10647 => "00000000",
	10648 => "00000000",
	10649 => "00000000",
	10650 => "00000000",
	10651 => "00000000",
	10652 => "00000000",
	10653 => "00000000",
	10654 => "00000000",
	10655 => "00000000",
	10656 => "11111111",
	10657 => "11111111",
	10658 => "11111111",
	10659 => "11111111",
	10660 => "11111111",
	10661 => "11111111",
	10662 => "11111111",
	10663 => "11111111",
	10664 => "11111111",
	10665 => "11111111",
	10666 => "11111111",
	10667 => "00000000",
	10668 => "00000000",
	10669 => "00000000",
	10670 => "00000000",
	10671 => "00000000",
	10672 => "00000000",
	10673 => "00000000",
	10674 => "00000000",
	10675 => "00000000",
	10676 => "00000000",
	10677 => "00000000",
	10678 => "00000000",
	10679 => "00000000",
	10680 => "00000000",
	10681 => "00000000",
	10682 => "00000000",
	10683 => "00000000",
	10684 => "00000000",
	10685 => "00000000",
	10686 => "00000000",
	10687 => "00000000",
	10688 => "00000000",
	10689 => "00000000",
	10690 => "00000000",
	10691 => "00000000",
	10692 => "00000000",
	10693 => "00000000",
	10694 => "00000000",
	10695 => "00000000",
	10696 => "00000000",
	10697 => "00000000",
	10698 => "00000000",
	10699 => "00000000",
	10700 => "00000000",
	10701 => "00000000",
	10702 => "11111111",
	10703 => "11111111",
	10704 => "11111111",
	10705 => "11111111",
	10706 => "11111111",
	10707 => "11111111",
	10708 => "11111111",
	10709 => "11111111",
	10710 => "11111111",
	10711 => "11111111",
	10712 => "11111111",
	10713 => "00000000",
	10714 => "00000000",
	10715 => "00000000",
	10716 => "00000000",
	10717 => "00000000",
	10718 => "00000000",
	10719 => "00000000",
	10720 => "00000000",
	10721 => "00000000",
	10722 => "00000000",
	10723 => "00000000",
	10724 => "00000000",
	10725 => "00000000",
	10726 => "00000000",
	10727 => "00000000",
	10728 => "00000000",
	10729 => "00000000",
	10730 => "00000000",
	10731 => "00000000",
	10732 => "00000000",
	10733 => "00000000",
	10734 => "00000000",
	10735 => "00000000",
	10736 => "00000000",
	10737 => "00000000",
	10738 => "00000000",
	10739 => "00000000",
	10740 => "00000000",
	10741 => "00000000",
	10742 => "00000000",
	10743 => "00000000",
	10752 => "00000000",
	10753 => "00000000",
	10754 => "00000000",
	10755 => "00000000",
	10756 => "00000000",
	10757 => "00000000",
	10758 => "00000000",
	10759 => "00000000",
	10760 => "00000000",
	10761 => "00000000",
	10762 => "00000000",
	10763 => "00000000",
	10764 => "00000000",
	10765 => "00000000",
	10766 => "00000000",
	10767 => "00000000",
	10768 => "00000000",
	10769 => "00000000",
	10770 => "00000000",
	10771 => "00000000",
	10772 => "00000000",
	10773 => "00000000",
	10774 => "00000000",
	10775 => "00000000",
	10776 => "00000000",
	10777 => "00000000",
	10778 => "00000000",
	10779 => "00000000",
	10780 => "00000000",
	10781 => "00000000",
	10782 => "00000000",
	10783 => "11111111",
	10784 => "11111111",
	10785 => "11111111",
	10786 => "11111111",
	10787 => "11111111",
	10788 => "11111111",
	10789 => "11111111",
	10790 => "11111111",
	10791 => "11111111",
	10792 => "11111111",
	10793 => "11111111",
	10794 => "00000000",
	10795 => "00000000",
	10796 => "00000000",
	10797 => "00000000",
	10798 => "00000000",
	10799 => "00000000",
	10800 => "00000000",
	10801 => "00000000",
	10802 => "00000000",
	10803 => "00000000",
	10804 => "00000000",
	10805 => "00000000",
	10806 => "00000000",
	10807 => "00000000",
	10808 => "00000000",
	10809 => "00000000",
	10810 => "00000000",
	10811 => "00000000",
	10812 => "00000000",
	10813 => "00000000",
	10814 => "00000000",
	10815 => "00000000",
	10816 => "00000000",
	10817 => "00000000",
	10818 => "00000000",
	10819 => "00000000",
	10820 => "00000000",
	10821 => "00000000",
	10822 => "00000000",
	10823 => "00000000",
	10824 => "00000000",
	10825 => "00000000",
	10826 => "00000000",
	10827 => "00000000",
	10828 => "00000000",
	10829 => "00000000",
	10830 => "00000000",
	10831 => "11111111",
	10832 => "11111111",
	10833 => "11111111",
	10834 => "11111111",
	10835 => "11111111",
	10836 => "11111111",
	10837 => "11111111",
	10838 => "11111111",
	10839 => "11111111",
	10840 => "11111111",
	10841 => "11111111",
	10842 => "00000000",
	10843 => "00000000",
	10844 => "00000000",
	10845 => "00000000",
	10846 => "00000000",
	10847 => "00000000",
	10848 => "00000000",
	10849 => "00000000",
	10850 => "00000000",
	10851 => "00000000",
	10852 => "00000000",
	10853 => "00000000",
	10854 => "00000000",
	10855 => "00000000",
	10856 => "00000000",
	10857 => "00000000",
	10858 => "00000000",
	10859 => "00000000",
	10860 => "00000000",
	10861 => "00000000",
	10862 => "00000000",
	10863 => "00000000",
	10864 => "00000000",
	10865 => "00000000",
	10866 => "00000000",
	10867 => "00000000",
	10868 => "00000000",
	10869 => "00000000",
	10870 => "00000000",
	10871 => "00000000",
	10880 => "00000000",
	10881 => "00000000",
	10882 => "00000000",
	10883 => "00000000",
	10884 => "00000000",
	10885 => "00000000",
	10886 => "00000000",
	10887 => "00000000",
	10888 => "00000000",
	10889 => "00000000",
	10890 => "00000000",
	10891 => "00000000",
	10892 => "00000000",
	10893 => "00000000",
	10894 => "00000000",
	10895 => "00000000",
	10896 => "00000000",
	10897 => "00000000",
	10898 => "00000000",
	10899 => "00000000",
	10900 => "00000000",
	10901 => "00000000",
	10902 => "00000000",
	10903 => "00000000",
	10904 => "00000000",
	10905 => "00000000",
	10906 => "00000000",
	10907 => "00000000",
	10908 => "00000000",
	10909 => "00000000",
	10910 => "11111111",
	10911 => "11111111",
	10912 => "11111111",
	10913 => "11111111",
	10914 => "11111111",
	10915 => "11111111",
	10916 => "11111111",
	10917 => "11111111",
	10918 => "11111111",
	10919 => "11111111",
	10920 => "11111111",
	10921 => "00000000",
	10922 => "00000000",
	10923 => "00000000",
	10924 => "00000000",
	10925 => "00000000",
	10926 => "00000000",
	10927 => "00000000",
	10928 => "00000000",
	10929 => "00000000",
	10930 => "00000000",
	10931 => "00000000",
	10932 => "00000000",
	10933 => "00000000",
	10934 => "00000000",
	10935 => "00000000",
	10936 => "00000000",
	10937 => "00000000",
	10938 => "00000000",
	10939 => "00000000",
	10940 => "00000000",
	10941 => "00000000",
	10942 => "00000000",
	10943 => "00000000",
	10944 => "00000000",
	10945 => "00000000",
	10946 => "00000000",
	10947 => "00000000",
	10948 => "00000000",
	10949 => "00000000",
	10950 => "00000000",
	10951 => "00000000",
	10952 => "00000000",
	10953 => "00000000",
	10954 => "00000000",
	10955 => "00000000",
	10956 => "00000000",
	10957 => "00000000",
	10958 => "00000000",
	10959 => "00000000",
	10960 => "11111111",
	10961 => "11111111",
	10962 => "11111111",
	10963 => "11111111",
	10964 => "11111111",
	10965 => "11111111",
	10966 => "11111111",
	10967 => "11111111",
	10968 => "11111111",
	10969 => "11111111",
	10970 => "11111111",
	10971 => "00000000",
	10972 => "00000000",
	10973 => "00000000",
	10974 => "00000000",
	10975 => "00000000",
	10976 => "00000000",
	10977 => "00000000",
	10978 => "00000000",
	10979 => "00000000",
	10980 => "00000000",
	10981 => "00000000",
	10982 => "00000000",
	10983 => "00000000",
	10984 => "00000000",
	10985 => "00000000",
	10986 => "00000000",
	10987 => "00000000",
	10988 => "00000000",
	10989 => "00000000",
	10990 => "00000000",
	10991 => "00000000",
	10992 => "00000000",
	10993 => "00000000",
	10994 => "00000000",
	10995 => "00000000",
	10996 => "00000000",
	10997 => "00000000",
	10998 => "00000000",
	10999 => "00000000",
	11008 => "00000000",
	11009 => "00000000",
	11010 => "00000000",
	11011 => "00000000",
	11012 => "00000000",
	11013 => "00000000",
	11014 => "00000000",
	11015 => "00000000",
	11016 => "00000000",
	11017 => "00000000",
	11018 => "00000000",
	11019 => "00000000",
	11020 => "00000000",
	11021 => "00000000",
	11022 => "00000000",
	11023 => "00000000",
	11024 => "00000000",
	11025 => "00000000",
	11026 => "00000000",
	11027 => "00000000",
	11028 => "00000000",
	11029 => "00000000",
	11030 => "00000000",
	11031 => "00000000",
	11032 => "00000000",
	11033 => "00000000",
	11034 => "00000000",
	11035 => "00000000",
	11036 => "00000000",
	11037 => "11111111",
	11038 => "11111111",
	11039 => "11111111",
	11040 => "11111111",
	11041 => "11111111",
	11042 => "11111111",
	11043 => "11111111",
	11044 => "11111111",
	11045 => "11111111",
	11046 => "11111111",
	11047 => "11111111",
	11048 => "00000000",
	11049 => "00000000",
	11050 => "00000000",
	11051 => "00000000",
	11052 => "00000000",
	11053 => "00000000",
	11054 => "00000000",
	11055 => "00000000",
	11056 => "00000000",
	11057 => "00000000",
	11058 => "00000000",
	11059 => "00000000",
	11060 => "00000000",
	11061 => "00000000",
	11062 => "00000000",
	11063 => "00000000",
	11064 => "00000000",
	11065 => "00000000",
	11066 => "00000000",
	11067 => "00000000",
	11068 => "00000000",
	11069 => "00000000",
	11070 => "00000000",
	11071 => "00000000",
	11072 => "00000000",
	11073 => "00000000",
	11074 => "00000000",
	11075 => "00000000",
	11076 => "00000000",
	11077 => "00000000",
	11078 => "00000000",
	11079 => "00000000",
	11080 => "00000000",
	11081 => "00000000",
	11082 => "00000000",
	11083 => "00000000",
	11084 => "00000000",
	11085 => "00000000",
	11086 => "00000000",
	11087 => "00000000",
	11088 => "00000000",
	11089 => "11111111",
	11090 => "11111111",
	11091 => "11111111",
	11092 => "11111111",
	11093 => "11111111",
	11094 => "11111111",
	11095 => "11111111",
	11096 => "11111111",
	11097 => "11111111",
	11098 => "11111111",
	11099 => "11111111",
	11100 => "00000000",
	11101 => "00000000",
	11102 => "00000000",
	11103 => "00000000",
	11104 => "00000000",
	11105 => "00000000",
	11106 => "00000000",
	11107 => "00000000",
	11108 => "00000000",
	11109 => "00000000",
	11110 => "00000000",
	11111 => "00000000",
	11112 => "00000000",
	11113 => "00000000",
	11114 => "00000000",
	11115 => "00000000",
	11116 => "00000000",
	11117 => "00000000",
	11118 => "00000000",
	11119 => "00000000",
	11120 => "00000000",
	11121 => "00000000",
	11122 => "00000000",
	11123 => "00000000",
	11124 => "00000000",
	11125 => "00000000",
	11126 => "00000000",
	11127 => "00000000",
	11136 => "00000000",
	11137 => "00000000",
	11138 => "00000000",
	11139 => "00000000",
	11140 => "00000000",
	11141 => "00000000",
	11142 => "00000000",
	11143 => "00000000",
	11144 => "00000000",
	11145 => "00000000",
	11146 => "00000000",
	11147 => "00000000",
	11148 => "00000000",
	11149 => "00000000",
	11150 => "00000000",
	11151 => "00000000",
	11152 => "00000000",
	11153 => "00000000",
	11154 => "00000000",
	11155 => "00000000",
	11156 => "00000000",
	11157 => "00000000",
	11158 => "00000000",
	11159 => "00000000",
	11160 => "00000000",
	11161 => "00000000",
	11162 => "00000000",
	11163 => "00000000",
	11164 => "11111111",
	11165 => "11111111",
	11166 => "11111111",
	11167 => "11111111",
	11168 => "11111111",
	11169 => "11111111",
	11170 => "11111111",
	11171 => "11111111",
	11172 => "11111111",
	11173 => "11111111",
	11174 => "11111111",
	11175 => "00000000",
	11176 => "00000000",
	11177 => "00000000",
	11178 => "00000000",
	11179 => "00000000",
	11180 => "00000000",
	11181 => "00000000",
	11182 => "00000000",
	11183 => "00000000",
	11184 => "00000000",
	11185 => "00000000",
	11186 => "00000000",
	11187 => "00000000",
	11188 => "00000000",
	11189 => "00000000",
	11190 => "00000000",
	11191 => "00000000",
	11192 => "00000000",
	11193 => "00000000",
	11194 => "00000000",
	11195 => "00000000",
	11196 => "00000000",
	11197 => "00000000",
	11198 => "00000000",
	11199 => "00000000",
	11200 => "00000000",
	11201 => "00000000",
	11202 => "00000000",
	11203 => "00000000",
	11204 => "00000000",
	11205 => "00000000",
	11206 => "00000000",
	11207 => "00000000",
	11208 => "00000000",
	11209 => "00000000",
	11210 => "00000000",
	11211 => "00000000",
	11212 => "00000000",
	11213 => "00000000",
	11214 => "00000000",
	11215 => "00000000",
	11216 => "00000000",
	11217 => "00000000",
	11218 => "11111111",
	11219 => "11111111",
	11220 => "11111111",
	11221 => "11111111",
	11222 => "11111111",
	11223 => "11111111",
	11224 => "11111111",
	11225 => "11111111",
	11226 => "11111111",
	11227 => "11111111",
	11228 => "11111111",
	11229 => "00000000",
	11230 => "00000000",
	11231 => "00000000",
	11232 => "00000000",
	11233 => "00000000",
	11234 => "00000000",
	11235 => "00000000",
	11236 => "00000000",
	11237 => "00000000",
	11238 => "00000000",
	11239 => "00000000",
	11240 => "00000000",
	11241 => "00000000",
	11242 => "00000000",
	11243 => "00000000",
	11244 => "00000000",
	11245 => "00000000",
	11246 => "00000000",
	11247 => "00000000",
	11248 => "00000000",
	11249 => "00000000",
	11250 => "00000000",
	11251 => "00000000",
	11252 => "00000000",
	11253 => "00000000",
	11254 => "00000000",
	11255 => "00000000",
	11264 => "00000000",
	11265 => "00000000",
	11266 => "00000000",
	11267 => "00000000",
	11268 => "00000000",
	11269 => "00000000",
	11270 => "00000000",
	11271 => "00000000",
	11272 => "00000000",
	11273 => "00000000",
	11274 => "00000000",
	11275 => "00000000",
	11276 => "00000000",
	11277 => "00000000",
	11278 => "00000000",
	11279 => "00000000",
	11280 => "00000000",
	11281 => "00000000",
	11282 => "00000000",
	11283 => "00000000",
	11284 => "00000000",
	11285 => "00000000",
	11286 => "00000000",
	11287 => "00000000",
	11288 => "00000000",
	11289 => "00000000",
	11290 => "00000000",
	11291 => "11111111",
	11292 => "11111111",
	11293 => "11111111",
	11294 => "11111111",
	11295 => "11111111",
	11296 => "11111111",
	11297 => "11111111",
	11298 => "11111111",
	11299 => "11111111",
	11300 => "11111111",
	11301 => "11111111",
	11302 => "00000000",
	11303 => "00000000",
	11304 => "00000000",
	11305 => "00000000",
	11306 => "00000000",
	11307 => "00000000",
	11308 => "00000000",
	11309 => "00000000",
	11310 => "00000000",
	11311 => "00000000",
	11312 => "00000000",
	11313 => "00000000",
	11314 => "00000000",
	11315 => "00000000",
	11316 => "00000000",
	11317 => "00000000",
	11318 => "00000000",
	11319 => "00000000",
	11320 => "00000000",
	11321 => "00000000",
	11322 => "00000000",
	11323 => "00000000",
	11324 => "00000000",
	11325 => "00000000",
	11326 => "00000000",
	11327 => "00000000",
	11328 => "00000000",
	11329 => "00000000",
	11330 => "00000000",
	11331 => "00000000",
	11332 => "00000000",
	11333 => "00000000",
	11334 => "00000000",
	11335 => "00000000",
	11336 => "00000000",
	11337 => "00000000",
	11338 => "00000000",
	11339 => "00000000",
	11340 => "00000000",
	11341 => "00000000",
	11342 => "00000000",
	11343 => "00000000",
	11344 => "00000000",
	11345 => "00000000",
	11346 => "00000000",
	11347 => "11111111",
	11348 => "11111111",
	11349 => "11111111",
	11350 => "11111111",
	11351 => "11111111",
	11352 => "11111111",
	11353 => "11111111",
	11354 => "11111111",
	11355 => "11111111",
	11356 => "11111111",
	11357 => "11111111",
	11358 => "00000000",
	11359 => "00000000",
	11360 => "00000000",
	11361 => "00000000",
	11362 => "00000000",
	11363 => "00000000",
	11364 => "00000000",
	11365 => "00000000",
	11366 => "00000000",
	11367 => "00000000",
	11368 => "00000000",
	11369 => "00000000",
	11370 => "00000000",
	11371 => "00000000",
	11372 => "00000000",
	11373 => "00000000",
	11374 => "00000000",
	11375 => "00000000",
	11376 => "00000000",
	11377 => "00000000",
	11378 => "00000000",
	11379 => "00000000",
	11380 => "00000000",
	11381 => "00000000",
	11382 => "00000000",
	11383 => "00000000",
	11392 => "00000000",
	11393 => "00000000",
	11394 => "00000000",
	11395 => "00000000",
	11396 => "00000000",
	11397 => "00000000",
	11398 => "00000000",
	11399 => "00000000",
	11400 => "00000000",
	11401 => "00000000",
	11402 => "00000000",
	11403 => "00000000",
	11404 => "00000000",
	11405 => "00000000",
	11406 => "00000000",
	11407 => "00000000",
	11408 => "00000000",
	11409 => "00000000",
	11410 => "00000000",
	11411 => "00000000",
	11412 => "00000000",
	11413 => "00000000",
	11414 => "00000000",
	11415 => "00000000",
	11416 => "00000000",
	11417 => "00000000",
	11418 => "11111111",
	11419 => "11111111",
	11420 => "11111111",
	11421 => "11111111",
	11422 => "11111111",
	11423 => "11111111",
	11424 => "11111111",
	11425 => "11111111",
	11426 => "11111111",
	11427 => "11111111",
	11428 => "11111111",
	11429 => "00000000",
	11430 => "00000000",
	11431 => "00000000",
	11432 => "00000000",
	11433 => "00000000",
	11434 => "00000000",
	11435 => "00000000",
	11436 => "00000000",
	11437 => "00000000",
	11438 => "00000000",
	11439 => "00000000",
	11440 => "00000000",
	11441 => "00000000",
	11442 => "00000000",
	11443 => "00000000",
	11444 => "00000000",
	11445 => "00000000",
	11446 => "00000000",
	11447 => "00000000",
	11448 => "00000000",
	11449 => "00000000",
	11450 => "00000000",
	11451 => "00000000",
	11452 => "00000000",
	11453 => "00000000",
	11454 => "00000000",
	11455 => "00000000",
	11456 => "00000000",
	11457 => "00000000",
	11458 => "00000000",
	11459 => "00000000",
	11460 => "00000000",
	11461 => "00000000",
	11462 => "00000000",
	11463 => "00000000",
	11464 => "00000000",
	11465 => "00000000",
	11466 => "00000000",
	11467 => "00000000",
	11468 => "00000000",
	11469 => "00000000",
	11470 => "00000000",
	11471 => "00000000",
	11472 => "00000000",
	11473 => "00000000",
	11474 => "00000000",
	11475 => "00000000",
	11476 => "11111111",
	11477 => "11111111",
	11478 => "11111111",
	11479 => "11111111",
	11480 => "11111111",
	11481 => "11111111",
	11482 => "11111111",
	11483 => "11111111",
	11484 => "11111111",
	11485 => "11111111",
	11486 => "11111111",
	11487 => "00000000",
	11488 => "00000000",
	11489 => "00000000",
	11490 => "00000000",
	11491 => "00000000",
	11492 => "00000000",
	11493 => "00000000",
	11494 => "00000000",
	11495 => "00000000",
	11496 => "00000000",
	11497 => "00000000",
	11498 => "00000000",
	11499 => "00000000",
	11500 => "00000000",
	11501 => "00000000",
	11502 => "00000000",
	11503 => "00000000",
	11504 => "00000000",
	11505 => "00000000",
	11506 => "00000000",
	11507 => "00000000",
	11508 => "00000000",
	11509 => "00000000",
	11510 => "00000000",
	11511 => "00000000",
	11520 => "00000000",
	11521 => "00000000",
	11522 => "00000000",
	11523 => "00000000",
	11524 => "00000000",
	11525 => "00000000",
	11526 => "00000000",
	11527 => "00000000",
	11528 => "00000000",
	11529 => "00000000",
	11530 => "00000000",
	11531 => "00000000",
	11532 => "00000000",
	11533 => "00000000",
	11534 => "00000000",
	11535 => "00000000",
	11536 => "00000000",
	11537 => "00000000",
	11538 => "00000000",
	11539 => "00000000",
	11540 => "00000000",
	11541 => "00000000",
	11542 => "00000000",
	11543 => "00000000",
	11544 => "00000000",
	11545 => "11111111",
	11546 => "11111111",
	11547 => "11111111",
	11548 => "11111111",
	11549 => "11111111",
	11550 => "11111111",
	11551 => "11111111",
	11552 => "11111111",
	11553 => "11111111",
	11554 => "11111111",
	11555 => "11111111",
	11556 => "00000000",
	11557 => "00000000",
	11558 => "00000000",
	11559 => "00000000",
	11560 => "00000000",
	11561 => "00000000",
	11562 => "00000000",
	11563 => "00000000",
	11564 => "00000000",
	11565 => "00000000",
	11566 => "00000000",
	11567 => "00000000",
	11568 => "00000000",
	11569 => "00000000",
	11570 => "00000000",
	11571 => "00000000",
	11572 => "00000000",
	11573 => "00000000",
	11574 => "00000000",
	11575 => "00000000",
	11576 => "00000000",
	11577 => "00000000",
	11578 => "00000000",
	11579 => "00000000",
	11580 => "00000000",
	11581 => "00000000",
	11582 => "00000000",
	11583 => "00000000",
	11584 => "00000000",
	11585 => "00000000",
	11586 => "00000000",
	11587 => "00000000",
	11588 => "00000000",
	11589 => "00000000",
	11590 => "00000000",
	11591 => "00000000",
	11592 => "00000000",
	11593 => "00000000",
	11594 => "00000000",
	11595 => "00000000",
	11596 => "00000000",
	11597 => "00000000",
	11598 => "00000000",
	11599 => "00000000",
	11600 => "00000000",
	11601 => "00000000",
	11602 => "00000000",
	11603 => "00000000",
	11604 => "00000000",
	11605 => "11111111",
	11606 => "11111111",
	11607 => "11111111",
	11608 => "11111111",
	11609 => "11111111",
	11610 => "11111111",
	11611 => "11111111",
	11612 => "11111111",
	11613 => "11111111",
	11614 => "11111111",
	11615 => "11111111",
	11616 => "00000000",
	11617 => "00000000",
	11618 => "00000000",
	11619 => "00000000",
	11620 => "00000000",
	11621 => "00000000",
	11622 => "00000000",
	11623 => "00000000",
	11624 => "00000000",
	11625 => "00000000",
	11626 => "00000000",
	11627 => "00000000",
	11628 => "00000000",
	11629 => "00000000",
	11630 => "00000000",
	11631 => "00000000",
	11632 => "00000000",
	11633 => "00000000",
	11634 => "00000000",
	11635 => "00000000",
	11636 => "00000000",
	11637 => "00000000",
	11638 => "00000000",
	11639 => "00000000",
	11648 => "00000000",
	11649 => "00000000",
	11650 => "00000000",
	11651 => "00000000",
	11652 => "00000000",
	11653 => "00000000",
	11654 => "00000000",
	11655 => "00000000",
	11656 => "00000000",
	11657 => "00000000",
	11658 => "00000000",
	11659 => "00000000",
	11660 => "00000000",
	11661 => "00000000",
	11662 => "00000000",
	11663 => "00000000",
	11664 => "00000000",
	11665 => "00000000",
	11666 => "00000000",
	11667 => "00000000",
	11668 => "00000000",
	11669 => "00000000",
	11670 => "00000000",
	11671 => "00000000",
	11672 => "11111111",
	11673 => "11111111",
	11674 => "11111111",
	11675 => "11111111",
	11676 => "11111111",
	11677 => "11111111",
	11678 => "11111111",
	11679 => "11111111",
	11680 => "11111111",
	11681 => "11111111",
	11682 => "11111111",
	11683 => "00000000",
	11684 => "00000000",
	11685 => "00000000",
	11686 => "00000000",
	11687 => "00000000",
	11688 => "00000000",
	11689 => "00000000",
	11690 => "00000000",
	11691 => "00000000",
	11692 => "00000000",
	11693 => "00000000",
	11694 => "00000000",
	11695 => "00000000",
	11696 => "00000000",
	11697 => "00000000",
	11698 => "00000000",
	11699 => "00000000",
	11700 => "00000000",
	11701 => "00000000",
	11702 => "00000000",
	11703 => "00000000",
	11704 => "00000000",
	11705 => "00000000",
	11706 => "00000000",
	11707 => "00000000",
	11708 => "00000000",
	11709 => "00000000",
	11710 => "00000000",
	11711 => "00000000",
	11712 => "00000000",
	11713 => "00000000",
	11714 => "00000000",
	11715 => "00000000",
	11716 => "00000000",
	11717 => "00000000",
	11718 => "00000000",
	11719 => "00000000",
	11720 => "00000000",
	11721 => "00000000",
	11722 => "00000000",
	11723 => "00000000",
	11724 => "00000000",
	11725 => "00000000",
	11726 => "00000000",
	11727 => "00000000",
	11728 => "00000000",
	11729 => "00000000",
	11730 => "00000000",
	11731 => "00000000",
	11732 => "00000000",
	11733 => "00000000",
	11734 => "11111111",
	11735 => "11111111",
	11736 => "11111111",
	11737 => "11111111",
	11738 => "11111111",
	11739 => "11111111",
	11740 => "11111111",
	11741 => "11111111",
	11742 => "11111111",
	11743 => "11111111",
	11744 => "11111111",
	11745 => "00000000",
	11746 => "00000000",
	11747 => "00000000",
	11748 => "00000000",
	11749 => "00000000",
	11750 => "00000000",
	11751 => "00000000",
	11752 => "00000000",
	11753 => "00000000",
	11754 => "00000000",
	11755 => "00000000",
	11756 => "00000000",
	11757 => "00000000",
	11758 => "00000000",
	11759 => "00000000",
	11760 => "00000000",
	11761 => "00000000",
	11762 => "00000000",
	11763 => "00000000",
	11764 => "00000000",
	11765 => "00000000",
	11766 => "00000000",
	11767 => "00000000",
	11776 => "00000000",
	11777 => "00000000",
	11778 => "00000000",
	11779 => "00000000",
	11780 => "00000000",
	11781 => "00000000",
	11782 => "00000000",
	11783 => "00000000",
	11784 => "00000000",
	11785 => "00000000",
	11786 => "00000000",
	11787 => "00000000",
	11788 => "00000000",
	11789 => "00000000",
	11790 => "00000000",
	11791 => "00000000",
	11792 => "00000000",
	11793 => "00000000",
	11794 => "00000000",
	11795 => "00000000",
	11796 => "00000000",
	11797 => "00000000",
	11798 => "00000000",
	11799 => "11111111",
	11800 => "11111111",
	11801 => "11111111",
	11802 => "11111111",
	11803 => "11111111",
	11804 => "11111111",
	11805 => "11111111",
	11806 => "11111111",
	11807 => "11111111",
	11808 => "11111111",
	11809 => "11111111",
	11810 => "00000000",
	11811 => "00000000",
	11812 => "00000000",
	11813 => "00000000",
	11814 => "00000000",
	11815 => "00000000",
	11816 => "00000000",
	11817 => "00000000",
	11818 => "00000000",
	11819 => "00000000",
	11820 => "00000000",
	11821 => "00000000",
	11822 => "00000000",
	11823 => "00000000",
	11824 => "00000000",
	11825 => "00000000",
	11826 => "00000000",
	11827 => "00000000",
	11828 => "00000000",
	11829 => "00000000",
	11830 => "00000000",
	11831 => "00000000",
	11832 => "00000000",
	11833 => "00000000",
	11834 => "00000000",
	11835 => "00000000",
	11836 => "00000000",
	11837 => "00000000",
	11838 => "00000000",
	11839 => "00000000",
	11840 => "00000000",
	11841 => "00000000",
	11842 => "00000000",
	11843 => "00000000",
	11844 => "00000000",
	11845 => "00000000",
	11846 => "00000000",
	11847 => "00000000",
	11848 => "00000000",
	11849 => "00000000",
	11850 => "00000000",
	11851 => "00000000",
	11852 => "00000000",
	11853 => "00000000",
	11854 => "00000000",
	11855 => "00000000",
	11856 => "00000000",
	11857 => "00000000",
	11858 => "00000000",
	11859 => "00000000",
	11860 => "00000000",
	11861 => "00000000",
	11862 => "00000000",
	11863 => "11111111",
	11864 => "11111111",
	11865 => "11111111",
	11866 => "11111111",
	11867 => "11111111",
	11868 => "11111111",
	11869 => "11111111",
	11870 => "11111111",
	11871 => "11111111",
	11872 => "11111111",
	11873 => "11111111",
	11874 => "00000000",
	11875 => "00000000",
	11876 => "00000000",
	11877 => "00000000",
	11878 => "00000000",
	11879 => "00000000",
	11880 => "00000000",
	11881 => "00000000",
	11882 => "00000000",
	11883 => "00000000",
	11884 => "00000000",
	11885 => "00000000",
	11886 => "00000000",
	11887 => "00000000",
	11888 => "00000000",
	11889 => "00000000",
	11890 => "00000000",
	11891 => "00000000",
	11892 => "00000000",
	11893 => "00000000",
	11894 => "00000000",
	11895 => "00000000",
	11904 => "00000000",
	11905 => "00000000",
	11906 => "00000000",
	11907 => "00000000",
	11908 => "00000000",
	11909 => "00000000",
	11910 => "00000000",
	11911 => "00000000",
	11912 => "00000000",
	11913 => "00000000",
	11914 => "00000000",
	11915 => "00000000",
	11916 => "00000000",
	11917 => "00000000",
	11918 => "00000000",
	11919 => "00000000",
	11920 => "00000000",
	11921 => "00000000",
	11922 => "00000000",
	11923 => "00000000",
	11924 => "00000000",
	11925 => "00000000",
	11926 => "11111111",
	11927 => "11111111",
	11928 => "11111111",
	11929 => "11111111",
	11930 => "11111111",
	11931 => "11111111",
	11932 => "11111111",
	11933 => "11111111",
	11934 => "11111111",
	11935 => "11111111",
	11936 => "11111111",
	11937 => "00000000",
	11938 => "00000000",
	11939 => "00000000",
	11940 => "00000000",
	11941 => "00000000",
	11942 => "00000000",
	11943 => "00000000",
	11944 => "00000000",
	11945 => "00000000",
	11946 => "00000000",
	11947 => "00000000",
	11948 => "00000000",
	11949 => "00000000",
	11950 => "00000000",
	11951 => "00000000",
	11952 => "00000000",
	11953 => "00000000",
	11954 => "00000000",
	11955 => "00000000",
	11956 => "00000000",
	11957 => "00000000",
	11958 => "00000000",
	11959 => "00000000",
	11960 => "00000000",
	11961 => "00000000",
	11962 => "00000000",
	11963 => "00000000",
	11964 => "00000000",
	11965 => "00000000",
	11966 => "00000000",
	11967 => "00000000",
	11968 => "00000000",
	11969 => "00000000",
	11970 => "00000000",
	11971 => "00000000",
	11972 => "00000000",
	11973 => "00000000",
	11974 => "00000000",
	11975 => "00000000",
	11976 => "00000000",
	11977 => "00000000",
	11978 => "00000000",
	11979 => "00000000",
	11980 => "00000000",
	11981 => "00000000",
	11982 => "00000000",
	11983 => "00000000",
	11984 => "00000000",
	11985 => "00000000",
	11986 => "00000000",
	11987 => "00000000",
	11988 => "00000000",
	11989 => "00000000",
	11990 => "00000000",
	11991 => "00000000",
	11992 => "11111111",
	11993 => "11111111",
	11994 => "11111111",
	11995 => "11111111",
	11996 => "11111111",
	11997 => "11111111",
	11998 => "11111111",
	11999 => "11111111",
	12000 => "11111111",
	12001 => "11111111",
	12002 => "11111111",
	12003 => "00000000",
	12004 => "00000000",
	12005 => "00000000",
	12006 => "00000000",
	12007 => "00000000",
	12008 => "00000000",
	12009 => "00000000",
	12010 => "00000000",
	12011 => "00000000",
	12012 => "00000000",
	12013 => "00000000",
	12014 => "00000000",
	12015 => "00000000",
	12016 => "00000000",
	12017 => "00000000",
	12018 => "00000000",
	12019 => "00000000",
	12020 => "00000000",
	12021 => "00000000",
	12022 => "00000000",
	12023 => "00000000",
	12032 => "00000000",
	12033 => "00000000",
	12034 => "00000000",
	12035 => "00000000",
	12036 => "00000000",
	12037 => "00000000",
	12038 => "00000000",
	12039 => "00000000",
	12040 => "00000000",
	12041 => "00000000",
	12042 => "00000000",
	12043 => "00000000",
	12044 => "00000000",
	12045 => "00000000",
	12046 => "00000000",
	12047 => "00000000",
	12048 => "00000000",
	12049 => "00000000",
	12050 => "00000000",
	12051 => "00000000",
	12052 => "00000000",
	12053 => "11111111",
	12054 => "11111111",
	12055 => "11111111",
	12056 => "11111111",
	12057 => "11111111",
	12058 => "11111111",
	12059 => "11111111",
	12060 => "11111111",
	12061 => "11111111",
	12062 => "11111111",
	12063 => "11111111",
	12064 => "00000000",
	12065 => "00000000",
	12066 => "00000000",
	12067 => "00000000",
	12068 => "00000000",
	12069 => "00000000",
	12070 => "00000000",
	12071 => "00000000",
	12072 => "00000000",
	12073 => "00000000",
	12074 => "00000000",
	12075 => "00000000",
	12076 => "00000000",
	12077 => "00000000",
	12078 => "00000000",
	12079 => "00000000",
	12080 => "00000000",
	12081 => "00000000",
	12082 => "00000000",
	12083 => "00000000",
	12084 => "00000000",
	12085 => "00000000",
	12086 => "00000000",
	12087 => "00000000",
	12088 => "00000000",
	12089 => "00000000",
	12090 => "00000000",
	12091 => "00000000",
	12092 => "00000000",
	12093 => "00000000",
	12094 => "00000000",
	12095 => "00000000",
	12096 => "00000000",
	12097 => "00000000",
	12098 => "00000000",
	12099 => "00000000",
	12100 => "00000000",
	12101 => "00000000",
	12102 => "00000000",
	12103 => "00000000",
	12104 => "00000000",
	12105 => "00000000",
	12106 => "00000000",
	12107 => "00000000",
	12108 => "00000000",
	12109 => "00000000",
	12110 => "00000000",
	12111 => "00000000",
	12112 => "00000000",
	12113 => "00000000",
	12114 => "00000000",
	12115 => "00000000",
	12116 => "00000000",
	12117 => "00000000",
	12118 => "00000000",
	12119 => "00000000",
	12120 => "00000000",
	12121 => "11111111",
	12122 => "11111111",
	12123 => "11111111",
	12124 => "11111111",
	12125 => "11111111",
	12126 => "11111111",
	12127 => "11111111",
	12128 => "11111111",
	12129 => "11111111",
	12130 => "11111111",
	12131 => "11111111",
	12132 => "00000000",
	12133 => "00000000",
	12134 => "00000000",
	12135 => "00000000",
	12136 => "00000000",
	12137 => "00000000",
	12138 => "00000000",
	12139 => "00000000",
	12140 => "00000000",
	12141 => "00000000",
	12142 => "00000000",
	12143 => "00000000",
	12144 => "00000000",
	12145 => "00000000",
	12146 => "00000000",
	12147 => "00000000",
	12148 => "00000000",
	12149 => "00000000",
	12150 => "00000000",
	12151 => "00000000",
	12160 => "00000000",
	12161 => "00000000",
	12162 => "00000000",
	12163 => "00000000",
	12164 => "00000000",
	12165 => "00000000",
	12166 => "00000000",
	12167 => "00000000",
	12168 => "00000000",
	12169 => "00000000",
	12170 => "00000000",
	12171 => "00000000",
	12172 => "00000000",
	12173 => "00000000",
	12174 => "00000000",
	12175 => "00000000",
	12176 => "00000000",
	12177 => "00000000",
	12178 => "00000000",
	12179 => "00000000",
	12180 => "11111111",
	12181 => "11111111",
	12182 => "11111111",
	12183 => "11111111",
	12184 => "11111111",
	12185 => "11111111",
	12186 => "11111111",
	12187 => "11111111",
	12188 => "11111111",
	12189 => "11111111",
	12190 => "11111111",
	12191 => "00000000",
	12192 => "00000000",
	12193 => "00000000",
	12194 => "00000000",
	12195 => "00000000",
	12196 => "00000000",
	12197 => "00000000",
	12198 => "00000000",
	12199 => "00000000",
	12200 => "00000000",
	12201 => "00000000",
	12202 => "00000000",
	12203 => "00000000",
	12204 => "00000000",
	12205 => "00000000",
	12206 => "00000000",
	12207 => "00000000",
	12208 => "00000000",
	12209 => "00000000",
	12210 => "00000000",
	12211 => "00000000",
	12212 => "00000000",
	12213 => "00000000",
	12214 => "00000000",
	12215 => "00000000",
	12216 => "00000000",
	12217 => "00000000",
	12218 => "00000000",
	12219 => "00000000",
	12220 => "00000000",
	12221 => "00000000",
	12222 => "00000000",
	12223 => "00000000",
	12224 => "00000000",
	12225 => "00000000",
	12226 => "00000000",
	12227 => "00000000",
	12228 => "00000000",
	12229 => "00000000",
	12230 => "00000000",
	12231 => "00000000",
	12232 => "00000000",
	12233 => "00000000",
	12234 => "00000000",
	12235 => "00000000",
	12236 => "00000000",
	12237 => "00000000",
	12238 => "00000000",
	12239 => "00000000",
	12240 => "00000000",
	12241 => "00000000",
	12242 => "00000000",
	12243 => "00000000",
	12244 => "00000000",
	12245 => "00000000",
	12246 => "00000000",
	12247 => "00000000",
	12248 => "00000000",
	12249 => "00000000",
	12250 => "11111111",
	12251 => "11111111",
	12252 => "11111111",
	12253 => "11111111",
	12254 => "11111111",
	12255 => "11111111",
	12256 => "11111111",
	12257 => "11111111",
	12258 => "11111111",
	12259 => "11111111",
	12260 => "11111111",
	12261 => "00000000",
	12262 => "00000000",
	12263 => "00000000",
	12264 => "00000000",
	12265 => "00000000",
	12266 => "00000000",
	12267 => "00000000",
	12268 => "00000000",
	12269 => "00000000",
	12270 => "00000000",
	12271 => "00000000",
	12272 => "00000000",
	12273 => "00000000",
	12274 => "00000000",
	12275 => "00000000",
	12276 => "00000000",
	12277 => "00000000",
	12278 => "00000000",
	12279 => "00000000",
	12288 => "00000000",
	12289 => "00000000",
	12290 => "00000000",
	12291 => "00000000",
	12292 => "00000000",
	12293 => "00000000",
	12294 => "00000000",
	12295 => "00000000",
	12296 => "00000000",
	12297 => "00000000",
	12298 => "00000000",
	12299 => "00000000",
	12300 => "00000000",
	12301 => "00000000",
	12302 => "00000000",
	12303 => "00000000",
	12304 => "00000000",
	12305 => "00000000",
	12306 => "00000000",
	12307 => "11111111",
	12308 => "11111111",
	12309 => "11111111",
	12310 => "11111111",
	12311 => "11111111",
	12312 => "11111111",
	12313 => "11111111",
	12314 => "11111111",
	12315 => "11111111",
	12316 => "11111111",
	12317 => "11111111",
	12318 => "00000000",
	12319 => "00000000",
	12320 => "00000000",
	12321 => "00000000",
	12322 => "00000000",
	12323 => "00000000",
	12324 => "00000000",
	12325 => "00000000",
	12326 => "00000000",
	12327 => "00000000",
	12328 => "00000000",
	12329 => "00000000",
	12330 => "00000000",
	12331 => "00000000",
	12332 => "00000000",
	12333 => "00000000",
	12334 => "00000000",
	12335 => "00000000",
	12336 => "00000000",
	12337 => "00000000",
	12338 => "00000000",
	12339 => "00000000",
	12340 => "00000000",
	12341 => "00000000",
	12342 => "00000000",
	12343 => "00000000",
	12344 => "00000000",
	12345 => "00000000",
	12346 => "00000000",
	12347 => "00000000",
	12348 => "00000000",
	12349 => "00000000",
	12350 => "00000000",
	12351 => "00000000",
	12352 => "00000000",
	12353 => "00000000",
	12354 => "00000000",
	12355 => "00000000",
	12356 => "00000000",
	12357 => "00000000",
	12358 => "00000000",
	12359 => "00000000",
	12360 => "00000000",
	12361 => "00000000",
	12362 => "00000000",
	12363 => "00000000",
	12364 => "00000000",
	12365 => "00000000",
	12366 => "00000000",
	12367 => "00000000",
	12368 => "00000000",
	12369 => "00000000",
	12370 => "00000000",
	12371 => "00000000",
	12372 => "00000000",
	12373 => "00000000",
	12374 => "00000000",
	12375 => "00000000",
	12376 => "00000000",
	12377 => "00000000",
	12378 => "00000000",
	12379 => "11111111",
	12380 => "11111111",
	12381 => "11111111",
	12382 => "11111111",
	12383 => "11111111",
	12384 => "11111111",
	12385 => "11111111",
	12386 => "11111111",
	12387 => "11111111",
	12388 => "11111111",
	12389 => "11111111",
	12390 => "00000000",
	12391 => "00000000",
	12392 => "00000000",
	12393 => "00000000",
	12394 => "00000000",
	12395 => "00000000",
	12396 => "00000000",
	12397 => "00000000",
	12398 => "00000000",
	12399 => "00000000",
	12400 => "00000000",
	12401 => "00000000",
	12402 => "00000000",
	12403 => "00000000",
	12404 => "00000000",
	12405 => "00000000",
	12406 => "00000000",
	12407 => "00000000",
	12416 => "00000000",
	12417 => "00000000",
	12418 => "00000000",
	12419 => "00000000",
	12420 => "00000000",
	12421 => "00000000",
	12422 => "00000000",
	12423 => "00000000",
	12424 => "00000000",
	12425 => "00000000",
	12426 => "00000000",
	12427 => "00000000",
	12428 => "00000000",
	12429 => "00000000",
	12430 => "00000000",
	12431 => "00000000",
	12432 => "00000000",
	12433 => "00000000",
	12434 => "11111111",
	12435 => "11111111",
	12436 => "11111111",
	12437 => "11111111",
	12438 => "11111111",
	12439 => "11111111",
	12440 => "11111111",
	12441 => "11111111",
	12442 => "11111111",
	12443 => "11111111",
	12444 => "11111111",
	12445 => "00000000",
	12446 => "00000000",
	12447 => "00000000",
	12448 => "00000000",
	12449 => "00000000",
	12450 => "00000000",
	12451 => "00000000",
	12452 => "00000000",
	12453 => "00000000",
	12454 => "00000000",
	12455 => "00000000",
	12456 => "00000000",
	12457 => "00000000",
	12458 => "00000000",
	12459 => "00000000",
	12460 => "00000000",
	12461 => "00000000",
	12462 => "00000000",
	12463 => "00000000",
	12464 => "00000000",
	12465 => "00000000",
	12466 => "00000000",
	12467 => "00000000",
	12468 => "00000000",
	12469 => "00000000",
	12470 => "00000000",
	12471 => "00000000",
	12472 => "00000000",
	12473 => "00000000",
	12474 => "00000000",
	12475 => "00000000",
	12476 => "00000000",
	12477 => "00000000",
	12478 => "00000000",
	12479 => "00000000",
	12480 => "00000000",
	12481 => "00000000",
	12482 => "00000000",
	12483 => "00000000",
	12484 => "00000000",
	12485 => "00000000",
	12486 => "00000000",
	12487 => "00000000",
	12488 => "00000000",
	12489 => "00000000",
	12490 => "00000000",
	12491 => "00000000",
	12492 => "00000000",
	12493 => "00000000",
	12494 => "00000000",
	12495 => "00000000",
	12496 => "00000000",
	12497 => "00000000",
	12498 => "00000000",
	12499 => "00000000",
	12500 => "00000000",
	12501 => "00000000",
	12502 => "00000000",
	12503 => "00000000",
	12504 => "00000000",
	12505 => "00000000",
	12506 => "00000000",
	12507 => "00000000",
	12508 => "11111111",
	12509 => "11111111",
	12510 => "11111111",
	12511 => "11111111",
	12512 => "11111111",
	12513 => "11111111",
	12514 => "11111111",
	12515 => "11111111",
	12516 => "11111111",
	12517 => "11111111",
	12518 => "11111111",
	12519 => "00000000",
	12520 => "00000000",
	12521 => "00000000",
	12522 => "00000000",
	12523 => "00000000",
	12524 => "00000000",
	12525 => "00000000",
	12526 => "00000000",
	12527 => "00000000",
	12528 => "00000000",
	12529 => "00000000",
	12530 => "00000000",
	12531 => "00000000",
	12532 => "00000000",
	12533 => "00000000",
	12534 => "00000000",
	12535 => "00000000",
	12544 => "00000000",
	12545 => "00000000",
	12546 => "00000000",
	12547 => "00000000",
	12548 => "00000000",
	12549 => "00000000",
	12550 => "00000000",
	12551 => "00000000",
	12552 => "00000000",
	12553 => "00000000",
	12554 => "00000000",
	12555 => "00000000",
	12556 => "00000000",
	12557 => "00000000",
	12558 => "00000000",
	12559 => "00000000",
	12560 => "00000000",
	12561 => "11111111",
	12562 => "11111111",
	12563 => "11111111",
	12564 => "11111111",
	12565 => "11111111",
	12566 => "11111111",
	12567 => "11111111",
	12568 => "11111111",
	12569 => "11111111",
	12570 => "11111111",
	12571 => "11111111",
	12572 => "00000000",
	12573 => "00000000",
	12574 => "00000000",
	12575 => "00000000",
	12576 => "00000000",
	12577 => "00000000",
	12578 => "00000000",
	12579 => "00000000",
	12580 => "00000000",
	12581 => "00000000",
	12582 => "00000000",
	12583 => "00000000",
	12584 => "00000000",
	12585 => "00000000",
	12586 => "00000000",
	12587 => "00000000",
	12588 => "00000000",
	12589 => "00000000",
	12590 => "00000000",
	12591 => "00000000",
	12592 => "00000000",
	12593 => "00000000",
	12594 => "00000000",
	12595 => "00000000",
	12596 => "00000000",
	12597 => "00000000",
	12598 => "00000000",
	12599 => "00000000",
	12600 => "00000000",
	12601 => "00000000",
	12602 => "00000000",
	12603 => "00000000",
	12604 => "00000000",
	12605 => "00000000",
	12606 => "00000000",
	12607 => "00000000",
	12608 => "00000000",
	12609 => "00000000",
	12610 => "00000000",
	12611 => "00000000",
	12612 => "00000000",
	12613 => "00000000",
	12614 => "00000000",
	12615 => "00000000",
	12616 => "00000000",
	12617 => "00000000",
	12618 => "00000000",
	12619 => "00000000",
	12620 => "00000000",
	12621 => "00000000",
	12622 => "00000000",
	12623 => "00000000",
	12624 => "00000000",
	12625 => "00000000",
	12626 => "00000000",
	12627 => "00000000",
	12628 => "00000000",
	12629 => "00000000",
	12630 => "00000000",
	12631 => "00000000",
	12632 => "00000000",
	12633 => "00000000",
	12634 => "00000000",
	12635 => "00000000",
	12636 => "00000000",
	12637 => "11111111",
	12638 => "11111111",
	12639 => "11111111",
	12640 => "11111111",
	12641 => "11111111",
	12642 => "11111111",
	12643 => "11111111",
	12644 => "11111111",
	12645 => "11111111",
	12646 => "11111111",
	12647 => "11111111",
	12648 => "00000000",
	12649 => "00000000",
	12650 => "00000000",
	12651 => "00000000",
	12652 => "00000000",
	12653 => "00000000",
	12654 => "00000000",
	12655 => "00000000",
	12656 => "00000000",
	12657 => "00000000",
	12658 => "00000000",
	12659 => "00000000",
	12660 => "00000000",
	12661 => "00000000",
	12662 => "00000000",
	12663 => "00000000",
	12672 => "00000000",
	12673 => "00000000",
	12674 => "00000000",
	12675 => "00000000",
	12676 => "00000000",
	12677 => "00000000",
	12678 => "00000000",
	12679 => "00000000",
	12680 => "00000000",
	12681 => "00000000",
	12682 => "00000000",
	12683 => "00000000",
	12684 => "00000000",
	12685 => "00000000",
	12686 => "00000000",
	12687 => "00000000",
	12688 => "00000000",
	12689 => "11111111",
	12690 => "11111111",
	12691 => "11111111",
	12692 => "11111111",
	12693 => "11111111",
	12694 => "11111111",
	12695 => "11111111",
	12696 => "11111111",
	12697 => "11111111",
	12698 => "11111111",
	12699 => "00000000",
	12700 => "00000000",
	12701 => "00000000",
	12702 => "00000000",
	12703 => "00000000",
	12704 => "00000000",
	12705 => "00000000",
	12706 => "00000000",
	12707 => "00000000",
	12708 => "00000000",
	12709 => "00000000",
	12710 => "00000000",
	12711 => "00000000",
	12712 => "00000000",
	12713 => "00000000",
	12714 => "00000000",
	12715 => "00000000",
	12716 => "00000000",
	12717 => "00000000",
	12718 => "00000000",
	12719 => "00000000",
	12720 => "00000000",
	12721 => "00000000",
	12722 => "00000000",
	12723 => "00000000",
	12724 => "00000000",
	12725 => "00000000",
	12726 => "00000000",
	12727 => "00000000",
	12728 => "00000000",
	12729 => "00000000",
	12730 => "00000000",
	12731 => "00000000",
	12732 => "00000000",
	12733 => "00000000",
	12734 => "00000000",
	12735 => "00000000",
	12736 => "00000000",
	12737 => "00000000",
	12738 => "00000000",
	12739 => "00000000",
	12740 => "00000000",
	12741 => "00000000",
	12742 => "00000000",
	12743 => "00000000",
	12744 => "00000000",
	12745 => "00000000",
	12746 => "00000000",
	12747 => "00000000",
	12748 => "00000000",
	12749 => "00000000",
	12750 => "00000000",
	12751 => "00000000",
	12752 => "00000000",
	12753 => "00000000",
	12754 => "00000000",
	12755 => "00000000",
	12756 => "00000000",
	12757 => "00000000",
	12758 => "00000000",
	12759 => "00000000",
	12760 => "00000000",
	12761 => "00000000",
	12762 => "00000000",
	12763 => "00000000",
	12764 => "00000000",
	12765 => "00000000",
	12766 => "11111111",
	12767 => "11111111",
	12768 => "11111111",
	12769 => "11111111",
	12770 => "11111111",
	12771 => "11111111",
	12772 => "11111111",
	12773 => "11111111",
	12774 => "11111111",
	12775 => "11111111",
	12776 => "00000000",
	12777 => "00000000",
	12778 => "00000000",
	12779 => "00000000",
	12780 => "00000000",
	12781 => "00000000",
	12782 => "00000000",
	12783 => "00000000",
	12784 => "00000000",
	12785 => "00000000",
	12786 => "00000000",
	12787 => "00000000",
	12788 => "00000000",
	12789 => "00000000",
	12790 => "00000000",
	12791 => "00000000",
	12800 => "00000000",
	12801 => "00000000",
	12802 => "00000000",
	12803 => "00000000",
	12804 => "00000000",
	12805 => "00000000",
	12806 => "00000000",
	12807 => "00000000",
	12808 => "00000000",
	12809 => "00000000",
	12810 => "00000000",
	12811 => "00000000",
	12812 => "00000000",
	12813 => "00000000",
	12814 => "00000000",
	12815 => "00000000",
	12816 => "00000000",
	12817 => "11111111",
	12818 => "11111111",
	12819 => "11111111",
	12820 => "11111111",
	12821 => "11111111",
	12822 => "11111111",
	12823 => "11111111",
	12824 => "11111111",
	12825 => "11111111",
	12826 => "00000000",
	12827 => "00000000",
	12828 => "00000000",
	12829 => "00000000",
	12830 => "00000000",
	12831 => "00000000",
	12832 => "00000000",
	12833 => "00000000",
	12834 => "00000000",
	12835 => "00000000",
	12836 => "00000000",
	12837 => "00000000",
	12838 => "00000000",
	12839 => "00000000",
	12840 => "00000000",
	12841 => "00000000",
	12842 => "00000000",
	12843 => "00000000",
	12844 => "00000000",
	12845 => "00000000",
	12846 => "00000000",
	12847 => "00000000",
	12848 => "00000000",
	12849 => "00000000",
	12850 => "00000000",
	12851 => "00000000",
	12852 => "00000000",
	12853 => "00000000",
	12854 => "00000000",
	12855 => "00000000",
	12856 => "00000000",
	12857 => "00000000",
	12858 => "00000000",
	12859 => "00000000",
	12860 => "00000000",
	12861 => "00000000",
	12862 => "00000000",
	12863 => "00000000",
	12864 => "00000000",
	12865 => "00000000",
	12866 => "00000000",
	12867 => "00000000",
	12868 => "00000000",
	12869 => "00000000",
	12870 => "00000000",
	12871 => "00000000",
	12872 => "00000000",
	12873 => "00000000",
	12874 => "00000000",
	12875 => "00000000",
	12876 => "00000000",
	12877 => "00000000",
	12878 => "00000000",
	12879 => "00000000",
	12880 => "00000000",
	12881 => "00000000",
	12882 => "00000000",
	12883 => "00000000",
	12884 => "00000000",
	12885 => "00000000",
	12886 => "00000000",
	12887 => "00000000",
	12888 => "00000000",
	12889 => "00000000",
	12890 => "00000000",
	12891 => "00000000",
	12892 => "00000000",
	12893 => "00000000",
	12894 => "00000000",
	12895 => "11111111",
	12896 => "11111111",
	12897 => "11111111",
	12898 => "11111111",
	12899 => "11111111",
	12900 => "11111111",
	12901 => "11111111",
	12902 => "11111111",
	12903 => "11111111",
	12904 => "11111111",
	12905 => "00000000",
	12906 => "00000000",
	12907 => "00000000",
	12908 => "00000000",
	12909 => "00000000",
	12910 => "00000000",
	12911 => "00000000",
	12912 => "00000000",
	12913 => "00000000",
	12914 => "00000000",
	12915 => "00000000",
	12916 => "00000000",
	12917 => "00000000",
	12918 => "00000000",
	12919 => "00000000",
	12928 => "00000000",
	12929 => "00000000",
	12930 => "00000000",
	12931 => "00000000",
	12932 => "00000000",
	12933 => "00000000",
	12934 => "00000000",
	12935 => "00000000",
	12936 => "00000000",
	12937 => "00000000",
	12938 => "00000000",
	12939 => "00000000",
	12940 => "00000000",
	12941 => "00000000",
	12942 => "00000000",
	12943 => "00000000",
	12944 => "00000000",
	12945 => "11111111",
	12946 => "11111111",
	12947 => "11111111",
	12948 => "11111111",
	12949 => "11111111",
	12950 => "11111111",
	12951 => "11111111",
	12952 => "11111111",
	12953 => "00000000",
	12954 => "00000000",
	12955 => "00000000",
	12956 => "00000000",
	12957 => "00000000",
	12958 => "00000000",
	12959 => "00000000",
	12960 => "00000000",
	12961 => "00000000",
	12962 => "00000000",
	12963 => "00000000",
	12964 => "00000000",
	12965 => "00000000",
	12966 => "00000000",
	12967 => "00000000",
	12968 => "00000000",
	12969 => "00000000",
	12970 => "00000000",
	12971 => "00000000",
	12972 => "00000000",
	12973 => "00000000",
	12974 => "00000000",
	12975 => "00000000",
	12976 => "00000000",
	12977 => "00000000",
	12978 => "00000000",
	12979 => "00000000",
	12980 => "00000000",
	12981 => "00000000",
	12982 => "00000000",
	12983 => "00000000",
	12984 => "00000000",
	12985 => "00000000",
	12986 => "00000000",
	12987 => "00000000",
	12988 => "00000000",
	12989 => "00000000",
	12990 => "00000000",
	12991 => "00000000",
	12992 => "00000000",
	12993 => "00000000",
	12994 => "00000000",
	12995 => "00000000",
	12996 => "00000000",
	12997 => "00000000",
	12998 => "00000000",
	12999 => "00000000",
	13000 => "00000000",
	13001 => "00000000",
	13002 => "00000000",
	13003 => "00000000",
	13004 => "00000000",
	13005 => "00000000",
	13006 => "00000000",
	13007 => "00000000",
	13008 => "00000000",
	13009 => "00000000",
	13010 => "00000000",
	13011 => "00000000",
	13012 => "00000000",
	13013 => "00000000",
	13014 => "00000000",
	13015 => "00000000",
	13016 => "00000000",
	13017 => "00000000",
	13018 => "00000000",
	13019 => "00000000",
	13020 => "00000000",
	13021 => "00000000",
	13022 => "00000000",
	13023 => "00000000",
	13024 => "11111111",
	13025 => "11111111",
	13026 => "11111111",
	13027 => "11111111",
	13028 => "11111111",
	13029 => "11111111",
	13030 => "11111111",
	13031 => "11111111",
	13032 => "00000000",
	13033 => "00000000",
	13034 => "00000000",
	13035 => "00000000",
	13036 => "00000000",
	13037 => "00000000",
	13038 => "00000000",
	13039 => "00000000",
	13040 => "00000000",
	13041 => "00000000",
	13042 => "00000000",
	13043 => "00000000",
	13044 => "00000000",
	13045 => "00000000",
	13046 => "00000000",
	13047 => "00000000",
	13056 => "00000000",
	13057 => "00000000",
	13058 => "00000000",
	13059 => "00000000",
	13060 => "00000000",
	13061 => "00000000",
	13062 => "00000000",
	13063 => "00000000",
	13064 => "00000000",
	13065 => "00000000",
	13066 => "00000000",
	13067 => "00000000",
	13068 => "00000000",
	13069 => "00000000",
	13070 => "00000000",
	13071 => "00000000",
	13072 => "00000000",
	13073 => "11111111",
	13074 => "11111111",
	13075 => "11111111",
	13076 => "11111111",
	13077 => "11111111",
	13078 => "11111111",
	13079 => "11111111",
	13080 => "00000000",
	13081 => "00000000",
	13082 => "00000000",
	13083 => "00000000",
	13084 => "00000000",
	13085 => "00000000",
	13086 => "00000000",
	13087 => "00000000",
	13088 => "00000000",
	13089 => "00000000",
	13090 => "00000000",
	13091 => "00000000",
	13092 => "00000000",
	13093 => "00000000",
	13094 => "00000000",
	13095 => "00000000",
	13096 => "00000000",
	13097 => "00000000",
	13098 => "00000000",
	13099 => "00000000",
	13100 => "00000000",
	13101 => "00000000",
	13102 => "00000000",
	13103 => "00000000",
	13104 => "00000000",
	13105 => "00000000",
	13106 => "00000000",
	13107 => "00000000",
	13108 => "00000000",
	13109 => "00000000",
	13110 => "00000000",
	13111 => "00000000",
	13112 => "00000000",
	13113 => "00000000",
	13114 => "00000000",
	13115 => "00000000",
	13116 => "00000000",
	13117 => "00000000",
	13118 => "00000000",
	13119 => "00000000",
	13120 => "00000000",
	13121 => "00000000",
	13122 => "00000000",
	13123 => "00000000",
	13124 => "00000000",
	13125 => "00000000",
	13126 => "00000000",
	13127 => "00000000",
	13128 => "00000000",
	13129 => "00000000",
	13130 => "00000000",
	13131 => "00000000",
	13132 => "00000000",
	13133 => "00000000",
	13134 => "00000000",
	13135 => "00000000",
	13136 => "00000000",
	13137 => "00000000",
	13138 => "00000000",
	13139 => "00000000",
	13140 => "00000000",
	13141 => "00000000",
	13142 => "00000000",
	13143 => "00000000",
	13144 => "00000000",
	13145 => "00000000",
	13146 => "00000000",
	13147 => "00000000",
	13148 => "00000000",
	13149 => "00000000",
	13150 => "00000000",
	13151 => "00000000",
	13152 => "00000000",
	13153 => "11111111",
	13154 => "11111111",
	13155 => "11111111",
	13156 => "11111111",
	13157 => "11111111",
	13158 => "11111111",
	13159 => "11111111",
	13160 => "00000000",
	13161 => "00000000",
	13162 => "00000000",
	13163 => "00000000",
	13164 => "00000000",
	13165 => "00000000",
	13166 => "00000000",
	13167 => "00000000",
	13168 => "00000000",
	13169 => "00000000",
	13170 => "00000000",
	13171 => "00000000",
	13172 => "00000000",
	13173 => "00000000",
	13174 => "00000000",
	13175 => "00000000",
	13184 => "00000000",
	13185 => "00000000",
	13186 => "00000000",
	13187 => "00000000",
	13188 => "00000000",
	13189 => "00000000",
	13190 => "00000000",
	13191 => "00000000",
	13192 => "00000000",
	13193 => "00000000",
	13194 => "00000000",
	13195 => "00000000",
	13196 => "00000000",
	13197 => "00000000",
	13198 => "00000000",
	13199 => "00000000",
	13200 => "00000000",
	13201 => "00000000",
	13202 => "11111111",
	13203 => "11111111",
	13204 => "11111111",
	13205 => "11111111",
	13206 => "11111111",
	13207 => "00000000",
	13208 => "00000000",
	13209 => "00000000",
	13210 => "00000000",
	13211 => "00000000",
	13212 => "00000000",
	13213 => "00000000",
	13214 => "00000000",
	13215 => "00000000",
	13216 => "00000000",
	13217 => "00000000",
	13218 => "00000000",
	13219 => "00000000",
	13220 => "00000000",
	13221 => "00000000",
	13222 => "00000000",
	13223 => "00000000",
	13224 => "00000000",
	13225 => "00000000",
	13226 => "00000000",
	13227 => "00000000",
	13228 => "00000000",
	13229 => "00000000",
	13230 => "00000000",
	13231 => "00000000",
	13232 => "00000000",
	13233 => "00000000",
	13234 => "00000000",
	13235 => "00000000",
	13236 => "00000000",
	13237 => "00000000",
	13238 => "00000000",
	13239 => "00000000",
	13240 => "00000000",
	13241 => "00000000",
	13242 => "00000000",
	13243 => "00000000",
	13244 => "00000000",
	13245 => "00000000",
	13246 => "00000000",
	13247 => "00000000",
	13248 => "00000000",
	13249 => "00000000",
	13250 => "00000000",
	13251 => "00000000",
	13252 => "00000000",
	13253 => "00000000",
	13254 => "00000000",
	13255 => "00000000",
	13256 => "00000000",
	13257 => "00000000",
	13258 => "00000000",
	13259 => "00000000",
	13260 => "00000000",
	13261 => "00000000",
	13262 => "00000000",
	13263 => "00000000",
	13264 => "00000000",
	13265 => "00000000",
	13266 => "00000000",
	13267 => "00000000",
	13268 => "00000000",
	13269 => "00000000",
	13270 => "00000000",
	13271 => "00000000",
	13272 => "00000000",
	13273 => "00000000",
	13274 => "00000000",
	13275 => "00000000",
	13276 => "00000000",
	13277 => "00000000",
	13278 => "00000000",
	13279 => "00000000",
	13280 => "00000000",
	13281 => "00000000",
	13282 => "11111111",
	13283 => "11111111",
	13284 => "11111111",
	13285 => "11111111",
	13286 => "11111111",
	13287 => "00000000",
	13288 => "00000000",
	13289 => "00000000",
	13290 => "00000000",
	13291 => "00000000",
	13292 => "00000000",
	13293 => "00000000",
	13294 => "00000000",
	13295 => "00000000",
	13296 => "00000000",
	13297 => "00000000",
	13298 => "00000000",
	13299 => "00000000",
	13300 => "00000000",
	13301 => "00000000",
	13302 => "00000000",
	13303 => "00000000",
	13312 => "00000000",
	13313 => "00000000",
	13314 => "00000000",
	13315 => "00000000",
	13316 => "00000000",
	13317 => "00000000",
	13318 => "00000000",
	13319 => "00000000",
	13320 => "00000000",
	13321 => "00000000",
	13322 => "00000000",
	13323 => "00000000",
	13324 => "00000000",
	13325 => "00000000",
	13326 => "00000000",
	13327 => "00000000",
	13328 => "00000000",
	13329 => "00000000",
	13330 => "00000000",
	13331 => "00000000",
	13332 => "11111111",
	13333 => "00000000",
	13334 => "00000000",
	13335 => "00000000",
	13336 => "00000000",
	13337 => "00000000",
	13338 => "00000000",
	13339 => "00000000",
	13340 => "00000000",
	13341 => "00000000",
	13342 => "00000000",
	13343 => "00000000",
	13344 => "00000000",
	13345 => "00000000",
	13346 => "00000000",
	13347 => "00000000",
	13348 => "00000000",
	13349 => "00000000",
	13350 => "00000000",
	13351 => "00000000",
	13352 => "00000000",
	13353 => "00000000",
	13354 => "00000000",
	13355 => "00000000",
	13356 => "00000000",
	13357 => "00000000",
	13358 => "00000000",
	13359 => "00000000",
	13360 => "00000000",
	13361 => "00000000",
	13362 => "00000000",
	13363 => "00000000",
	13364 => "00000000",
	13365 => "00000000",
	13366 => "00000000",
	13367 => "00000000",
	13368 => "00000000",
	13369 => "00000000",
	13370 => "00000000",
	13371 => "00000000",
	13372 => "00000000",
	13373 => "00000000",
	13374 => "00000000",
	13375 => "00000000",
	13376 => "00000000",
	13377 => "00000000",
	13378 => "00000000",
	13379 => "00000000",
	13380 => "00000000",
	13381 => "00000000",
	13382 => "00000000",
	13383 => "00000000",
	13384 => "00000000",
	13385 => "00000000",
	13386 => "00000000",
	13387 => "00000000",
	13388 => "00000000",
	13389 => "00000000",
	13390 => "00000000",
	13391 => "00000000",
	13392 => "00000000",
	13393 => "00000000",
	13394 => "00000000",
	13395 => "00000000",
	13396 => "00000000",
	13397 => "00000000",
	13398 => "00000000",
	13399 => "00000000",
	13400 => "00000000",
	13401 => "00000000",
	13402 => "00000000",
	13403 => "00000000",
	13404 => "00000000",
	13405 => "00000000",
	13406 => "00000000",
	13407 => "00000000",
	13408 => "00000000",
	13409 => "00000000",
	13410 => "00000000",
	13411 => "00000000",
	13412 => "11111111",
	13413 => "00000000",
	13414 => "00000000",
	13415 => "00000000",
	13416 => "00000000",
	13417 => "00000000",
	13418 => "00000000",
	13419 => "00000000",
	13420 => "00000000",
	13421 => "00000000",
	13422 => "00000000",
	13423 => "00000000",
	13424 => "00000000",
	13425 => "00000000",
	13426 => "00000000",
	13427 => "00000000",
	13428 => "00000000",
	13429 => "00000000",
	13430 => "00000000",
	13431 => "00000000",
	13440 => "00000000",
	13441 => "00000000",
	13442 => "00000000",
	13443 => "00000000",
	13444 => "00000000",
	13445 => "00000000",
	13446 => "00000000",
	13447 => "00000000",
	13448 => "00000000",
	13449 => "00000000",
	13450 => "00000000",
	13451 => "00000000",
	13452 => "00000000",
	13453 => "00000000",
	13454 => "00000000",
	13455 => "00000000",
	13456 => "00000000",
	13457 => "00000000",
	13458 => "00000000",
	13459 => "00000000",
	13460 => "00000000",
	13461 => "00000000",
	13462 => "00000000",
	13463 => "00000000",
	13464 => "00000000",
	13465 => "00000000",
	13466 => "00000000",
	13467 => "00000000",
	13468 => "00000000",
	13469 => "00000000",
	13470 => "00000000",
	13471 => "00000000",
	13472 => "00000000",
	13473 => "00000000",
	13474 => "00000000",
	13475 => "00000000",
	13476 => "00000000",
	13477 => "00000000",
	13478 => "00000000",
	13479 => "00000000",
	13480 => "00000000",
	13481 => "00000000",
	13482 => "00000000",
	13483 => "00000000",
	13484 => "00000000",
	13485 => "00000000",
	13486 => "00000000",
	13487 => "00000000",
	13488 => "00000000",
	13489 => "00000000",
	13490 => "00000000",
	13491 => "00000000",
	13492 => "00000000",
	13493 => "00000000",
	13494 => "00000000",
	13495 => "00000000",
	13496 => "00000000",
	13497 => "00000000",
	13498 => "00000000",
	13499 => "00000000",
	13500 => "00000000",
	13501 => "00000000",
	13502 => "00000000",
	13503 => "00000000",
	13504 => "00000000",
	13505 => "00000000",
	13506 => "00000000",
	13507 => "00000000",
	13508 => "00000000",
	13509 => "00000000",
	13510 => "00000000",
	13511 => "00000000",
	13512 => "00000000",
	13513 => "00000000",
	13514 => "00000000",
	13515 => "00000000",
	13516 => "00000000",
	13517 => "00000000",
	13518 => "00000000",
	13519 => "00000000",
	13520 => "00000000",
	13521 => "00000000",
	13522 => "00000000",
	13523 => "00000000",
	13524 => "00000000",
	13525 => "00000000",
	13526 => "00000000",
	13527 => "00000000",
	13528 => "00000000",
	13529 => "00000000",
	13530 => "00000000",
	13531 => "00000000",
	13532 => "00000000",
	13533 => "00000000",
	13534 => "00000000",
	13535 => "00000000",
	13536 => "00000000",
	13537 => "00000000",
	13538 => "00000000",
	13539 => "00000000",
	13540 => "00000000",
	13541 => "00000000",
	13542 => "00000000",
	13543 => "00000000",
	13544 => "00000000",
	13545 => "00000000",
	13546 => "00000000",
	13547 => "00000000",
	13548 => "00000000",
	13549 => "00000000",
	13550 => "00000000",
	13551 => "00000000",
	13552 => "00000000",
	13553 => "00000000",
	13554 => "00000000",
	13555 => "00000000",
	13556 => "00000000",
	13557 => "00000000",
	13558 => "00000000",
	13559 => "00000000",
	13568 => "00000000",
	13569 => "00000000",
	13570 => "00000000",
	13571 => "00000000",
	13572 => "00000000",
	13573 => "00000000",
	13574 => "00000000",
	13575 => "00000000",
	13576 => "00000000",
	13577 => "00000000",
	13578 => "00000000",
	13579 => "00000000",
	13580 => "00000000",
	13581 => "00000000",
	13582 => "00000000",
	13583 => "00000000",
	13584 => "00000000",
	13585 => "00000000",
	13586 => "00000000",
	13587 => "00000000",
	13588 => "00000000",
	13589 => "00000000",
	13590 => "00000000",
	13591 => "00000000",
	13592 => "00000000",
	13593 => "00000000",
	13594 => "00000000",
	13595 => "00000000",
	13596 => "00000000",
	13597 => "00000000",
	13598 => "00000000",
	13599 => "00000000",
	13600 => "00000000",
	13601 => "00000000",
	13602 => "00000000",
	13603 => "00000000",
	13604 => "00000000",
	13605 => "00000000",
	13606 => "00000000",
	13607 => "00000000",
	13608 => "00000000",
	13609 => "00000000",
	13610 => "00000000",
	13611 => "00000000",
	13612 => "00000000",
	13613 => "00000000",
	13614 => "00000000",
	13615 => "00000000",
	13616 => "00000000",
	13617 => "00000000",
	13618 => "00000000",
	13619 => "00000000",
	13620 => "00000000",
	13621 => "00000000",
	13622 => "00000000",
	13623 => "00000000",
	13624 => "00000000",
	13625 => "00000000",
	13626 => "00000000",
	13627 => "00000000",
	13628 => "00000000",
	13629 => "00000000",
	13630 => "00000000",
	13631 => "00000000",
	13632 => "00000000",
	13633 => "00000000",
	13634 => "00000000",
	13635 => "00000000",
	13636 => "00000000",
	13637 => "00000000",
	13638 => "00000000",
	13639 => "00000000",
	13640 => "00000000",
	13641 => "00000000",
	13642 => "00000000",
	13643 => "00000000",
	13644 => "00000000",
	13645 => "00000000",
	13646 => "00000000",
	13647 => "00000000",
	13648 => "00000000",
	13649 => "00000000",
	13650 => "00000000",
	13651 => "00000000",
	13652 => "00000000",
	13653 => "00000000",
	13654 => "00000000",
	13655 => "00000000",
	13656 => "00000000",
	13657 => "00000000",
	13658 => "00000000",
	13659 => "00000000",
	13660 => "00000000",
	13661 => "00000000",
	13662 => "00000000",
	13663 => "00000000",
	13664 => "00000000",
	13665 => "00000000",
	13666 => "00000000",
	13667 => "00000000",
	13668 => "00000000",
	13669 => "00000000",
	13670 => "00000000",
	13671 => "00000000",
	13672 => "00000000",
	13673 => "00000000",
	13674 => "00000000",
	13675 => "00000000",
	13676 => "00000000",
	13677 => "00000000",
	13678 => "00000000",
	13679 => "00000000",
	13680 => "00000000",
	13681 => "00000000",
	13682 => "00000000",
	13683 => "00000000",
	13684 => "00000000",
	13685 => "00000000",
	13686 => "00000000",
	13687 => "00000000",
	13696 => "00000000",
	13697 => "00000000",
	13698 => "00000000",
	13699 => "00000000",
	13700 => "00000000",
	13701 => "00000000",
	13702 => "00000000",
	13703 => "00000000",
	13704 => "00000000",
	13705 => "00000000",
	13706 => "00000000",
	13707 => "00000000",
	13708 => "00000000",
	13709 => "00000000",
	13710 => "00000000",
	13711 => "00000000",
	13712 => "00000000",
	13713 => "00000000",
	13714 => "00000000",
	13715 => "00000000",
	13716 => "00000000",
	13717 => "00000000",
	13718 => "00000000",
	13719 => "00000000",
	13720 => "00000000",
	13721 => "00000000",
	13722 => "00000000",
	13723 => "00000000",
	13724 => "00000000",
	13725 => "00000000",
	13726 => "00000000",
	13727 => "00000000",
	13728 => "00000000",
	13729 => "00000000",
	13730 => "00000000",
	13731 => "00000000",
	13732 => "00000000",
	13733 => "00000000",
	13734 => "00000000",
	13735 => "00000000",
	13736 => "00000000",
	13737 => "00000000",
	13738 => "00000000",
	13739 => "00000000",
	13740 => "00000000",
	13741 => "00000000",
	13742 => "00000000",
	13743 => "00000000",
	13744 => "00000000",
	13745 => "00000000",
	13746 => "00000000",
	13747 => "00000000",
	13748 => "00000000",
	13749 => "00000000",
	13750 => "00000000",
	13751 => "00000000",
	13752 => "00000000",
	13753 => "00000000",
	13754 => "00000000",
	13755 => "00000000",
	13756 => "00000000",
	13757 => "00000000",
	13758 => "00000000",
	13759 => "00000000",
	13760 => "00000000",
	13761 => "00000000",
	13762 => "00000000",
	13763 => "00000000",
	13764 => "00000000",
	13765 => "00000000",
	13766 => "00000000",
	13767 => "00000000",
	13768 => "00000000",
	13769 => "00000000",
	13770 => "00000000",
	13771 => "00000000",
	13772 => "00000000",
	13773 => "00000000",
	13774 => "00000000",
	13775 => "00000000",
	13776 => "00000000",
	13777 => "00000000",
	13778 => "00000000",
	13779 => "00000000",
	13780 => "00000000",
	13781 => "00000000",
	13782 => "00000000",
	13783 => "00000000",
	13784 => "00000000",
	13785 => "00000000",
	13786 => "00000000",
	13787 => "00000000",
	13788 => "00000000",
	13789 => "00000000",
	13790 => "00000000",
	13791 => "00000000",
	13792 => "00000000",
	13793 => "00000000",
	13794 => "00000000",
	13795 => "00000000",
	13796 => "00000000",
	13797 => "00000000",
	13798 => "00000000",
	13799 => "00000000",
	13800 => "00000000",
	13801 => "00000000",
	13802 => "00000000",
	13803 => "00000000",
	13804 => "00000000",
	13805 => "00000000",
	13806 => "00000000",
	13807 => "00000000",
	13808 => "00000000",
	13809 => "00000000",
	13810 => "00000000",
	13811 => "00000000",
	13812 => "00000000",
	13813 => "00000000",
	13814 => "00000000",
	13815 => "00000000",
	13824 => "00000000",
	13825 => "00000000",
	13826 => "00000000",
	13827 => "00000000",
	13828 => "00000000",
	13829 => "00000000",
	13830 => "00000000",
	13831 => "00000000",
	13832 => "00000000",
	13833 => "00000000",
	13834 => "00000000",
	13835 => "00000000",
	13836 => "00000000",
	13837 => "00000000",
	13838 => "00000000",
	13839 => "00000000",
	13840 => "00000000",
	13841 => "00000000",
	13842 => "00000000",
	13843 => "00000000",
	13844 => "00000000",
	13845 => "00000000",
	13846 => "00000000",
	13847 => "00000000",
	13848 => "00000000",
	13849 => "00000000",
	13850 => "00000000",
	13851 => "00000000",
	13852 => "00000000",
	13853 => "00000000",
	13854 => "00000000",
	13855 => "00000000",
	13856 => "00000000",
	13857 => "00000000",
	13858 => "00000000",
	13859 => "00000000",
	13860 => "00000000",
	13861 => "00000000",
	13862 => "00000000",
	13863 => "00000000",
	13864 => "00000000",
	13865 => "00000000",
	13866 => "00000000",
	13867 => "00000000",
	13868 => "00000000",
	13869 => "00000000",
	13870 => "00000000",
	13871 => "00000000",
	13872 => "00000000",
	13873 => "00000000",
	13874 => "00000000",
	13875 => "00000000",
	13876 => "00000000",
	13877 => "00000000",
	13878 => "00000000",
	13879 => "00000000",
	13880 => "00000000",
	13881 => "00000000",
	13882 => "00000000",
	13883 => "00000000",
	13884 => "00000000",
	13885 => "00000000",
	13886 => "00000000",
	13887 => "00000000",
	13888 => "00000000",
	13889 => "00000000",
	13890 => "00000000",
	13891 => "00000000",
	13892 => "00000000",
	13893 => "00000000",
	13894 => "00000000",
	13895 => "00000000",
	13896 => "00000000",
	13897 => "00000000",
	13898 => "00000000",
	13899 => "00000000",
	13900 => "00000000",
	13901 => "00000000",
	13902 => "00000000",
	13903 => "00000000",
	13904 => "00000000",
	13905 => "00000000",
	13906 => "00000000",
	13907 => "00000000",
	13908 => "00000000",
	13909 => "00000000",
	13910 => "00000000",
	13911 => "00000000",
	13912 => "00000000",
	13913 => "00000000",
	13914 => "00000000",
	13915 => "00000000",
	13916 => "00000000",
	13917 => "00000000",
	13918 => "00000000",
	13919 => "00000000",
	13920 => "00000000",
	13921 => "00000000",
	13922 => "00000000",
	13923 => "00000000",
	13924 => "00000000",
	13925 => "00000000",
	13926 => "00000000",
	13927 => "00000000",
	13928 => "00000000",
	13929 => "00000000",
	13930 => "00000000",
	13931 => "00000000",
	13932 => "00000000",
	13933 => "00000000",
	13934 => "00000000",
	13935 => "00000000",
	13936 => "00000000",
	13937 => "00000000",
	13938 => "00000000",
	13939 => "00000000",
	13940 => "00000000",
	13941 => "00000000",
	13942 => "00000000",
	13943 => "00000000",
	13952 => "00000000",
	13953 => "00000000",
	13954 => "00000000",
	13955 => "00000000",
	13956 => "00000000",
	13957 => "00000000",
	13958 => "00000000",
	13959 => "00000000",
	13960 => "00000000",
	13961 => "00000000",
	13962 => "00000000",
	13963 => "00000000",
	13964 => "00000000",
	13965 => "00000000",
	13966 => "00000000",
	13967 => "00000000",
	13968 => "00000000",
	13969 => "00000000",
	13970 => "00000000",
	13971 => "00000000",
	13972 => "00000000",
	13973 => "00000000",
	13974 => "00000000",
	13975 => "00000000",
	13976 => "00000000",
	13977 => "00000000",
	13978 => "00000000",
	13979 => "00000000",
	13980 => "00000000",
	13981 => "00000000",
	13982 => "00000000",
	13983 => "00000000",
	13984 => "00000000",
	13985 => "00000000",
	13986 => "00000000",
	13987 => "00000000",
	13988 => "00000000",
	13989 => "00000000",
	13990 => "00000000",
	13991 => "00000000",
	13992 => "00000000",
	13993 => "00000000",
	13994 => "00000000",
	13995 => "00000000",
	13996 => "00000000",
	13997 => "00000000",
	13998 => "00000000",
	13999 => "00000000",
	14000 => "00000000",
	14001 => "00000000",
	14002 => "00000000",
	14003 => "00000000",
	14004 => "00000000",
	14005 => "00000000",
	14006 => "00000000",
	14007 => "00000000",
	14008 => "00000000",
	14009 => "00000000",
	14010 => "00000000",
	14011 => "00000000",
	14012 => "00000000",
	14013 => "00000000",
	14014 => "00000000",
	14015 => "00000000",
	14016 => "00000000",
	14017 => "00000000",
	14018 => "00000000",
	14019 => "00000000",
	14020 => "00000000",
	14021 => "00000000",
	14022 => "00000000",
	14023 => "00000000",
	14024 => "00000000",
	14025 => "00000000",
	14026 => "00000000",
	14027 => "00000000",
	14028 => "00000000",
	14029 => "00000000",
	14030 => "00000000",
	14031 => "00000000",
	14032 => "00000000",
	14033 => "00000000",
	14034 => "00000000",
	14035 => "00000000",
	14036 => "00000000",
	14037 => "00000000",
	14038 => "00000000",
	14039 => "00000000",
	14040 => "00000000",
	14041 => "00000000",
	14042 => "00000000",
	14043 => "00000000",
	14044 => "00000000",
	14045 => "00000000",
	14046 => "00000000",
	14047 => "00000000",
	14048 => "00000000",
	14049 => "00000000",
	14050 => "00000000",
	14051 => "00000000",
	14052 => "00000000",
	14053 => "00000000",
	14054 => "00000000",
	14055 => "00000000",
	14056 => "00000000",
	14057 => "00000000",
	14058 => "00000000",
	14059 => "00000000",
	14060 => "00000000",
	14061 => "00000000",
	14062 => "00000000",
	14063 => "00000000",
	14064 => "00000000",
	14065 => "00000000",
	14066 => "00000000",
	14067 => "00000000",
	14068 => "00000000",
	14069 => "00000000",
	14070 => "00000000",
	14071 => "00000000",
	14080 => "00000000",
	14081 => "00000000",
	14082 => "00000000",
	14083 => "00000000",
	14084 => "00000000",
	14085 => "00000000",
	14086 => "00000000",
	14087 => "00000000",
	14088 => "00000000",
	14089 => "00000000",
	14090 => "00000000",
	14091 => "00000000",
	14092 => "00000000",
	14093 => "00000000",
	14094 => "00000000",
	14095 => "00000000",
	14096 => "00000000",
	14097 => "00000000",
	14098 => "00000000",
	14099 => "00000000",
	14100 => "00000000",
	14101 => "00000000",
	14102 => "00000000",
	14103 => "00000000",
	14104 => "00000000",
	14105 => "00000000",
	14106 => "00000000",
	14107 => "00000000",
	14108 => "00000000",
	14109 => "00000000",
	14110 => "00000000",
	14111 => "00000000",
	14112 => "00000000",
	14113 => "00000000",
	14114 => "00000000",
	14115 => "00000000",
	14116 => "00000000",
	14117 => "00000000",
	14118 => "00000000",
	14119 => "00000000",
	14120 => "00000000",
	14121 => "00000000",
	14122 => "00000000",
	14123 => "00000000",
	14124 => "00000000",
	14125 => "00000000",
	14126 => "00000000",
	14127 => "00000000",
	14128 => "00000000",
	14129 => "00000000",
	14130 => "00000000",
	14131 => "00000000",
	14132 => "00000000",
	14133 => "00000000",
	14134 => "00000000",
	14135 => "00000000",
	14136 => "00000000",
	14137 => "00000000",
	14138 => "00000000",
	14139 => "00000000",
	14140 => "00000000",
	14141 => "00000000",
	14142 => "00000000",
	14143 => "00000000",
	14144 => "00000000",
	14145 => "00000000",
	14146 => "00000000",
	14147 => "00000000",
	14148 => "00000000",
	14149 => "00000000",
	14150 => "00000000",
	14151 => "00000000",
	14152 => "00000000",
	14153 => "00000000",
	14154 => "00000000",
	14155 => "00000000",
	14156 => "00000000",
	14157 => "00000000",
	14158 => "00000000",
	14159 => "00000000",
	14160 => "00000000",
	14161 => "00000000",
	14162 => "00000000",
	14163 => "00000000",
	14164 => "00000000",
	14165 => "00000000",
	14166 => "00000000",
	14167 => "00000000",
	14168 => "00000000",
	14169 => "00000000",
	14170 => "00000000",
	14171 => "00000000",
	14172 => "00000000",
	14173 => "00000000",
	14174 => "00000000",
	14175 => "00000000",
	14176 => "00000000",
	14177 => "00000000",
	14178 => "00000000",
	14179 => "00000000",
	14180 => "00000000",
	14181 => "00000000",
	14182 => "00000000",
	14183 => "00000000",
	14184 => "00000000",
	14185 => "00000000",
	14186 => "00000000",
	14187 => "00000000",
	14188 => "00000000",
	14189 => "00000000",
	14190 => "00000000",
	14191 => "00000000",
	14192 => "00000000",
	14193 => "00000000",
	14194 => "00000000",
	14195 => "00000000",
	14196 => "00000000",
	14197 => "00000000",
	14198 => "00000000",
	14199 => "00000000",
	14208 => "00000000",
	14209 => "00000000",
	14210 => "00000000",
	14211 => "00000000",
	14212 => "00000000",
	14213 => "00000000",
	14214 => "00000000",
	14215 => "00000000",
	14216 => "00000000",
	14217 => "00000000",
	14218 => "00000000",
	14219 => "00000000",
	14220 => "00000000",
	14221 => "00000000",
	14222 => "00000000",
	14223 => "00000000",
	14224 => "00000000",
	14225 => "00000000",
	14226 => "00000000",
	14227 => "00000000",
	14228 => "00000000",
	14229 => "00000000",
	14230 => "00000000",
	14231 => "00000000",
	14232 => "00000000",
	14233 => "00000000",
	14234 => "00000000",
	14235 => "00000000",
	14236 => "00000000",
	14237 => "00000000",
	14238 => "00000000",
	14239 => "00000000",
	14240 => "00000000",
	14241 => "00000000",
	14242 => "00000000",
	14243 => "00000000",
	14244 => "00000000",
	14245 => "00000000",
	14246 => "00000000",
	14247 => "00000000",
	14248 => "00000000",
	14249 => "00000000",
	14250 => "00000000",
	14251 => "00000000",
	14252 => "00000000",
	14253 => "00000000",
	14254 => "00000000",
	14255 => "00000000",
	14256 => "00000000",
	14257 => "00000000",
	14258 => "00000000",
	14259 => "00000000",
	14260 => "00000000",
	14261 => "00000000",
	14262 => "00000000",
	14263 => "00000000",
	14264 => "00000000",
	14265 => "00000000",
	14266 => "00000000",
	14267 => "00000000",
	14268 => "00000000",
	14269 => "00000000",
	14270 => "00000000",
	14271 => "00000000",
	14272 => "00000000",
	14273 => "00000000",
	14274 => "00000000",
	14275 => "00000000",
	14276 => "00000000",
	14277 => "00000000",
	14278 => "00000000",
	14279 => "00000000",
	14280 => "00000000",
	14281 => "00000000",
	14282 => "00000000",
	14283 => "00000000",
	14284 => "00000000",
	14285 => "00000000",
	14286 => "00000000",
	14287 => "00000000",
	14288 => "00000000",
	14289 => "00000000",
	14290 => "00000000",
	14291 => "00000000",
	14292 => "00000000",
	14293 => "00000000",
	14294 => "00000000",
	14295 => "00000000",
	14296 => "00000000",
	14297 => "00000000",
	14298 => "00000000",
	14299 => "00000000",
	14300 => "00000000",
	14301 => "00000000",
	14302 => "00000000",
	14303 => "00000000",
	14304 => "00000000",
	14305 => "00000000",
	14306 => "00000000",
	14307 => "00000000",
	14308 => "00000000",
	14309 => "00000000",
	14310 => "00000000",
	14311 => "00000000",
	14312 => "00000000",
	14313 => "00000000",
	14314 => "00000000",
	14315 => "00000000",
	14316 => "00000000",
	14317 => "00000000",
	14318 => "00000000",
	14319 => "00000000",
	14320 => "00000000",
	14321 => "00000000",
	14322 => "00000000",
	14323 => "00000000",
	14324 => "00000000",
	14325 => "00000000",
	14326 => "00000000",
	14327 => "00000000",
	14336 => "00000000",
	14337 => "00000000",
	14338 => "00000000",
	14339 => "00000000",
	14340 => "00000000",
	14341 => "00000000",
	14342 => "00000000",
	14343 => "00000000",
	14344 => "00000000",
	14345 => "00000000",
	14346 => "00000000",
	14347 => "00000000",
	14348 => "00000000",
	14349 => "00000000",
	14350 => "00000000",
	14351 => "00000000",
	14352 => "00000000",
	14353 => "00000000",
	14354 => "00000000",
	14355 => "00000000",
	14356 => "00000000",
	14357 => "00000000",
	14358 => "00000000",
	14359 => "00000000",
	14360 => "00000000",
	14361 => "00000000",
	14362 => "00000000",
	14363 => "00000000",
	14364 => "00000000",
	14365 => "00000000",
	14366 => "00000000",
	14367 => "00000000",
	14368 => "00000000",
	14369 => "00000000",
	14370 => "00000000",
	14371 => "00000000",
	14372 => "00000000",
	14373 => "00000000",
	14374 => "00000000",
	14375 => "00000000",
	14376 => "00000000",
	14377 => "00000000",
	14378 => "00000000",
	14379 => "00000000",
	14380 => "00000000",
	14381 => "00000000",
	14382 => "00000000",
	14383 => "00000000",
	14384 => "00000000",
	14385 => "00000000",
	14386 => "00000000",
	14387 => "00000000",
	14388 => "00000000",
	14389 => "00000000",
	14390 => "00000000",
	14391 => "00000000",
	14392 => "00000000",
	14393 => "00000000",
	14394 => "00000000",
	14395 => "00000000",
	14396 => "00000000",
	14397 => "00000000",
	14398 => "00000000",
	14399 => "00000000",
	14400 => "00000000",
	14401 => "00000000",
	14402 => "00000000",
	14403 => "00000000",
	14404 => "00000000",
	14405 => "00000000",
	14406 => "00000000",
	14407 => "00000000",
	14408 => "00000000",
	14409 => "00000000",
	14410 => "00000000",
	14411 => "00000000",
	14412 => "00000000",
	14413 => "00000000",
	14414 => "00000000",
	14415 => "00000000",
	14416 => "00000000",
	14417 => "00000000",
	14418 => "00000000",
	14419 => "00000000",
	14420 => "00000000",
	14421 => "00000000",
	14422 => "00000000",
	14423 => "00000000",
	14424 => "00000000",
	14425 => "00000000",
	14426 => "00000000",
	14427 => "00000000",
	14428 => "00000000",
	14429 => "00000000",
	14430 => "00000000",
	14431 => "00000000",
	14432 => "00000000",
	14433 => "00000000",
	14434 => "00000000",
	14435 => "00000000",
	14436 => "00000000",
	14437 => "00000000",
	14438 => "00000000",
	14439 => "00000000",
	14440 => "00000000",
	14441 => "00000000",
	14442 => "00000000",
	14443 => "00000000",
	14444 => "00000000",
	14445 => "00000000",
	14446 => "00000000",
	14447 => "00000000",
	14448 => "00000000",
	14449 => "00000000",
	14450 => "00000000",
	14451 => "00000000",
	14452 => "00000000",
	14453 => "00000000",
	14454 => "00000000",
	14455 => "00000000",
	14464 => "00000000",
	14465 => "00000000",
	14466 => "00000000",
	14467 => "00000000",
	14468 => "00000000",
	14469 => "00000000",
	14470 => "00000000",
	14471 => "00000000",
	14472 => "00000000",
	14473 => "00000000",
	14474 => "00000000",
	14475 => "00000000",
	14476 => "00000000",
	14477 => "00000000",
	14478 => "00000000",
	14479 => "00000000",
	14480 => "00000000",
	14481 => "00000000",
	14482 => "00000000",
	14483 => "00000000",
	14484 => "00000000",
	14485 => "00000000",
	14486 => "00000000",
	14487 => "00000000",
	14488 => "00000000",
	14489 => "00000000",
	14490 => "00000000",
	14491 => "00000000",
	14492 => "00000000",
	14493 => "00000000",
	14494 => "00000000",
	14495 => "00000000",
	14496 => "00000000",
	14497 => "00000000",
	14498 => "00000000",
	14499 => "00000000",
	14500 => "00000000",
	14501 => "00000000",
	14502 => "00000000",
	14503 => "00000000",
	14504 => "00000000",
	14505 => "00000000",
	14506 => "00000000",
	14507 => "00000000",
	14508 => "00000000",
	14509 => "00000000",
	14510 => "00000000",
	14511 => "00000000",
	14512 => "00000000",
	14513 => "00000000",
	14514 => "00000000",
	14515 => "00000000",
	14516 => "00000000",
	14517 => "00000000",
	14518 => "00000000",
	14519 => "00000000",
	14520 => "00000000",
	14521 => "00000000",
	14522 => "00000000",
	14523 => "00000000",
	14524 => "00000000",
	14525 => "00000000",
	14526 => "00000000",
	14527 => "00000000",
	14528 => "00000000",
	14529 => "00000000",
	14530 => "00000000",
	14531 => "00000000",
	14532 => "00000000",
	14533 => "00000000",
	14534 => "00000000",
	14535 => "00000000",
	14536 => "00000000",
	14537 => "00000000",
	14538 => "00000000",
	14539 => "00000000",
	14540 => "00000000",
	14541 => "00000000",
	14542 => "00000000",
	14543 => "00000000",
	14544 => "00000000",
	14545 => "00000000",
	14546 => "00000000",
	14547 => "00000000",
	14548 => "00000000",
	14549 => "00000000",
	14550 => "00000000",
	14551 => "00000000",
	14552 => "00000000",
	14553 => "00000000",
	14554 => "00000000",
	14555 => "00000000",
	14556 => "00000000",
	14557 => "00000000",
	14558 => "00000000",
	14559 => "00000000",
	14560 => "00000000",
	14561 => "00000000",
	14562 => "00000000",
	14563 => "00000000",
	14564 => "00000000",
	14565 => "00000000",
	14566 => "00000000",
	14567 => "00000000",
	14568 => "00000000",
	14569 => "00000000",
	14570 => "00000000",
	14571 => "00000000",
	14572 => "00000000",
	14573 => "00000000",
	14574 => "00000000",
	14575 => "00000000",
	14576 => "00000000",
	14577 => "00000000",
	14578 => "00000000",
	14579 => "00000000",
	14580 => "00000000",
	14581 => "00000000",
	14582 => "00000000",
	14583 => "00000000",
	14592 => "00000000",
	14593 => "00000000",
	14594 => "00000000",
	14595 => "00000000",
	14596 => "00000000",
	14597 => "00000000",
	14598 => "00000000",
	14599 => "00000000",
	14600 => "00000000",
	14601 => "00000000",
	14602 => "00000000",
	14603 => "00000000",
	14604 => "00000000",
	14605 => "00000000",
	14606 => "00000000",
	14607 => "00000000",
	14608 => "00000000",
	14609 => "00000000",
	14610 => "00000000",
	14611 => "00000000",
	14612 => "00000000",
	14613 => "00000000",
	14614 => "00000000",
	14615 => "00000000",
	14616 => "00000000",
	14617 => "00000000",
	14618 => "00000000",
	14619 => "00000000",
	14620 => "00000000",
	14621 => "00000000",
	14622 => "00000000",
	14623 => "00000000",
	14624 => "00000000",
	14625 => "00000000",
	14626 => "00000000",
	14627 => "00000000",
	14628 => "00000000",
	14629 => "00000000",
	14630 => "00000000",
	14631 => "00000000",
	14632 => "00000000",
	14633 => "00000000",
	14634 => "00000000",
	14635 => "00000000",
	14636 => "00000000",
	14637 => "00000000",
	14638 => "00000000",
	14639 => "00000000",
	14640 => "00000000",
	14641 => "00000000",
	14642 => "00000000",
	14643 => "00000000",
	14644 => "00000000",
	14645 => "00000000",
	14646 => "00000000",
	14647 => "00000000",
	14648 => "00000000",
	14649 => "00000000",
	14650 => "00000000",
	14651 => "00000000",
	14652 => "00000000",
	14653 => "00000000",
	14654 => "00000000",
	14655 => "00000000",
	14656 => "00000000",
	14657 => "00000000",
	14658 => "00000000",
	14659 => "00000000",
	14660 => "00000000",
	14661 => "00000000",
	14662 => "00000000",
	14663 => "00000000",
	14664 => "00000000",
	14665 => "00000000",
	14666 => "00000000",
	14667 => "00000000",
	14668 => "00000000",
	14669 => "00000000",
	14670 => "00000000",
	14671 => "00000000",
	14672 => "00000000",
	14673 => "00000000",
	14674 => "00000000",
	14675 => "00000000",
	14676 => "00000000",
	14677 => "00000000",
	14678 => "00000000",
	14679 => "00000000",
	14680 => "00000000",
	14681 => "00000000",
	14682 => "00000000",
	14683 => "00000000",
	14684 => "00000000",
	14685 => "00000000",
	14686 => "00000000",
	14687 => "00000000",
	14688 => "00000000",
	14689 => "00000000",
	14690 => "00000000",
	14691 => "00000000",
	14692 => "00000000",
	14693 => "00000000",
	14694 => "00000000",
	14695 => "00000000",
	14696 => "00000000",
	14697 => "00000000",
	14698 => "00000000",
	14699 => "00000000",
	14700 => "00000000",
	14701 => "00000000",
	14702 => "00000000",
	14703 => "00000000",
	14704 => "00000000",
	14705 => "00000000",
	14706 => "00000000",
	14707 => "00000000",
	14708 => "00000000",
	14709 => "00000000",
	14710 => "00000000",
	14711 => "00000000",
	14720 => "00000000",
	14721 => "00000000",
	14722 => "00000000",
	14723 => "00000000",
	14724 => "00000000",
	14725 => "00000000",
	14726 => "00000000",
	14727 => "00000000",
	14728 => "00000000",
	14729 => "00000000",
	14730 => "00000000",
	14731 => "00000000",
	14732 => "00000000",
	14733 => "00000000",
	14734 => "00000000",
	14735 => "00000000",
	14736 => "00000000",
	14737 => "00000000",
	14738 => "00000000",
	14739 => "00000000",
	14740 => "00000000",
	14741 => "00000000",
	14742 => "00000000",
	14743 => "00000000",
	14744 => "00000000",
	14745 => "00000000",
	14746 => "00000000",
	14747 => "00000000",
	14748 => "00000000",
	14749 => "00000000",
	14750 => "00000000",
	14751 => "00000000",
	14752 => "00000000",
	14753 => "00000000",
	14754 => "00000000",
	14755 => "00000000",
	14756 => "00000000",
	14757 => "00000000",
	14758 => "00000000",
	14759 => "00000000",
	14760 => "00000000",
	14761 => "00000000",
	14762 => "00000000",
	14763 => "00000000",
	14764 => "00000000",
	14765 => "00000000",
	14766 => "00000000",
	14767 => "00000000",
	14768 => "00000000",
	14769 => "00000000",
	14770 => "00000000",
	14771 => "00000000",
	14772 => "00000000",
	14773 => "00000000",
	14774 => "00000000",
	14775 => "00000000",
	14776 => "00000000",
	14777 => "00000000",
	14778 => "00000000",
	14779 => "00000000",
	14780 => "00000000",
	14781 => "00000000",
	14782 => "00000000",
	14783 => "00000000",
	14784 => "00000000",
	14785 => "00000000",
	14786 => "00000000",
	14787 => "00000000",
	14788 => "00000000",
	14789 => "00000000",
	14790 => "00000000",
	14791 => "00000000",
	14792 => "00000000",
	14793 => "00000000",
	14794 => "00000000",
	14795 => "00000000",
	14796 => "00000000",
	14797 => "00000000",
	14798 => "00000000",
	14799 => "00000000",
	14800 => "00000000",
	14801 => "00000000",
	14802 => "00000000",
	14803 => "00000000",
	14804 => "00000000",
	14805 => "00000000",
	14806 => "00000000",
	14807 => "00000000",
	14808 => "00000000",
	14809 => "00000000",
	14810 => "00000000",
	14811 => "00000000",
	14812 => "00000000",
	14813 => "00000000",
	14814 => "00000000",
	14815 => "00000000",
	14816 => "00000000",
	14817 => "00000000",
	14818 => "00000000",
	14819 => "00000000",
	14820 => "00000000",
	14821 => "00000000",
	14822 => "00000000",
	14823 => "00000000",
	14824 => "00000000",
	14825 => "00000000",
	14826 => "00000000",
	14827 => "00000000",
	14828 => "00000000",
	14829 => "00000000",
	14830 => "00000000",
	14831 => "00000000",
	14832 => "00000000",
	14833 => "00000000",
	14834 => "00000000",
	14835 => "00000000",
	14836 => "00000000",
	14837 => "00000000",
	14838 => "00000000",
	14839 => "00000000",
	14848 => "00000000",
	14849 => "00000000",
	14850 => "00000000",
	14851 => "00000000",
	14852 => "00000000",
	14853 => "00000000",
	14854 => "00000000",
	14855 => "00000000",
	14856 => "00000000",
	14857 => "00000000",
	14858 => "00000000",
	14859 => "00000000",
	14860 => "00000000",
	14861 => "00000000",
	14862 => "00000000",
	14863 => "00000000",
	14864 => "00000000",
	14865 => "00000000",
	14866 => "00000000",
	14867 => "00000000",
	14868 => "00000000",
	14869 => "00000000",
	14870 => "00000000",
	14871 => "00000000",
	14872 => "00000000",
	14873 => "00000000",
	14874 => "00000000",
	14875 => "00000000",
	14876 => "00000000",
	14877 => "00000000",
	14878 => "00000000",
	14879 => "00000000",
	14880 => "00000000",
	14881 => "00000000",
	14882 => "00000000",
	14883 => "00000000",
	14884 => "00000000",
	14885 => "00000000",
	14886 => "00000000",
	14887 => "00000000",
	14888 => "00000000",
	14889 => "00000000",
	14890 => "00000000",
	14891 => "00000000",
	14892 => "00000000",
	14893 => "00000000",
	14894 => "00000000",
	14895 => "00000000",
	14896 => "00000000",
	14897 => "00000000",
	14898 => "00000000",
	14899 => "00000000",
	14900 => "00000000",
	14901 => "00000000",
	14902 => "00000000",
	14903 => "00000000",
	14904 => "00000000",
	14905 => "00000000",
	14906 => "00000000",
	14907 => "00000000",
	14908 => "00000000",
	14909 => "00000000",
	14910 => "00000000",
	14911 => "00000000",
	14912 => "00000000",
	14913 => "00000000",
	14914 => "00000000",
	14915 => "00000000",
	14916 => "00000000",
	14917 => "00000000",
	14918 => "00000000",
	14919 => "00000000",
	14920 => "00000000",
	14921 => "00000000",
	14922 => "00000000",
	14923 => "00000000",
	14924 => "00000000",
	14925 => "00000000",
	14926 => "00000000",
	14927 => "00000000",
	14928 => "00000000",
	14929 => "00000000",
	14930 => "00000000",
	14931 => "00000000",
	14932 => "00000000",
	14933 => "00000000",
	14934 => "00000000",
	14935 => "00000000",
	14936 => "00000000",
	14937 => "00000000",
	14938 => "00000000",
	14939 => "00000000",
	14940 => "00000000",
	14941 => "00000000",
	14942 => "00000000",
	14943 => "00000000",
	14944 => "00000000",
	14945 => "00000000",
	14946 => "00000000",
	14947 => "00000000",
	14948 => "00000000",
	14949 => "00000000",
	14950 => "00000000",
	14951 => "00000000",
	14952 => "00000000",
	14953 => "00000000",
	14954 => "00000000",
	14955 => "00000000",
	14956 => "00000000",
	14957 => "00000000",
	14958 => "00000000",
	14959 => "00000000",
	14960 => "00000000",
	14961 => "00000000",
	14962 => "00000000",
	14963 => "00000000",
	14964 => "00000000",
	14965 => "00000000",
	14966 => "00000000",
	14967 => "00000000",
	14976 => "00000000",
	14977 => "00000000",
	14978 => "00000000",
	14979 => "00000000",
	14980 => "00000000",
	14981 => "00000000",
	14982 => "00000000",
	14983 => "00000000",
	14984 => "00000000",
	14985 => "00000000",
	14986 => "00000000",
	14987 => "00000000",
	14988 => "00000000",
	14989 => "00000000",
	14990 => "00000000",
	14991 => "00000000",
	14992 => "00000000",
	14993 => "00000000",
	14994 => "00000000",
	14995 => "00000000",
	14996 => "00000000",
	14997 => "00000000",
	14998 => "00000000",
	14999 => "00000000",
	15000 => "00000000",
	15001 => "00000000",
	15002 => "00000000",
	15003 => "00000000",
	15004 => "00000000",
	15005 => "00000000",
	15006 => "00000000",
	15007 => "00000000",
	15008 => "00000000",
	15009 => "00000000",
	15010 => "00000000",
	15011 => "00000000",
	15012 => "00000000",
	15013 => "00000000",
	15014 => "00000000",
	15015 => "00000000",
	15016 => "00000000",
	15017 => "00000000",
	15018 => "00000000",
	15019 => "00000000",
	15020 => "00000000",
	15021 => "00000000",
	15022 => "00000000",
	15023 => "00000000",
	15024 => "00000000",
	15025 => "00000000",
	15026 => "00000000",
	15027 => "00000000",
	15028 => "00000000",
	15029 => "00000000",
	15030 => "00000000",
	15031 => "00000000",
	15032 => "00000000",
	15033 => "00000000",
	15034 => "00000000",
	15035 => "00000000",
	15036 => "00000000",
	15037 => "00000000",
	15038 => "00000000",
	15039 => "00000000",
	15040 => "00000000",
	15041 => "00000000",
	15042 => "00000000",
	15043 => "00000000",
	15044 => "00000000",
	15045 => "00000000",
	15046 => "00000000",
	15047 => "00000000",
	15048 => "00000000",
	15049 => "00000000",
	15050 => "00000000",
	15051 => "00000000",
	15052 => "00000000",
	15053 => "00000000",
	15054 => "00000000",
	15055 => "00000000",
	15056 => "00000000",
	15057 => "00000000",
	15058 => "00000000",
	15059 => "00000000",
	15060 => "00000000",
	15061 => "00000000",
	15062 => "00000000",
	15063 => "00000000",
	15064 => "00000000",
	15065 => "00000000",
	15066 => "00000000",
	15067 => "00000000",
	15068 => "00000000",
	15069 => "00000000",
	15070 => "00000000",
	15071 => "00000000",
	15072 => "00000000",
	15073 => "00000000",
	15074 => "00000000",
	15075 => "00000000",
	15076 => "00000000",
	15077 => "00000000",
	15078 => "00000000",
	15079 => "00000000",
	15080 => "00000000",
	15081 => "00000000",
	15082 => "00000000",
	15083 => "00000000",
	15084 => "00000000",
	15085 => "00000000",
	15086 => "00000000",
	15087 => "00000000",
	15088 => "00000000",
	15089 => "00000000",
	15090 => "00000000",
	15091 => "00000000",
	15092 => "00000000",
	15093 => "00000000",
	15094 => "00000000",
	15095 => "00000000",
	15104 => "00000000",
	15105 => "00000000",
	15106 => "00000000",
	15107 => "00000000",
	15108 => "00000000",
	15109 => "00000000",
	15110 => "00000000",
	15111 => "00000000",
	15112 => "00000000",
	15113 => "00000000",
	15114 => "00000000",
	15115 => "00000000",
	15116 => "00000000",
	15117 => "00000000",
	15118 => "00000000",
	15119 => "00000000",
	15120 => "00000000",
	15121 => "00000000",
	15122 => "00000000",
	15123 => "00000000",
	15124 => "00000000",
	15125 => "00000000",
	15126 => "00000000",
	15127 => "00000000",
	15128 => "00000000",
	15129 => "00000000",
	15130 => "00000000",
	15131 => "00000000",
	15132 => "00000000",
	15133 => "00000000",
	15134 => "00000000",
	15135 => "00000000",
	15136 => "00000000",
	15137 => "00000000",
	15138 => "00000000",
	15139 => "00000000",
	15140 => "00000000",
	15141 => "00000000",
	15142 => "00000000",
	15143 => "00000000",
	15144 => "00000000",
	15145 => "00000000",
	15146 => "00000000",
	15147 => "00000000",
	15148 => "00000000",
	15149 => "00000000",
	15150 => "00000000",
	15151 => "00000000",
	15152 => "00000000",
	15153 => "00000000",
	15154 => "00000000",
	15155 => "00000000",
	15156 => "00000000",
	15157 => "00000000",
	15158 => "00000000",
	15159 => "00000000",
	15160 => "00000000",
	15161 => "00000000",
	15162 => "00000000",
	15163 => "00000000",
	15164 => "00000000",
	15165 => "00000000",
	15166 => "00000000",
	15167 => "00000000",
	15168 => "00000000",
	15169 => "00000000",
	15170 => "00000000",
	15171 => "00000000",
	15172 => "00000000",
	15173 => "00000000",
	15174 => "00000000",
	15175 => "00000000",
	15176 => "00000000",
	15177 => "00000000",
	15178 => "00000000",
	15179 => "00000000",
	15180 => "00000000",
	15181 => "00000000",
	15182 => "00000000",
	15183 => "00000000",
	15184 => "00000000",
	15185 => "00000000",
	15186 => "00000000",
	15187 => "00000000",
	15188 => "00000000",
	15189 => "00000000",
	15190 => "00000000",
	15191 => "00000000",
	15192 => "00000000",
	15193 => "00000000",
	15194 => "00000000",
	15195 => "00000000",
	15196 => "00000000",
	15197 => "00000000",
	15198 => "00000000",
	15199 => "00000000",
	15200 => "00000000",
	15201 => "00000000",
	15202 => "00000000",
	15203 => "00000000",
	15204 => "00000000",
	15205 => "00000000",
	15206 => "00000000",
	15207 => "00000000",
	15208 => "00000000",
	15209 => "00000000",
	15210 => "00000000",
	15211 => "00000000",
	15212 => "00000000",
	15213 => "00000000",
	15214 => "00000000",
	15215 => "00000000",
	15216 => "00000000",
	15217 => "00000000",
	15218 => "00000000",
	15219 => "00000000",
	15220 => "00000000",
	15221 => "00000000",
	15222 => "00000000",
	15223 => "00000000",
	15232 => "00000000",
	15233 => "00000000",
	15234 => "00000000",
	15235 => "00000000",
	15236 => "00000000",
	15237 => "00000000",
	15238 => "00000000",
	15239 => "00000000",
	15240 => "00000000",
	15241 => "00000000",
	15242 => "00000000",
	15243 => "00000000",
	15244 => "00000000",
	15245 => "00000000",
	15246 => "00000000",
	15247 => "00000000",
	15248 => "00000000",
	15249 => "00000000",
	15250 => "00000000",
	15251 => "00000000",
	15252 => "00000000",
	15253 => "00000000",
	15254 => "00000000",
	15255 => "00000000",
	15256 => "00000000",
	15257 => "00000000",
	15258 => "00000000",
	15259 => "00000000",
	15260 => "00000000",
	15261 => "00000000",
	15262 => "00000000",
	15263 => "00000000",
	15264 => "00000000",
	15265 => "00000000",
	15266 => "00000000",
	15267 => "00000000",
	15268 => "00000000",
	15269 => "00000000",
	15270 => "00000000",
	15271 => "00000000",
	15272 => "00000000",
	15273 => "00000000",
	15274 => "00000000",
	15275 => "00000000",
	15276 => "00000000",
	15277 => "00000000",
	15278 => "00000000",
	15279 => "00000000",
	15280 => "00000000",
	15281 => "00000000",
	15282 => "00000000",
	15283 => "00000000",
	15284 => "00000000",
	15285 => "00000000",
	15286 => "00000000",
	15287 => "00000000",
	15288 => "00000000",
	15289 => "00000000",
	15290 => "00000000",
	15291 => "00000000",
	15292 => "00000000",
	15293 => "00000000",
	15294 => "00000000",
	15295 => "00000000",
	15296 => "00000000",
	15297 => "00000000",
	15298 => "00000000",
	15299 => "00000000",
	15300 => "00000000",
	15301 => "00000000",
	15302 => "00000000",
	15303 => "00000000",
	15304 => "00000000",
	15305 => "00000000",
	15306 => "00000000",
	15307 => "00000000",
	15308 => "00000000",
	15309 => "00000000",
	15310 => "00000000",
	15311 => "00000000",
	15312 => "00000000",
	15313 => "00000000",
	15314 => "00000000",
	15315 => "00000000",
	15316 => "00000000",
	15317 => "00000000",
	15318 => "00000000",
	15319 => "00000000",
	15320 => "00000000",
	15321 => "00000000",
	15322 => "00000000",
	15323 => "00000000",
	15324 => "00000000",
	15325 => "00000000",
	15326 => "00000000",
	15327 => "00000000",
	15328 => "00000000",
	15329 => "00000000",
	15330 => "00000000",
	15331 => "00000000",
	15332 => "00000000",
	15333 => "00000000",
	15334 => "00000000",
	15335 => "00000000",
	15336 => "00000000",
	15337 => "00000000",
	15338 => "00000000",
	15339 => "00000000",
	15340 => "00000000",
	15341 => "00000000",
	15342 => "00000000",
	15343 => "00000000",
	15344 => "00000000",
	15345 => "00000000",
	15346 => "00000000",
	15347 => "00000000",
	15348 => "00000000",
	15349 => "00000000",
	15350 => "00000000",
	15351 => "00000000",

	others => (others => '0')
);

begin
	
	-- process ROM
	process (CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (EN = '1') then
				DATA <= ROM(conv_integer(ADDR));
			end if;
		end if;
	end process;
	
end Behavioral;

