----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:16:29 04/19/2013 
-- Design Name: 
-- Module Name:    VRAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity VRAM is
	port (Clk		: in 	std_logic;
			CE			: in 	std_logic;
			Enable_w	: in 	std_logic;
			Addr_w	: in 	std_logic_vector	(18 downto 0);
			Addr_r	: in 	std_logic_vector	(18 downto 0);
			Data_in	: in 	std_logic_vector	(7 downto 0);
			Data_out	: out std_logic_vector	(7 downto 0));
end VRAM;

architecture Behavioral of VRAM is
	type ram_type is array ((2**17)-1 downto 0) of std_logic_vector (7 downto 0);
	signal VRAM: ram_type := (
		9225 to 9318 => "11111111",
		10249 to 10249 => "11111111",
		10280 to 10280 => "11111111",
		10311 to 10311 => "11111111",
		10342 to 10342 => "11111111",
		11273 to 11273 => "11111111",
		11304 to 11304 => "11111111",
		11335 to 11335 => "11111111",
		11366 to 11366 => "11111111",
		12297 to 12297 => "11111111",
		12328 to 12328 => "11111111",
		12359 to 12359 => "11111111",
		12390 to 12390 => "11111111",
		13321 to 13321 => "11111111",
		13352 to 13352 => "11111111",
		13383 to 13383 => "11111111",
		13414 to 13414 => "11111111",
		14345 to 14345 => "11111111",
		14376 to 14376 => "11111111",
		14407 to 14407 => "11111111",
		14438 to 14438 => "11111111",
		15369 to 15369 => "11111111",
		15400 to 15400 => "11111111",
		15431 to 15431 => "11111111",
		15462 to 15462 => "11111111",
		16393 to 16393 => "11111111",
		16424 to 16424 => "11111111",
		16455 to 16455 => "11111111",
		16486 to 16486 => "11111111",
		17417 to 17417 => "11111111",
		17448 to 17448 => "11111111",
		17479 to 17479 => "11111111",
		17510 to 17510 => "11111111",
		18441 to 18441 => "11111111",
		18472 to 18472 => "11111111",
		18503 to 18503 => "11111111",
		18534 to 18534 => "11111111",
		19465 to 19465 => "11111111",
		19496 to 19496 => "11111111",
		19527 to 19527 => "11111111",
		19558 to 19558 => "11111111",
		20489 to 20489 => "11111111",
		20520 to 20520 => "11111111",
		20551 to 20551 => "11111111",
		20582 to 20582 => "11111111",
		21513 to 21513 => "11111111",
		21544 to 21544 => "11111111",
		21575 to 21575 => "11111111",
		21606 to 21606 => "11111111",
		22537 to 22537 => "11111111",
		22568 to 22568 => "11111111",
		22599 to 22599 => "11111111",
		22630 to 22630 => "11111111",
		23561 to 23561 => "11111111",
		23592 to 23592 => "11111111",
		23623 to 23623 => "11111111",
		23654 to 23654 => "11111111",
		24585 to 24585 => "11111111",
		24616 to 24616 => "11111111",
		24647 to 24647 => "11111111",
		24678 to 24678 => "11111111",
		25609 to 25609 => "11111111",
		25640 to 25640 => "11111111",
		25671 to 25671 => "11111111",
		25702 to 25702 => "11111111",
		26633 to 26633 => "11111111",
		26664 to 26664 => "11111111",
		26695 to 26695 => "11111111",
		26726 to 26726 => "11111111",
		27657 to 27657 => "11111111",
		27688 to 27688 => "11111111",
		27719 to 27719 => "11111111",
		27750 to 27750 => "11111111",
		28681 to 28681 => "11111111",
		28712 to 28712 => "11111111",
		28743 to 28743 => "11111111",
		28774 to 28774 => "11111111",
		29705 to 29705 => "11111111",
		29736 to 29736 => "11111111",
		29767 to 29767 => "11111111",
		29798 to 29798 => "11111111",
		30729 to 30729 => "11111111",
		30760 to 30760 => "11111111",
		30791 to 30791 => "11111111",
		30822 to 30822 => "11111111",
		31753 to 31753 => "11111111",
		31784 to 31784 => "11111111",
		31815 to 31815 => "11111111",
		31846 to 31846 => "11111111",
		32777 to 32777 => "11111111",
		32808 to 32808 => "11111111",
		32839 to 32839 => "11111111",
		32870 to 32870 => "11111111",
		33801 to 33801 => "11111111",
		33832 to 33832 => "11111111",
		33863 to 33863 => "11111111",
		33894 to 33894 => "11111111",
		34825 to 34825 => "11111111",
		34856 to 34856 => "11111111",
		34887 to 34887 => "11111111",
		34918 to 34918 => "11111111",
		35849 to 35849 => "11111111",
		35880 to 35880 => "11111111",
		35911 to 35911 => "11111111",
		35942 to 35942 => "11111111",
		36873 to 36873 => "11111111",
		36904 to 36904 => "11111111",
		36935 to 36935 => "11111111",
		36966 to 36966 => "11111111",
		37897 to 37897 => "11111111",
		37928 to 37928 => "11111111",
		37959 to 37959 => "11111111",
		37990 to 37990 => "11111111",
		38921 to 38921 => "11111111",
		38952 to 38952 => "11111111",
		38983 to 38983 => "11111111",
		39014 to 39014 => "11111111",
		39945 to 39945 => "11111111",
		39976 to 39976 => "11111111",
		40007 to 40007 => "11111111",
		40038 to 40038 => "11111111",
		40969 to 41062 => "11111111",
		41993 to 41993 => "11111111",
		42024 to 42024 => "11111111",
		42055 to 42055 => "11111111",
		42086 to 42086 => "11111111",
		43017 to 43017 => "11111111",
		43048 to 43048 => "11111111",
		43079 to 43079 => "11111111",
		43110 to 43110 => "11111111",
		44041 to 44041 => "11111111",
		44072 to 44072 => "11111111",
		44103 to 44103 => "11111111",
		44134 to 44134 => "11111111",
		45065 to 45065 => "11111111",
		45096 to 45096 => "11111111",
		45127 to 45127 => "11111111",
		45158 to 45158 => "11111111",
		46089 to 46089 => "11111111",
		46120 to 46120 => "11111111",
		46151 to 46151 => "11111111",
		46182 to 46182 => "11111111",
		47113 to 47113 => "11111111",
		47144 to 47144 => "11111111",
		47175 to 47175 => "11111111",
		47206 to 47206 => "11111111",
		48137 to 48137 => "11111111",
		48168 to 48168 => "11111111",
		48199 to 48199 => "11111111",
		48230 to 48230 => "11111111",
		49161 to 49161 => "11111111",
		49192 to 49192 => "11111111",
		49223 to 49223 => "11111111",
		49254 to 49254 => "11111111",
		50185 to 50185 => "11111111",
		50216 to 50216 => "11111111",
		50247 to 50247 => "11111111",
		50278 to 50278 => "11111111",
		51209 to 51209 => "11111111",
		51240 to 51240 => "11111111",
		51271 to 51271 => "11111111",
		51302 to 51302 => "11111111",
		52233 to 52233 => "11111111",
		52264 to 52264 => "11111111",
		52295 to 52295 => "11111111",
		52326 to 52326 => "11111111",
		53257 to 53257 => "11111111",
		53288 to 53288 => "11111111",
		53319 to 53319 => "11111111",
		53350 to 53350 => "11111111",
		54281 to 54281 => "11111111",
		54312 to 54312 => "11111111",
		54343 to 54343 => "11111111",
		54374 to 54374 => "11111111",
		55305 to 55305 => "11111111",
		55336 to 55336 => "11111111",
		55367 to 55367 => "11111111",
		55398 to 55398 => "11111111",
		56329 to 56329 => "11111111",
		56360 to 56360 => "11111111",
		56391 to 56391 => "11111111",
		56422 to 56422 => "11111111",
		57353 to 57353 => "11111111",
		57384 to 57384 => "11111111",
		57415 to 57415 => "11111111",
		57446 to 57446 => "11111111",
		58377 to 58377 => "11111111",
		58408 to 58408 => "11111111",
		58439 to 58439 => "11111111",
		58470 to 58470 => "11111111",
		59401 to 59401 => "11111111",
		59432 to 59432 => "11111111",
		59463 to 59463 => "11111111",
		59494 to 59494 => "11111111",
		60425 to 60425 => "11111111",
		60456 to 60456 => "11111111",
		60487 to 60487 => "11111111",
		60518 to 60518 => "11111111",
		61449 to 61449 => "11111111",
		61480 to 61480 => "11111111",
		61511 to 61511 => "11111111",
		61542 to 61542 => "11111111",
		62473 to 62473 => "11111111",
		62504 to 62504 => "11111111",
		62535 to 62535 => "11111111",
		62566 to 62566 => "11111111",
		63497 to 63497 => "11111111",
		63528 to 63528 => "11111111",
		63559 to 63559 => "11111111",
		63590 to 63590 => "11111111",
		64521 to 64521 => "11111111",
		64552 to 64552 => "11111111",
		64583 to 64583 => "11111111",
		64614 to 64614 => "11111111",
		65545 to 65545 => "11111111",
		65576 to 65576 => "11111111",
		65607 to 65607 => "11111111",
		65638 to 65638 => "11111111",
		66569 to 66569 => "11111111",
		66600 to 66600 => "11111111",
		66631 to 66631 => "11111111",
		66662 to 66662 => "11111111",
		67593 to 67593 => "11111111",
		67624 to 67624 => "11111111",
		67655 to 67655 => "11111111",
		67686 to 67686 => "11111111",
		68617 to 68617 => "11111111",
		68648 to 68648 => "11111111",
		68679 to 68679 => "11111111",
		68710 to 68710 => "11111111",
		69641 to 69641 => "11111111",
		69672 to 69672 => "11111111",
		69703 to 69703 => "11111111",
		69734 to 69734 => "11111111",
		70665 to 70665 => "11111111",
		70696 to 70696 => "11111111",
		70727 to 70727 => "11111111",
		70758 to 70758 => "11111111",
		71689 to 71689 => "11111111",
		71720 to 71720 => "11111111",
		71751 to 71751 => "11111111",
		71782 to 71782 => "11111111",
		72713 to 72806 => "11111111",
		73737 to 73737 => "11111111",
		73768 to 73768 => "11111111",
		73799 to 73799 => "11111111",
		73830 to 73830 => "11111111",
		74761 to 74761 => "11111111",
		74792 to 74792 => "11111111",
		74823 to 74823 => "11111111",
		74854 to 74854 => "11111111",
		75785 to 75785 => "11111111",
		75816 to 75816 => "11111111",
		75847 to 75847 => "11111111",
		75878 to 75878 => "11111111",
		76809 to 76809 => "11111111",
		76840 to 76840 => "11111111",
		76871 to 76871 => "11111111",
		76902 to 76902 => "11111111",
		77833 to 77833 => "11111111",
		77864 to 77864 => "11111111",
		77895 to 77895 => "11111111",
		77926 to 77926 => "11111111",
		78857 to 78857 => "11111111",
		78888 to 78888 => "11111111",
		78919 to 78919 => "11111111",
		78950 to 78950 => "11111111",
		79881 to 79881 => "11111111",
		79912 to 79912 => "11111111",
		79943 to 79943 => "11111111",
		79974 to 79974 => "11111111",
		80905 to 80905 => "11111111",
		80936 to 80936 => "11111111",
		80967 to 80967 => "11111111",
		80998 to 80998 => "11111111",
		81929 to 81929 => "11111111",
		81960 to 81960 => "11111111",
		81991 to 81991 => "11111111",
		82022 to 82022 => "11111111",
		82953 to 82953 => "11111111",
		82984 to 82984 => "11111111",
		83015 to 83015 => "11111111",
		83046 to 83046 => "11111111",
		83977 to 83977 => "11111111",
		84008 to 84008 => "11111111",
		84039 to 84039 => "11111111",
		84070 to 84070 => "11111111",
		85001 to 85001 => "11111111",
		85032 to 85032 => "11111111",
		85063 to 85063 => "11111111",
		85094 to 85094 => "11111111",
		86025 to 86025 => "11111111",
		86056 to 86056 => "11111111",
		86087 to 86087 => "11111111",
		86118 to 86118 => "11111111",
		87049 to 87049 => "11111111",
		87080 to 87080 => "11111111",
		87111 to 87111 => "11111111",
		87142 to 87142 => "11111111",
		88073 to 88073 => "11111111",
		88104 to 88104 => "11111111",
		88135 to 88135 => "11111111",
		88166 to 88166 => "11111111",
		89097 to 89097 => "11111111",
		89128 to 89128 => "11111111",
		89159 to 89159 => "11111111",
		89190 to 89190 => "11111111",
		90121 to 90121 => "11111111",
		90152 to 90152 => "11111111",
		90183 to 90183 => "11111111",
		90214 to 90214 => "11111111",
		91145 to 91145 => "11111111",
		91176 to 91176 => "11111111",
		91207 to 91207 => "11111111",
		91238 to 91238 => "11111111",
		92169 to 92169 => "11111111",
		92200 to 92200 => "11111111",
		92231 to 92231 => "11111111",
		92262 to 92262 => "11111111",
		93193 to 93193 => "11111111",
		93224 to 93224 => "11111111",
		93255 to 93255 => "11111111",
		93286 to 93286 => "11111111",
		94217 to 94217 => "11111111",
		94248 to 94248 => "11111111",
		94279 to 94279 => "11111111",
		94310 to 94310 => "11111111",
		95241 to 95241 => "11111111",
		95272 to 95272 => "11111111",
		95303 to 95303 => "11111111",
		95334 to 95334 => "11111111",
		96265 to 96265 => "11111111",
		96296 to 96296 => "11111111",
		96327 to 96327 => "11111111",
		96358 to 96358 => "11111111",
		97289 to 97289 => "11111111",
		97320 to 97320 => "11111111",
		97351 to 97351 => "11111111",
		97382 to 97382 => "11111111",
		98313 to 98313 => "11111111",
		98344 to 98344 => "11111111",
		98375 to 98375 => "11111111",
		98406 to 98406 => "11111111",
		99337 to 99337 => "11111111",
		99368 to 99368 => "11111111",
		99399 to 99399 => "11111111",
		99430 to 99430 => "11111111",
		100361 to 100361 => "11111111",
		100392 to 100392 => "11111111",
		100423 to 100423 => "11111111",
		100454 to 100454 => "11111111",
		101385 to 101385 => "11111111",
		101416 to 101416 => "11111111",
		101447 to 101447 => "11111111",
		101478 to 101478 => "11111111",
		102409 to 102409 => "11111111",
		102440 to 102440 => "11111111",
		102471 to 102471 => "11111111",
		102502 to 102502 => "11111111",
		103433 to 103433 => "11111111",
		103464 to 103464 => "11111111",
		103495 to 103495 => "11111111",
		103526 to 103526 => "11111111",
		104457 to 104550 => "11111111",
		others=> "00000000");
begin

	process (Clk)
	begin
		if (Clk'event and Clk = '1') then
			if (CE = '1') then
				if (Enable_w = '1') then
					VRAM (to_integer(unsigned(Addr_w))) <= Data_in;
				end if;
				Data_out <= VRAM(to_integer(unsigned(Addr_r)));
			else
				NULL;
			end if;
		end if;
	end process;

end Behavioral;

					
