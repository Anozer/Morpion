library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity ROM_victoire is
	port (CLK : in std_logic;
		  EN : in std_logic;
		  ADDR : in std_logic_vector(13 downto 0);
		  DATA : out std_logic);
end ROM_victoire;

architecture Behavioral of ROM_victoire is

type zone_memoire is array ((2**14)-1 downto 0) of std_logic;
constant ROM: zone_memoire := (
		0 => '1',
		1 => '1',
		2 => '1',
		3 => '1',
		4 => '1',
		5 => '1',
		6 => '1',
		7 => '1',
		8 => '1',
		9 => '1',
		10 => '1',
		11 => '1',
		12 => '1',
		13 => '0',
		14 => '0',
		15 => '1',
		16 => '1',
		17 => '1',
		18 => '1',
		19 => '1',
		20 => '1',
		21 => '1',
		22 => '1',
		23 => '0',
		24 => '0',
		25 => '1',
		26 => '1',
		27 => '1',
		28 => '1',
		29 => '1',
		30 => '1',
		31 => '1',
		32 => '1',
		33 => '1',
		34 => '1',
		35 => '1',
		36 => '1',
		37 => '1',
		38 => '0',
		39 => '0',
		40 => '1',
		41 => '1',
		42 => '1',
		43 => '1',
		44 => '1',
		45 => '1',
		46 => '1',
		47 => '1',
		48 => '1',
		49 => '1',
		50 => '1',
		51 => '1',
		52 => '1',
		53 => '0',
		54 => '0',
		55 => '1',
		56 => '1',
		57 => '1',
		58 => '1',
		59 => '1',
		60 => '1',
		61 => '1',
		62 => '1',
		63 => '1',
		64 => '1',
		65 => '1',
		66 => '1',
		67 => '1',
		68 => '0',
		69 => '0',
		70 => '1',
		71 => '1',
		72 => '1',
		73 => '1',
		74 => '1',
		75 => '1',
		76 => '1',
		77 => '1',
		78 => '0',
		79 => '0',
		80 => '1',
		81 => '1',
		82 => '1',
		83 => '1',
		84 => '1',
		85 => '1',
		86 => '1',
		87 => '1',
		88 => '1',
		89 => '1',
		90 => '1',
		91 => '1',
		92 => '1',
		93 => '0',
		94 => '0',
		95 => '1',
		96 => '1',
		97 => '1',
		98 => '1',
		99 => '1',
		100 => '1',
		101 => '1',
		102 => '1',
		103 => '1',
		104 => '1',
		105 => '1',
		106 => '1',
		107 => '1',
		108 => '0',
		109 => '0',
		110 => '1',
		111 => '1',
		112 => '1',
		113 => '1',
		114 => '1',
		115 => '1',
		116 => '1',
		117 => '1',
		118 => '0',
		119 => '0',
		128 => '1',
		129 => '1',
		130 => '1',
		131 => '1',
		132 => '1',
		133 => '1',
		134 => '1',
		135 => '1',
		136 => '1',
		137 => '1',
		138 => '1',
		139 => '1',
		140 => '1',
		141 => '0',
		142 => '0',
		143 => '1',
		144 => '1',
		145 => '1',
		146 => '1',
		147 => '1',
		148 => '1',
		149 => '1',
		150 => '1',
		151 => '0',
		152 => '0',
		153 => '1',
		154 => '1',
		155 => '1',
		156 => '1',
		157 => '1',
		158 => '1',
		159 => '1',
		160 => '1',
		161 => '1',
		162 => '1',
		163 => '1',
		164 => '1',
		165 => '1',
		166 => '0',
		167 => '0',
		168 => '1',
		169 => '1',
		170 => '1',
		171 => '1',
		172 => '1',
		173 => '1',
		174 => '1',
		175 => '1',
		176 => '1',
		177 => '1',
		178 => '1',
		179 => '1',
		180 => '1',
		181 => '0',
		182 => '0',
		183 => '1',
		184 => '1',
		185 => '1',
		186 => '1',
		187 => '1',
		188 => '1',
		189 => '1',
		190 => '1',
		191 => '1',
		192 => '1',
		193 => '1',
		194 => '1',
		195 => '1',
		196 => '0',
		197 => '0',
		198 => '1',
		199 => '1',
		200 => '1',
		201 => '1',
		202 => '1',
		203 => '1',
		204 => '1',
		205 => '1',
		206 => '0',
		207 => '0',
		208 => '1',
		209 => '1',
		210 => '1',
		211 => '1',
		212 => '1',
		213 => '1',
		214 => '1',
		215 => '1',
		216 => '1',
		217 => '1',
		218 => '1',
		219 => '1',
		220 => '1',
		221 => '0',
		222 => '0',
		223 => '1',
		224 => '1',
		225 => '1',
		226 => '1',
		227 => '1',
		228 => '1',
		229 => '1',
		230 => '1',
		231 => '1',
		232 => '1',
		233 => '1',
		234 => '1',
		235 => '1',
		236 => '0',
		237 => '0',
		238 => '1',
		239 => '1',
		240 => '1',
		241 => '1',
		242 => '1',
		243 => '1',
		244 => '1',
		245 => '1',
		246 => '0',
		247 => '0',
		256 => '1',
		257 => '1',
		258 => '1',
		259 => '1',
		260 => '1',
		261 => '1',
		262 => '1',
		263 => '1',
		264 => '1',
		265 => '1',
		266 => '1',
		267 => '1',
		268 => '1',
		269 => '0',
		270 => '0',
		271 => '1',
		272 => '1',
		273 => '1',
		274 => '1',
		275 => '1',
		276 => '1',
		277 => '1',
		278 => '1',
		279 => '0',
		280 => '0',
		281 => '1',
		282 => '1',
		283 => '1',
		284 => '1',
		285 => '1',
		286 => '1',
		287 => '1',
		288 => '1',
		289 => '1',
		290 => '1',
		291 => '1',
		292 => '1',
		293 => '1',
		294 => '0',
		295 => '0',
		296 => '1',
		297 => '1',
		298 => '1',
		299 => '1',
		300 => '1',
		301 => '1',
		302 => '1',
		303 => '1',
		304 => '1',
		305 => '1',
		306 => '1',
		307 => '1',
		308 => '1',
		309 => '0',
		310 => '0',
		311 => '1',
		312 => '1',
		313 => '1',
		314 => '1',
		315 => '1',
		316 => '1',
		317 => '1',
		318 => '1',
		319 => '1',
		320 => '1',
		321 => '1',
		322 => '1',
		323 => '1',
		324 => '0',
		325 => '0',
		326 => '1',
		327 => '1',
		328 => '1',
		329 => '1',
		330 => '1',
		331 => '1',
		332 => '1',
		333 => '1',
		334 => '0',
		335 => '0',
		336 => '1',
		337 => '1',
		338 => '1',
		339 => '1',
		340 => '1',
		341 => '1',
		342 => '1',
		343 => '1',
		344 => '1',
		345 => '1',
		346 => '1',
		347 => '1',
		348 => '1',
		349 => '0',
		350 => '0',
		351 => '1',
		352 => '1',
		353 => '1',
		354 => '1',
		355 => '1',
		356 => '1',
		357 => '1',
		358 => '1',
		359 => '1',
		360 => '1',
		361 => '1',
		362 => '1',
		363 => '1',
		364 => '0',
		365 => '0',
		366 => '1',
		367 => '1',
		368 => '1',
		369 => '1',
		370 => '1',
		371 => '1',
		372 => '1',
		373 => '1',
		374 => '0',
		375 => '0',
		384 => '1',
		385 => '1',
		386 => '1',
		387 => '0',
		388 => '0',
		389 => '1',
		390 => '1',
		391 => '1',
		392 => '0',
		393 => '0',
		394 => '1',
		395 => '1',
		396 => '1',
		397 => '0',
		398 => '0',
		399 => '1',
		400 => '1',
		401 => '1',
		402 => '0',
		403 => '0',
		404 => '1',
		405 => '1',
		406 => '1',
		407 => '0',
		408 => '0',
		409 => '1',
		410 => '1',
		411 => '1',
		412 => '0',
		413 => '0',
		414 => '0',
		415 => '0',
		416 => '0',
		417 => '0',
		418 => '0',
		419 => '1',
		420 => '1',
		421 => '1',
		422 => '0',
		423 => '0',
		424 => '1',
		425 => '1',
		426 => '1',
		427 => '0',
		428 => '0',
		429 => '0',
		430 => '0',
		431 => '0',
		432 => '0',
		433 => '0',
		434 => '1',
		435 => '1',
		436 => '1',
		437 => '0',
		438 => '0',
		439 => '1',
		440 => '1',
		441 => '1',
		442 => '0',
		443 => '0',
		444 => '0',
		445 => '0',
		446 => '0',
		447 => '0',
		448 => '0',
		449 => '1',
		450 => '1',
		451 => '1',
		452 => '0',
		453 => '0',
		454 => '1',
		455 => '1',
		456 => '1',
		457 => '0',
		458 => '0',
		459 => '1',
		460 => '1',
		461 => '1',
		462 => '0',
		463 => '0',
		464 => '1',
		465 => '1',
		466 => '1',
		467 => '0',
		468 => '0',
		469 => '0',
		470 => '0',
		471 => '0',
		472 => '0',
		473 => '0',
		474 => '1',
		475 => '1',
		476 => '1',
		477 => '0',
		478 => '0',
		479 => '1',
		480 => '1',
		481 => '1',
		482 => '0',
		483 => '0',
		484 => '0',
		485 => '0',
		486 => '0',
		487 => '0',
		488 => '0',
		489 => '1',
		490 => '1',
		491 => '1',
		492 => '0',
		493 => '0',
		494 => '1',
		495 => '1',
		496 => '1',
		497 => '0',
		498 => '0',
		499 => '1',
		500 => '1',
		501 => '1',
		502 => '0',
		503 => '0',
		512 => '1',
		513 => '1',
		514 => '1',
		515 => '0',
		516 => '0',
		517 => '1',
		518 => '1',
		519 => '1',
		520 => '0',
		521 => '0',
		522 => '1',
		523 => '1',
		524 => '1',
		525 => '0',
		526 => '0',
		527 => '1',
		528 => '1',
		529 => '1',
		530 => '0',
		531 => '0',
		532 => '1',
		533 => '1',
		534 => '1',
		535 => '0',
		536 => '0',
		537 => '1',
		538 => '1',
		539 => '1',
		540 => '0',
		541 => '0',
		542 => '0',
		543 => '0',
		544 => '0',
		545 => '0',
		546 => '0',
		547 => '1',
		548 => '1',
		549 => '1',
		550 => '0',
		551 => '0',
		552 => '1',
		553 => '1',
		554 => '1',
		555 => '0',
		556 => '0',
		557 => '0',
		558 => '0',
		559 => '0',
		560 => '0',
		561 => '0',
		562 => '1',
		563 => '1',
		564 => '1',
		565 => '0',
		566 => '0',
		567 => '1',
		568 => '1',
		569 => '1',
		570 => '0',
		571 => '0',
		572 => '0',
		573 => '0',
		574 => '0',
		575 => '0',
		576 => '0',
		577 => '1',
		578 => '1',
		579 => '1',
		580 => '0',
		581 => '0',
		582 => '1',
		583 => '1',
		584 => '1',
		585 => '0',
		586 => '0',
		587 => '1',
		588 => '1',
		589 => '1',
		590 => '0',
		591 => '0',
		592 => '1',
		593 => '1',
		594 => '1',
		595 => '0',
		596 => '0',
		597 => '0',
		598 => '0',
		599 => '0',
		600 => '0',
		601 => '0',
		602 => '1',
		603 => '1',
		604 => '1',
		605 => '0',
		606 => '0',
		607 => '1',
		608 => '1',
		609 => '1',
		610 => '0',
		611 => '0',
		612 => '0',
		613 => '0',
		614 => '0',
		615 => '0',
		616 => '0',
		617 => '1',
		618 => '1',
		619 => '1',
		620 => '0',
		621 => '0',
		622 => '1',
		623 => '1',
		624 => '1',
		625 => '0',
		626 => '0',
		627 => '1',
		628 => '1',
		629 => '1',
		630 => '0',
		631 => '0',
		640 => '1',
		641 => '1',
		642 => '1',
		643 => '0',
		644 => '0',
		645 => '1',
		646 => '1',
		647 => '1',
		648 => '0',
		649 => '0',
		650 => '1',
		651 => '1',
		652 => '1',
		653 => '0',
		654 => '0',
		655 => '1',
		656 => '1',
		657 => '1',
		658 => '0',
		659 => '0',
		660 => '1',
		661 => '1',
		662 => '1',
		663 => '0',
		664 => '0',
		665 => '1',
		666 => '1',
		667 => '1',
		668 => '0',
		669 => '0',
		670 => '0',
		671 => '0',
		672 => '0',
		673 => '0',
		674 => '0',
		675 => '1',
		676 => '1',
		677 => '1',
		678 => '0',
		679 => '0',
		680 => '1',
		681 => '1',
		682 => '1',
		683 => '1',
		684 => '1',
		685 => '1',
		686 => '0',
		687 => '1',
		688 => '1',
		689 => '1',
		690 => '1',
		691 => '1',
		692 => '1',
		693 => '0',
		694 => '0',
		695 => '1',
		696 => '1',
		697 => '1',
		698 => '0',
		699 => '0',
		700 => '0',
		701 => '0',
		702 => '0',
		703 => '0',
		704 => '0',
		705 => '1',
		706 => '1',
		707 => '1',
		708 => '0',
		709 => '0',
		710 => '1',
		711 => '1',
		712 => '1',
		713 => '0',
		714 => '0',
		715 => '1',
		716 => '1',
		717 => '1',
		718 => '0',
		719 => '0',
		720 => '1',
		721 => '1',
		722 => '1',
		723 => '0',
		724 => '0',
		725 => '1',
		726 => '1',
		727 => '1',
		728 => '0',
		729 => '0',
		730 => '1',
		731 => '1',
		732 => '1',
		733 => '0',
		734 => '0',
		735 => '1',
		736 => '1',
		737 => '1',
		738 => '0',
		739 => '0',
		740 => '1',
		741 => '1',
		742 => '1',
		743 => '1',
		744 => '1',
		745 => '1',
		746 => '1',
		747 => '1',
		748 => '0',
		749 => '0',
		750 => '1',
		751 => '1',
		752 => '1',
		753 => '0',
		754 => '0',
		755 => '1',
		756 => '1',
		757 => '1',
		758 => '0',
		759 => '0',
		768 => '1',
		769 => '1',
		770 => '1',
		771 => '0',
		772 => '0',
		773 => '1',
		774 => '1',
		775 => '1',
		776 => '0',
		777 => '0',
		778 => '1',
		779 => '1',
		780 => '1',
		781 => '0',
		782 => '0',
		783 => '1',
		784 => '1',
		785 => '1',
		786 => '0',
		787 => '0',
		788 => '1',
		789 => '1',
		790 => '1',
		791 => '0',
		792 => '0',
		793 => '1',
		794 => '1',
		795 => '1',
		796 => '0',
		797 => '0',
		798 => '1',
		799 => '1',
		800 => '1',
		801 => '0',
		802 => '0',
		803 => '1',
		804 => '1',
		805 => '1',
		806 => '0',
		807 => '0',
		808 => '1',
		809 => '1',
		810 => '1',
		811 => '1',
		812 => '1',
		813 => '1',
		814 => '0',
		815 => '1',
		816 => '1',
		817 => '1',
		818 => '1',
		819 => '1',
		820 => '1',
		821 => '0',
		822 => '0',
		823 => '1',
		824 => '1',
		825 => '1',
		826 => '0',
		827 => '0',
		828 => '1',
		829 => '1',
		830 => '1',
		831 => '0',
		832 => '0',
		833 => '1',
		834 => '1',
		835 => '1',
		836 => '0',
		837 => '0',
		838 => '1',
		839 => '1',
		840 => '1',
		841 => '0',
		842 => '0',
		843 => '1',
		844 => '1',
		845 => '1',
		846 => '0',
		847 => '0',
		848 => '1',
		849 => '1',
		850 => '1',
		851 => '0',
		852 => '0',
		853 => '1',
		854 => '1',
		855 => '1',
		856 => '0',
		857 => '0',
		858 => '1',
		859 => '1',
		860 => '1',
		861 => '0',
		862 => '0',
		863 => '1',
		864 => '1',
		865 => '1',
		866 => '0',
		867 => '0',
		868 => '1',
		869 => '1',
		870 => '1',
		871 => '1',
		872 => '1',
		873 => '1',
		874 => '1',
		875 => '1',
		876 => '0',
		877 => '0',
		878 => '1',
		879 => '1',
		880 => '1',
		881 => '0',
		882 => '0',
		883 => '1',
		884 => '1',
		885 => '1',
		886 => '0',
		887 => '0',
		896 => '1',
		897 => '1',
		898 => '1',
		899 => '0',
		900 => '0',
		901 => '1',
		902 => '1',
		903 => '1',
		904 => '0',
		905 => '0',
		906 => '1',
		907 => '1',
		908 => '1',
		909 => '0',
		910 => '0',
		911 => '1',
		912 => '1',
		913 => '1',
		914 => '0',
		915 => '0',
		916 => '1',
		917 => '1',
		918 => '1',
		919 => '0',
		920 => '0',
		921 => '1',
		922 => '1',
		923 => '1',
		924 => '0',
		925 => '0',
		926 => '1',
		927 => '1',
		928 => '1',
		929 => '0',
		930 => '0',
		931 => '1',
		932 => '1',
		933 => '1',
		934 => '0',
		935 => '0',
		936 => '1',
		937 => '1',
		938 => '1',
		939 => '1',
		940 => '1',
		941 => '1',
		942 => '0',
		943 => '1',
		944 => '1',
		945 => '1',
		946 => '1',
		947 => '1',
		948 => '1',
		949 => '0',
		950 => '0',
		951 => '1',
		952 => '1',
		953 => '1',
		954 => '0',
		955 => '0',
		956 => '1',
		957 => '1',
		958 => '1',
		959 => '0',
		960 => '0',
		961 => '1',
		962 => '1',
		963 => '1',
		964 => '0',
		965 => '0',
		966 => '1',
		967 => '1',
		968 => '1',
		969 => '0',
		970 => '0',
		971 => '1',
		972 => '1',
		973 => '1',
		974 => '0',
		975 => '0',
		976 => '1',
		977 => '1',
		978 => '1',
		979 => '0',
		980 => '0',
		981 => '1',
		982 => '1',
		983 => '1',
		984 => '0',
		985 => '0',
		986 => '1',
		987 => '1',
		988 => '1',
		989 => '0',
		990 => '0',
		991 => '1',
		992 => '1',
		993 => '1',
		994 => '0',
		995 => '0',
		996 => '1',
		997 => '1',
		998 => '1',
		999 => '1',
		1000 => '1',
		1001 => '1',
		1002 => '1',
		1003 => '1',
		1004 => '0',
		1005 => '0',
		1006 => '1',
		1007 => '1',
		1008 => '1',
		1009 => '0',
		1010 => '0',
		1011 => '1',
		1012 => '1',
		1013 => '1',
		1014 => '0',
		1015 => '0',
		1024 => '1',
		1025 => '1',
		1026 => '1',
		1027 => '0',
		1028 => '0',
		1029 => '1',
		1030 => '1',
		1031 => '1',
		1032 => '0',
		1033 => '0',
		1034 => '1',
		1035 => '1',
		1036 => '1',
		1037 => '0',
		1038 => '0',
		1039 => '1',
		1040 => '1',
		1041 => '1',
		1042 => '0',
		1043 => '0',
		1044 => '1',
		1045 => '1',
		1046 => '1',
		1047 => '0',
		1048 => '0',
		1049 => '1',
		1050 => '1',
		1051 => '1',
		1052 => '0',
		1053 => '0',
		1054 => '1',
		1055 => '1',
		1056 => '1',
		1057 => '1',
		1058 => '1',
		1059 => '1',
		1060 => '1',
		1061 => '1',
		1062 => '0',
		1063 => '0',
		1064 => '0',
		1065 => '0',
		1066 => '0',
		1067 => '1',
		1068 => '1',
		1069 => '1',
		1070 => '0',
		1071 => '1',
		1072 => '1',
		1073 => '1',
		1074 => '0',
		1075 => '0',
		1076 => '0',
		1077 => '0',
		1078 => '0',
		1079 => '1',
		1080 => '1',
		1081 => '1',
		1082 => '0',
		1083 => '0',
		1084 => '1',
		1085 => '1',
		1086 => '1',
		1087 => '0',
		1088 => '0',
		1089 => '1',
		1090 => '1',
		1091 => '1',
		1092 => '0',
		1093 => '0',
		1094 => '1',
		1095 => '1',
		1096 => '1',
		1097 => '0',
		1098 => '0',
		1099 => '1',
		1100 => '1',
		1101 => '1',
		1102 => '0',
		1103 => '0',
		1104 => '1',
		1105 => '1',
		1106 => '1',
		1107 => '0',
		1108 => '0',
		1109 => '0',
		1110 => '0',
		1111 => '0',
		1112 => '1',
		1113 => '1',
		1114 => '1',
		1115 => '1',
		1116 => '1',
		1117 => '0',
		1118 => '0',
		1119 => '1',
		1120 => '1',
		1121 => '1',
		1122 => '0',
		1123 => '0',
		1124 => '0',
		1125 => '0',
		1126 => '0',
		1127 => '0',
		1128 => '0',
		1129 => '1',
		1130 => '1',
		1131 => '1',
		1132 => '0',
		1133 => '0',
		1134 => '1',
		1135 => '1',
		1136 => '1',
		1137 => '0',
		1138 => '0',
		1139 => '1',
		1140 => '1',
		1141 => '1',
		1142 => '0',
		1143 => '0',
		1152 => '1',
		1153 => '1',
		1154 => '1',
		1155 => '0',
		1156 => '0',
		1157 => '1',
		1158 => '1',
		1159 => '1',
		1160 => '0',
		1161 => '0',
		1162 => '1',
		1163 => '1',
		1164 => '1',
		1165 => '0',
		1166 => '0',
		1167 => '1',
		1168 => '1',
		1169 => '1',
		1170 => '0',
		1171 => '0',
		1172 => '1',
		1173 => '1',
		1174 => '1',
		1175 => '0',
		1176 => '0',
		1177 => '1',
		1178 => '1',
		1179 => '1',
		1180 => '0',
		1181 => '0',
		1182 => '1',
		1183 => '1',
		1184 => '1',
		1185 => '1',
		1186 => '1',
		1187 => '1',
		1188 => '1',
		1189 => '1',
		1190 => '0',
		1191 => '0',
		1192 => '0',
		1193 => '0',
		1194 => '0',
		1195 => '1',
		1196 => '1',
		1197 => '1',
		1198 => '0',
		1199 => '1',
		1200 => '1',
		1201 => '1',
		1202 => '0',
		1203 => '0',
		1204 => '0',
		1205 => '0',
		1206 => '0',
		1207 => '1',
		1208 => '1',
		1209 => '1',
		1210 => '0',
		1211 => '0',
		1212 => '1',
		1213 => '1',
		1214 => '1',
		1215 => '0',
		1216 => '0',
		1217 => '1',
		1218 => '1',
		1219 => '1',
		1220 => '0',
		1221 => '0',
		1222 => '1',
		1223 => '1',
		1224 => '1',
		1225 => '0',
		1226 => '0',
		1227 => '1',
		1228 => '1',
		1229 => '1',
		1230 => '0',
		1231 => '0',
		1232 => '1',
		1233 => '1',
		1234 => '1',
		1235 => '0',
		1236 => '0',
		1237 => '0',
		1238 => '0',
		1239 => '0',
		1240 => '1',
		1241 => '1',
		1242 => '1',
		1243 => '1',
		1244 => '1',
		1245 => '0',
		1246 => '0',
		1247 => '1',
		1248 => '1',
		1249 => '1',
		1250 => '0',
		1251 => '0',
		1252 => '0',
		1253 => '0',
		1254 => '0',
		1255 => '0',
		1256 => '0',
		1257 => '1',
		1258 => '1',
		1259 => '1',
		1260 => '0',
		1261 => '0',
		1262 => '1',
		1263 => '1',
		1264 => '1',
		1265 => '0',
		1266 => '0',
		1267 => '1',
		1268 => '1',
		1269 => '1',
		1270 => '0',
		1271 => '0',
		1280 => '1',
		1281 => '1',
		1282 => '1',
		1283 => '0',
		1284 => '0',
		1285 => '1',
		1286 => '1',
		1287 => '1',
		1288 => '0',
		1289 => '0',
		1290 => '1',
		1291 => '1',
		1292 => '1',
		1293 => '0',
		1294 => '0',
		1295 => '1',
		1296 => '1',
		1297 => '1',
		1298 => '0',
		1299 => '0',
		1300 => '1',
		1301 => '1',
		1302 => '1',
		1303 => '0',
		1304 => '0',
		1305 => '1',
		1306 => '1',
		1307 => '1',
		1308 => '0',
		1309 => '0',
		1310 => '1',
		1311 => '1',
		1312 => '1',
		1313 => '1',
		1314 => '1',
		1315 => '1',
		1316 => '1',
		1317 => '1',
		1318 => '0',
		1319 => '0',
		1320 => '0',
		1321 => '0',
		1322 => '0',
		1323 => '1',
		1324 => '1',
		1325 => '1',
		1326 => '0',
		1327 => '1',
		1328 => '1',
		1329 => '1',
		1330 => '0',
		1331 => '0',
		1332 => '0',
		1333 => '0',
		1334 => '0',
		1335 => '1',
		1336 => '1',
		1337 => '1',
		1338 => '0',
		1339 => '0',
		1340 => '1',
		1341 => '1',
		1342 => '1',
		1343 => '0',
		1344 => '0',
		1345 => '1',
		1346 => '1',
		1347 => '1',
		1348 => '0',
		1349 => '0',
		1350 => '1',
		1351 => '1',
		1352 => '1',
		1353 => '0',
		1354 => '0',
		1355 => '1',
		1356 => '1',
		1357 => '1',
		1358 => '0',
		1359 => '0',
		1360 => '1',
		1361 => '1',
		1362 => '1',
		1363 => '0',
		1364 => '0',
		1365 => '1',
		1366 => '1',
		1367 => '1',
		1368 => '1',
		1369 => '1',
		1370 => '1',
		1371 => '1',
		1372 => '1',
		1373 => '0',
		1374 => '0',
		1375 => '1',
		1376 => '1',
		1377 => '1',
		1378 => '0',
		1379 => '0',
		1380 => '1',
		1381 => '1',
		1382 => '1',
		1383 => '1',
		1384 => '1',
		1385 => '1',
		1386 => '1',
		1387 => '1',
		1388 => '0',
		1389 => '0',
		1390 => '1',
		1391 => '1',
		1392 => '1',
		1393 => '1',
		1394 => '1',
		1395 => '1',
		1396 => '1',
		1397 => '1',
		1398 => '0',
		1399 => '0',
		1408 => '1',
		1409 => '1',
		1410 => '1',
		1411 => '0',
		1412 => '0',
		1413 => '1',
		1414 => '1',
		1415 => '1',
		1416 => '0',
		1417 => '0',
		1418 => '1',
		1419 => '1',
		1420 => '1',
		1421 => '0',
		1422 => '0',
		1423 => '1',
		1424 => '1',
		1425 => '1',
		1426 => '0',
		1427 => '0',
		1428 => '1',
		1429 => '1',
		1430 => '1',
		1431 => '0',
		1432 => '0',
		1433 => '1',
		1434 => '1',
		1435 => '1',
		1436 => '0',
		1437 => '0',
		1438 => '1',
		1439 => '1',
		1440 => '1',
		1441 => '0',
		1442 => '0',
		1443 => '1',
		1444 => '1',
		1445 => '1',
		1446 => '0',
		1447 => '0',
		1448 => '0',
		1449 => '0',
		1450 => '0',
		1451 => '1',
		1452 => '1',
		1453 => '1',
		1454 => '0',
		1455 => '1',
		1456 => '1',
		1457 => '1',
		1458 => '0',
		1459 => '0',
		1460 => '0',
		1461 => '0',
		1462 => '0',
		1463 => '1',
		1464 => '1',
		1465 => '1',
		1466 => '0',
		1467 => '0',
		1468 => '1',
		1469 => '1',
		1470 => '1',
		1471 => '0',
		1472 => '0',
		1473 => '1',
		1474 => '1',
		1475 => '1',
		1476 => '0',
		1477 => '0',
		1478 => '1',
		1479 => '1',
		1480 => '1',
		1481 => '0',
		1482 => '0',
		1483 => '1',
		1484 => '1',
		1485 => '1',
		1486 => '0',
		1487 => '0',
		1488 => '1',
		1489 => '1',
		1490 => '1',
		1491 => '0',
		1492 => '0',
		1493 => '1',
		1494 => '1',
		1495 => '1',
		1496 => '0',
		1497 => '0',
		1498 => '1',
		1499 => '1',
		1500 => '1',
		1501 => '0',
		1502 => '0',
		1503 => '1',
		1504 => '1',
		1505 => '1',
		1506 => '0',
		1507 => '0',
		1508 => '1',
		1509 => '1',
		1510 => '1',
		1511 => '1',
		1512 => '1',
		1513 => '1',
		1514 => '1',
		1515 => '1',
		1516 => '0',
		1517 => '0',
		1518 => '1',
		1519 => '1',
		1520 => '1',
		1521 => '1',
		1522 => '1',
		1523 => '1',
		1524 => '1',
		1525 => '1',
		1526 => '0',
		1527 => '0',
		1536 => '1',
		1537 => '1',
		1538 => '1',
		1539 => '0',
		1540 => '0',
		1541 => '1',
		1542 => '1',
		1543 => '1',
		1544 => '0',
		1545 => '0',
		1546 => '1',
		1547 => '1',
		1548 => '1',
		1549 => '0',
		1550 => '0',
		1551 => '1',
		1552 => '1',
		1553 => '1',
		1554 => '0',
		1555 => '0',
		1556 => '1',
		1557 => '1',
		1558 => '1',
		1559 => '0',
		1560 => '0',
		1561 => '1',
		1562 => '1',
		1563 => '1',
		1564 => '0',
		1565 => '0',
		1566 => '1',
		1567 => '1',
		1568 => '1',
		1569 => '0',
		1570 => '0',
		1571 => '1',
		1572 => '1',
		1573 => '1',
		1574 => '0',
		1575 => '0',
		1576 => '0',
		1577 => '0',
		1578 => '0',
		1579 => '1',
		1580 => '1',
		1581 => '1',
		1582 => '0',
		1583 => '1',
		1584 => '1',
		1585 => '1',
		1586 => '0',
		1587 => '0',
		1588 => '0',
		1589 => '0',
		1590 => '0',
		1591 => '1',
		1592 => '1',
		1593 => '1',
		1594 => '0',
		1595 => '0',
		1596 => '1',
		1597 => '1',
		1598 => '1',
		1599 => '0',
		1600 => '0',
		1601 => '1',
		1602 => '1',
		1603 => '1',
		1604 => '0',
		1605 => '0',
		1606 => '1',
		1607 => '1',
		1608 => '1',
		1609 => '0',
		1610 => '0',
		1611 => '1',
		1612 => '1',
		1613 => '1',
		1614 => '0',
		1615 => '0',
		1616 => '1',
		1617 => '1',
		1618 => '1',
		1619 => '0',
		1620 => '0',
		1621 => '1',
		1622 => '1',
		1623 => '1',
		1624 => '0',
		1625 => '0',
		1626 => '1',
		1627 => '1',
		1628 => '1',
		1629 => '0',
		1630 => '0',
		1631 => '1',
		1632 => '1',
		1633 => '1',
		1634 => '0',
		1635 => '0',
		1636 => '1',
		1637 => '1',
		1638 => '1',
		1639 => '1',
		1640 => '1',
		1641 => '1',
		1642 => '1',
		1643 => '1',
		1644 => '0',
		1645 => '0',
		1646 => '1',
		1647 => '1',
		1648 => '1',
		1649 => '1',
		1650 => '1',
		1651 => '1',
		1652 => '1',
		1653 => '1',
		1654 => '0',
		1655 => '0',
		1664 => '1',
		1665 => '1',
		1666 => '1',
		1667 => '1',
		1668 => '1',
		1669 => '0',
		1670 => '0',
		1671 => '0',
		1672 => '1',
		1673 => '1',
		1674 => '1',
		1675 => '1',
		1676 => '1',
		1677 => '0',
		1678 => '0',
		1679 => '1',
		1680 => '1',
		1681 => '1',
		1682 => '0',
		1683 => '0',
		1684 => '1',
		1685 => '1',
		1686 => '1',
		1687 => '0',
		1688 => '0',
		1689 => '1',
		1690 => '1',
		1691 => '1',
		1692 => '0',
		1693 => '0',
		1694 => '0',
		1695 => '0',
		1696 => '0',
		1697 => '0',
		1698 => '0',
		1699 => '1',
		1700 => '1',
		1701 => '1',
		1702 => '0',
		1703 => '0',
		1704 => '0',
		1705 => '0',
		1706 => '0',
		1707 => '1',
		1708 => '1',
		1709 => '1',
		1710 => '0',
		1711 => '1',
		1712 => '1',
		1713 => '1',
		1714 => '0',
		1715 => '0',
		1716 => '0',
		1717 => '0',
		1718 => '0',
		1719 => '1',
		1720 => '1',
		1721 => '1',
		1722 => '0',
		1723 => '0',
		1724 => '0',
		1725 => '0',
		1726 => '0',
		1727 => '0',
		1728 => '0',
		1729 => '1',
		1730 => '1',
		1731 => '1',
		1732 => '0',
		1733 => '0',
		1734 => '1',
		1735 => '1',
		1736 => '1',
		1737 => '0',
		1738 => '0',
		1739 => '1',
		1740 => '1',
		1741 => '1',
		1742 => '0',
		1743 => '0',
		1744 => '1',
		1745 => '1',
		1746 => '1',
		1747 => '0',
		1748 => '0',
		1749 => '1',
		1750 => '1',
		1751 => '1',
		1752 => '0',
		1753 => '0',
		1754 => '1',
		1755 => '1',
		1756 => '1',
		1757 => '0',
		1758 => '0',
		1759 => '1',
		1760 => '1',
		1761 => '1',
		1762 => '0',
		1763 => '0',
		1764 => '0',
		1765 => '0',
		1766 => '0',
		1767 => '0',
		1768 => '0',
		1769 => '1',
		1770 => '1',
		1771 => '1',
		1772 => '0',
		1773 => '0',
		1774 => '1',
		1775 => '1',
		1776 => '1',
		1777 => '0',
		1778 => '0',
		1779 => '1',
		1780 => '1',
		1781 => '1',
		1782 => '0',
		1783 => '0',
		1792 => '1',
		1793 => '1',
		1794 => '1',
		1795 => '1',
		1796 => '1',
		1797 => '0',
		1798 => '0',
		1799 => '0',
		1800 => '1',
		1801 => '1',
		1802 => '1',
		1803 => '1',
		1804 => '1',
		1805 => '0',
		1806 => '0',
		1807 => '1',
		1808 => '1',
		1809 => '1',
		1810 => '0',
		1811 => '0',
		1812 => '1',
		1813 => '1',
		1814 => '1',
		1815 => '0',
		1816 => '0',
		1817 => '1',
		1818 => '1',
		1819 => '1',
		1820 => '0',
		1821 => '0',
		1822 => '0',
		1823 => '0',
		1824 => '0',
		1825 => '0',
		1826 => '0',
		1827 => '1',
		1828 => '1',
		1829 => '1',
		1830 => '0',
		1831 => '0',
		1832 => '0',
		1833 => '0',
		1834 => '0',
		1835 => '1',
		1836 => '1',
		1837 => '1',
		1838 => '0',
		1839 => '1',
		1840 => '1',
		1841 => '1',
		1842 => '0',
		1843 => '0',
		1844 => '0',
		1845 => '0',
		1846 => '0',
		1847 => '1',
		1848 => '1',
		1849 => '1',
		1850 => '0',
		1851 => '0',
		1852 => '0',
		1853 => '0',
		1854 => '0',
		1855 => '0',
		1856 => '0',
		1857 => '1',
		1858 => '1',
		1859 => '1',
		1860 => '0',
		1861 => '0',
		1862 => '1',
		1863 => '1',
		1864 => '1',
		1865 => '0',
		1866 => '0',
		1867 => '1',
		1868 => '1',
		1869 => '1',
		1870 => '0',
		1871 => '0',
		1872 => '1',
		1873 => '1',
		1874 => '1',
		1875 => '0',
		1876 => '0',
		1877 => '1',
		1878 => '1',
		1879 => '1',
		1880 => '0',
		1881 => '0',
		1882 => '1',
		1883 => '1',
		1884 => '1',
		1885 => '0',
		1886 => '0',
		1887 => '1',
		1888 => '1',
		1889 => '1',
		1890 => '0',
		1891 => '0',
		1892 => '0',
		1893 => '0',
		1894 => '0',
		1895 => '0',
		1896 => '0',
		1897 => '1',
		1898 => '1',
		1899 => '1',
		1900 => '0',
		1901 => '0',
		1902 => '1',
		1903 => '1',
		1904 => '1',
		1905 => '0',
		1906 => '0',
		1907 => '1',
		1908 => '1',
		1909 => '1',
		1910 => '0',
		1911 => '0',
		1920 => '0',
		1921 => '0',
		1922 => '0',
		1923 => '1',
		1924 => '1',
		1925 => '1',
		1926 => '1',
		1927 => '1',
		1928 => '1',
		1929 => '1',
		1930 => '0',
		1931 => '0',
		1932 => '0',
		1933 => '0',
		1934 => '0',
		1935 => '1',
		1936 => '1',
		1937 => '1',
		1938 => '1',
		1939 => '1',
		1940 => '1',
		1941 => '1',
		1942 => '1',
		1943 => '0',
		1944 => '0',
		1945 => '1',
		1946 => '1',
		1947 => '1',
		1948 => '1',
		1949 => '1',
		1950 => '1',
		1951 => '1',
		1952 => '1',
		1953 => '1',
		1954 => '1',
		1955 => '1',
		1956 => '1',
		1957 => '1',
		1958 => '0',
		1959 => '0',
		1960 => '0',
		1961 => '0',
		1962 => '0',
		1963 => '1',
		1964 => '1',
		1965 => '1',
		1966 => '1',
		1967 => '1',
		1968 => '1',
		1969 => '1',
		1970 => '0',
		1971 => '0',
		1972 => '0',
		1973 => '0',
		1974 => '0',
		1975 => '1',
		1976 => '1',
		1977 => '1',
		1978 => '1',
		1979 => '1',
		1980 => '1',
		1981 => '1',
		1982 => '1',
		1983 => '1',
		1984 => '1',
		1985 => '1',
		1986 => '1',
		1987 => '1',
		1988 => '0',
		1989 => '0',
		1990 => '1',
		1991 => '1',
		1992 => '1',
		1993 => '1',
		1994 => '1',
		1995 => '1',
		1996 => '1',
		1997 => '1',
		1998 => '0',
		1999 => '0',
		2000 => '1',
		2001 => '1',
		2002 => '1',
		2003 => '1',
		2004 => '1',
		2005 => '1',
		2006 => '1',
		2007 => '1',
		2008 => '1',
		2009 => '1',
		2010 => '1',
		2011 => '1',
		2012 => '1',
		2013 => '0',
		2014 => '0',
		2015 => '1',
		2016 => '1',
		2017 => '1',
		2018 => '1',
		2019 => '1',
		2020 => '1',
		2021 => '1',
		2022 => '1',
		2023 => '1',
		2024 => '1',
		2025 => '1',
		2026 => '1',
		2027 => '1',
		2028 => '0',
		2029 => '0',
		2030 => '1',
		2031 => '1',
		2032 => '1',
		2033 => '1',
		2034 => '1',
		2035 => '1',
		2036 => '1',
		2037 => '1',
		2038 => '0',
		2039 => '0',
		2048 => '0',
		2049 => '0',
		2050 => '0',
		2051 => '1',
		2052 => '1',
		2053 => '1',
		2054 => '1',
		2055 => '1',
		2056 => '1',
		2057 => '1',
		2058 => '0',
		2059 => '0',
		2060 => '0',
		2061 => '0',
		2062 => '0',
		2063 => '1',
		2064 => '1',
		2065 => '1',
		2066 => '1',
		2067 => '1',
		2068 => '1',
		2069 => '1',
		2070 => '1',
		2071 => '0',
		2072 => '0',
		2073 => '1',
		2074 => '1',
		2075 => '1',
		2076 => '1',
		2077 => '1',
		2078 => '1',
		2079 => '1',
		2080 => '1',
		2081 => '1',
		2082 => '1',
		2083 => '1',
		2084 => '1',
		2085 => '1',
		2086 => '0',
		2087 => '0',
		2088 => '0',
		2089 => '0',
		2090 => '0',
		2091 => '1',
		2092 => '1',
		2093 => '1',
		2094 => '1',
		2095 => '1',
		2096 => '1',
		2097 => '1',
		2098 => '0',
		2099 => '0',
		2100 => '0',
		2101 => '0',
		2102 => '0',
		2103 => '1',
		2104 => '1',
		2105 => '1',
		2106 => '1',
		2107 => '1',
		2108 => '1',
		2109 => '1',
		2110 => '1',
		2111 => '1',
		2112 => '1',
		2113 => '1',
		2114 => '1',
		2115 => '1',
		2116 => '0',
		2117 => '0',
		2118 => '1',
		2119 => '1',
		2120 => '1',
		2121 => '1',
		2122 => '1',
		2123 => '1',
		2124 => '1',
		2125 => '1',
		2126 => '0',
		2127 => '0',
		2128 => '1',
		2129 => '1',
		2130 => '1',
		2131 => '1',
		2132 => '1',
		2133 => '1',
		2134 => '1',
		2135 => '1',
		2136 => '1',
		2137 => '1',
		2138 => '1',
		2139 => '1',
		2140 => '1',
		2141 => '0',
		2142 => '0',
		2143 => '1',
		2144 => '1',
		2145 => '1',
		2146 => '1',
		2147 => '1',
		2148 => '1',
		2149 => '1',
		2150 => '1',
		2151 => '1',
		2152 => '1',
		2153 => '1',
		2154 => '1',
		2155 => '1',
		2156 => '0',
		2157 => '0',
		2158 => '1',
		2159 => '1',
		2160 => '1',
		2161 => '1',
		2162 => '1',
		2163 => '1',
		2164 => '1',
		2165 => '1',
		2166 => '0',
		2167 => '0',
		2176 => '0',
		2177 => '0',
		2178 => '0',
		2179 => '1',
		2180 => '1',
		2181 => '1',
		2182 => '1',
		2183 => '1',
		2184 => '1',
		2185 => '1',
		2186 => '0',
		2187 => '0',
		2188 => '0',
		2189 => '0',
		2190 => '0',
		2191 => '1',
		2192 => '1',
		2193 => '1',
		2194 => '1',
		2195 => '1',
		2196 => '1',
		2197 => '1',
		2198 => '1',
		2199 => '0',
		2200 => '0',
		2201 => '1',
		2202 => '1',
		2203 => '1',
		2204 => '1',
		2205 => '1',
		2206 => '1',
		2207 => '1',
		2208 => '1',
		2209 => '1',
		2210 => '1',
		2211 => '1',
		2212 => '1',
		2213 => '1',
		2214 => '0',
		2215 => '0',
		2216 => '0',
		2217 => '0',
		2218 => '0',
		2219 => '1',
		2220 => '1',
		2221 => '1',
		2222 => '1',
		2223 => '1',
		2224 => '1',
		2225 => '1',
		2226 => '0',
		2227 => '0',
		2228 => '0',
		2229 => '0',
		2230 => '0',
		2231 => '1',
		2232 => '1',
		2233 => '1',
		2234 => '1',
		2235 => '1',
		2236 => '1',
		2237 => '1',
		2238 => '1',
		2239 => '1',
		2240 => '1',
		2241 => '1',
		2242 => '1',
		2243 => '1',
		2244 => '0',
		2245 => '0',
		2246 => '1',
		2247 => '1',
		2248 => '1',
		2249 => '1',
		2250 => '1',
		2251 => '1',
		2252 => '1',
		2253 => '1',
		2254 => '0',
		2255 => '0',
		2256 => '1',
		2257 => '1',
		2258 => '1',
		2259 => '1',
		2260 => '1',
		2261 => '1',
		2262 => '1',
		2263 => '1',
		2264 => '1',
		2265 => '1',
		2266 => '1',
		2267 => '1',
		2268 => '1',
		2269 => '0',
		2270 => '0',
		2271 => '1',
		2272 => '1',
		2273 => '1',
		2274 => '1',
		2275 => '1',
		2276 => '1',
		2277 => '1',
		2278 => '1',
		2279 => '1',
		2280 => '1',
		2281 => '1',
		2282 => '1',
		2283 => '1',
		2284 => '0',
		2285 => '0',
		2286 => '1',
		2287 => '1',
		2288 => '1',
		2289 => '1',
		2290 => '1',
		2291 => '1',
		2292 => '1',
		2293 => '1',
		2294 => '0',
		2295 => '0',
		2304 => '0',
		2305 => '0',
		2306 => '0',
		2307 => '0',
		2308 => '0',
		2309 => '0',
		2310 => '0',
		2311 => '0',
		2312 => '0',
		2313 => '0',
		2314 => '0',
		2315 => '0',
		2316 => '0',
		2317 => '0',
		2318 => '0',
		2319 => '0',
		2320 => '0',
		2321 => '0',
		2322 => '0',
		2323 => '0',
		2324 => '0',
		2325 => '0',
		2326 => '0',
		2327 => '0',
		2328 => '0',
		2329 => '0',
		2330 => '0',
		2331 => '0',
		2332 => '0',
		2333 => '0',
		2334 => '0',
		2335 => '0',
		2336 => '0',
		2337 => '0',
		2338 => '0',
		2339 => '0',
		2340 => '0',
		2341 => '0',
		2342 => '0',
		2343 => '0',
		2344 => '0',
		2345 => '0',
		2346 => '0',
		2347 => '0',
		2348 => '0',
		2349 => '0',
		2350 => '0',
		2351 => '0',
		2352 => '0',
		2353 => '0',
		2354 => '0',
		2355 => '0',
		2356 => '0',
		2357 => '0',
		2358 => '0',
		2359 => '0',
		2360 => '0',
		2361 => '0',
		2362 => '0',
		2363 => '0',
		2364 => '0',
		2365 => '0',
		2366 => '0',
		2367 => '0',
		2368 => '0',
		2369 => '0',
		2370 => '0',
		2371 => '0',
		2372 => '0',
		2373 => '0',
		2374 => '0',
		2375 => '0',
		2376 => '0',
		2377 => '0',
		2378 => '0',
		2379 => '0',
		2380 => '0',
		2381 => '0',
		2382 => '0',
		2383 => '0',
		2384 => '0',
		2385 => '0',
		2386 => '0',
		2387 => '0',
		2388 => '0',
		2389 => '0',
		2390 => '0',
		2391 => '0',
		2392 => '0',
		2393 => '0',
		2394 => '0',
		2395 => '0',
		2396 => '0',
		2397 => '0',
		2398 => '0',
		2399 => '0',
		2400 => '0',
		2401 => '0',
		2402 => '0',
		2403 => '0',
		2404 => '0',
		2405 => '0',
		2406 => '0',
		2407 => '0',
		2408 => '0',
		2409 => '0',
		2410 => '0',
		2411 => '0',
		2412 => '0',
		2413 => '0',
		2414 => '0',
		2415 => '0',
		2416 => '0',
		2417 => '0',
		2418 => '0',
		2419 => '0',
		2420 => '0',
		2421 => '0',
		2422 => '0',
		2423 => '0',
		2432 => '0',
		2433 => '0',
		2434 => '0',
		2435 => '0',
		2436 => '0',
		2437 => '0',
		2438 => '0',
		2439 => '0',
		2440 => '0',
		2441 => '0',
		2442 => '0',
		2443 => '0',
		2444 => '0',
		2445 => '0',
		2446 => '0',
		2447 => '0',
		2448 => '0',
		2449 => '0',
		2450 => '0',
		2451 => '0',
		2452 => '0',
		2453 => '0',
		2454 => '0',
		2455 => '0',
		2456 => '0',
		2457 => '0',
		2458 => '0',
		2459 => '0',
		2460 => '0',
		2461 => '0',
		2462 => '0',
		2463 => '0',
		2464 => '0',
		2465 => '0',
		2466 => '0',
		2467 => '0',
		2468 => '0',
		2469 => '0',
		2470 => '0',
		2471 => '0',
		2472 => '0',
		2473 => '0',
		2474 => '0',
		2475 => '0',
		2476 => '0',
		2477 => '0',
		2478 => '0',
		2479 => '0',
		2480 => '0',
		2481 => '0',
		2482 => '0',
		2483 => '0',
		2484 => '0',
		2485 => '0',
		2486 => '0',
		2487 => '0',
		2488 => '0',
		2489 => '0',
		2490 => '0',
		2491 => '0',
		2492 => '0',
		2493 => '0',
		2494 => '0',
		2495 => '0',
		2496 => '0',
		2497 => '0',
		2498 => '0',
		2499 => '0',
		2500 => '0',
		2501 => '0',
		2502 => '0',
		2503 => '0',
		2504 => '0',
		2505 => '0',
		2506 => '0',
		2507 => '0',
		2508 => '0',
		2509 => '0',
		2510 => '0',
		2511 => '0',
		2512 => '0',
		2513 => '0',
		2514 => '0',
		2515 => '0',
		2516 => '0',
		2517 => '0',
		2518 => '0',
		2519 => '0',
		2520 => '0',
		2521 => '0',
		2522 => '0',
		2523 => '0',
		2524 => '0',
		2525 => '0',
		2526 => '0',
		2527 => '0',
		2528 => '0',
		2529 => '0',
		2530 => '0',
		2531 => '0',
		2532 => '0',
		2533 => '0',
		2534 => '0',
		2535 => '0',
		2536 => '0',
		2537 => '0',
		2538 => '0',
		2539 => '0',
		2540 => '0',
		2541 => '0',
		2542 => '0',
		2543 => '0',
		2544 => '0',
		2545 => '0',
		2546 => '0',
		2547 => '0',
		2548 => '0',
		2549 => '0',
		2550 => '0',
		2551 => '0',
		2560 => '0',
		2561 => '0',
		2562 => '0',
		2563 => '0',
		2564 => '0',
		2565 => '0',
		2566 => '0',
		2567 => '0',
		2568 => '0',
		2569 => '0',
		2570 => '0',
		2571 => '0',
		2572 => '0',
		2573 => '0',
		2574 => '0',
		2575 => '0',
		2576 => '0',
		2577 => '0',
		2578 => '0',
		2579 => '0',
		2580 => '0',
		2581 => '0',
		2582 => '0',
		2583 => '0',
		2584 => '0',
		2585 => '0',
		2586 => '0',
		2587 => '0',
		2588 => '0',
		2589 => '0',
		2590 => '0',
		2591 => '0',
		2592 => '0',
		2593 => '0',
		2594 => '0',
		2595 => '0',
		2596 => '0',
		2597 => '0',
		2598 => '0',
		2599 => '0',
		2600 => '0',
		2601 => '0',
		2602 => '0',
		2603 => '0',
		2604 => '0',
		2605 => '0',
		2606 => '0',
		2607 => '0',
		2608 => '0',
		2609 => '0',
		2610 => '0',
		2611 => '0',
		2612 => '0',
		2613 => '0',
		2614 => '0',
		2615 => '0',
		2616 => '0',
		2617 => '0',
		2618 => '0',
		2619 => '0',
		2620 => '0',
		2621 => '0',
		2622 => '0',
		2623 => '0',
		2624 => '0',
		2625 => '0',
		2626 => '0',
		2627 => '0',
		2628 => '0',
		2629 => '0',
		2630 => '0',
		2631 => '0',
		2632 => '0',
		2633 => '0',
		2634 => '0',
		2635 => '0',
		2636 => '0',
		2637 => '0',
		2638 => '0',
		2639 => '0',
		2640 => '0',
		2641 => '0',
		2642 => '0',
		2643 => '0',
		2644 => '0',
		2645 => '0',
		2646 => '0',
		2647 => '0',
		2648 => '0',
		2649 => '0',
		2650 => '0',
		2651 => '0',
		2652 => '0',
		2653 => '0',
		2654 => '0',
		2655 => '0',
		2656 => '0',
		2657 => '0',
		2658 => '0',
		2659 => '0',
		2660 => '0',
		2661 => '0',
		2662 => '0',
		2663 => '0',
		2664 => '0',
		2665 => '0',
		2666 => '0',
		2667 => '0',
		2668 => '0',
		2669 => '0',
		2670 => '0',
		2671 => '0',
		2672 => '0',
		2673 => '0',
		2674 => '0',
		2675 => '0',
		2676 => '0',
		2677 => '0',
		2678 => '0',
		2679 => '0',
		2688 => '0',
		2689 => '0',
		2690 => '0',
		2691 => '0',
		2692 => '0',
		2693 => '0',
		2694 => '0',
		2695 => '0',
		2696 => '0',
		2697 => '0',
		2698 => '0',
		2699 => '0',
		2700 => '0',
		2701 => '0',
		2702 => '0',
		2703 => '0',
		2704 => '0',
		2705 => '0',
		2706 => '0',
		2707 => '0',
		2708 => '0',
		2709 => '0',
		2710 => '0',
		2711 => '0',
		2712 => '0',
		2713 => '0',
		2714 => '0',
		2715 => '0',
		2716 => '0',
		2717 => '0',
		2718 => '0',
		2719 => '0',
		2720 => '0',
		2721 => '0',
		2722 => '0',
		2723 => '0',
		2724 => '0',
		2725 => '0',
		2726 => '0',
		2727 => '0',
		2728 => '0',
		2729 => '0',
		2730 => '0',
		2731 => '0',
		2732 => '0',
		2733 => '0',
		2734 => '0',
		2735 => '0',
		2736 => '0',
		2737 => '0',
		2738 => '0',
		2739 => '0',
		2740 => '0',
		2741 => '0',
		2742 => '0',
		2743 => '0',
		2744 => '0',
		2745 => '0',
		2746 => '0',
		2747 => '0',
		2748 => '0',
		2749 => '0',
		2750 => '0',
		2751 => '0',
		2752 => '0',
		2753 => '0',
		2754 => '0',
		2755 => '0',
		2756 => '0',
		2757 => '0',
		2758 => '0',
		2759 => '0',
		2760 => '0',
		2761 => '0',
		2762 => '0',
		2763 => '0',
		2764 => '0',
		2765 => '0',
		2766 => '0',
		2767 => '0',
		2768 => '0',
		2769 => '0',
		2770 => '0',
		2771 => '0',
		2772 => '0',
		2773 => '0',
		2774 => '0',
		2775 => '0',
		2776 => '0',
		2777 => '0',
		2778 => '0',
		2779 => '0',
		2780 => '0',
		2781 => '0',
		2782 => '0',
		2783 => '0',
		2784 => '0',
		2785 => '0',
		2786 => '0',
		2787 => '0',
		2788 => '0',
		2789 => '0',
		2790 => '0',
		2791 => '0',
		2792 => '0',
		2793 => '0',
		2794 => '0',
		2795 => '0',
		2796 => '0',
		2797 => '0',
		2798 => '0',
		2799 => '0',
		2800 => '0',
		2801 => '0',
		2802 => '0',
		2803 => '0',
		2804 => '0',
		2805 => '0',
		2806 => '0',
		2807 => '0',
		2816 => '0',
		2817 => '0',
		2818 => '0',
		2819 => '0',
		2820 => '0',
		2821 => '0',
		2822 => '0',
		2823 => '0',
		2824 => '0',
		2825 => '0',
		2826 => '0',
		2827 => '0',
		2828 => '0',
		2829 => '0',
		2830 => '0',
		2831 => '0',
		2832 => '0',
		2833 => '0',
		2834 => '0',
		2835 => '0',
		2836 => '0',
		2837 => '0',
		2838 => '0',
		2839 => '0',
		2840 => '0',
		2841 => '0',
		2842 => '0',
		2843 => '0',
		2844 => '0',
		2845 => '0',
		2846 => '0',
		2847 => '0',
		2848 => '0',
		2849 => '0',
		2850 => '0',
		2851 => '0',
		2852 => '0',
		2853 => '0',
		2854 => '0',
		2855 => '0',
		2856 => '0',
		2857 => '0',
		2858 => '0',
		2859 => '0',
		2860 => '0',
		2861 => '0',
		2862 => '0',
		2863 => '0',
		2864 => '0',
		2865 => '0',
		2866 => '0',
		2867 => '0',
		2868 => '0',
		2869 => '0',
		2870 => '0',
		2871 => '0',
		2872 => '0',
		2873 => '0',
		2874 => '0',
		2875 => '0',
		2876 => '0',
		2877 => '0',
		2878 => '0',
		2879 => '0',
		2880 => '0',
		2881 => '0',
		2882 => '0',
		2883 => '0',
		2884 => '0',
		2885 => '0',
		2886 => '0',
		2887 => '0',
		2888 => '0',
		2889 => '0',
		2890 => '0',
		2891 => '0',
		2892 => '0',
		2893 => '0',
		2894 => '0',
		2895 => '0',
		2896 => '0',
		2897 => '0',
		2898 => '0',
		2899 => '0',
		2900 => '0',
		2901 => '0',
		2902 => '0',
		2903 => '0',
		2904 => '0',
		2905 => '0',
		2906 => '0',
		2907 => '0',
		2908 => '0',
		2909 => '0',
		2910 => '0',
		2911 => '0',
		2912 => '0',
		2913 => '0',
		2914 => '0',
		2915 => '0',
		2916 => '0',
		2917 => '0',
		2918 => '0',
		2919 => '0',
		2920 => '0',
		2921 => '0',
		2922 => '0',
		2923 => '0',
		2924 => '0',
		2925 => '0',
		2926 => '0',
		2927 => '0',
		2928 => '0',
		2929 => '0',
		2930 => '0',
		2931 => '0',
		2932 => '0',
		2933 => '0',
		2934 => '0',
		2935 => '0',
		2944 => '0',
		2945 => '0',
		2946 => '0',
		2947 => '0',
		2948 => '0',
		2949 => '0',
		2950 => '0',
		2951 => '0',
		2952 => '0',
		2953 => '0',
		2954 => '0',
		2955 => '0',
		2956 => '0',
		2957 => '0',
		2958 => '0',
		2959 => '0',
		2960 => '0',
		2961 => '0',
		2962 => '0',
		2963 => '0',
		2964 => '0',
		2965 => '0',
		2966 => '0',
		2967 => '0',
		2968 => '0',
		2969 => '0',
		2970 => '0',
		2971 => '0',
		2972 => '0',
		2973 => '0',
		2974 => '0',
		2975 => '0',
		2976 => '0',
		2977 => '0',
		2978 => '0',
		2979 => '0',
		2980 => '0',
		2981 => '0',
		2982 => '0',
		2983 => '0',
		2984 => '0',
		2985 => '0',
		2986 => '0',
		2987 => '0',
		2988 => '0',
		2989 => '0',
		2990 => '0',
		2991 => '0',
		2992 => '0',
		2993 => '0',
		2994 => '0',
		2995 => '0',
		2996 => '0',
		2997 => '0',
		2998 => '0',
		2999 => '0',
		3000 => '0',
		3001 => '0',
		3002 => '0',
		3003 => '0',
		3004 => '0',
		3005 => '0',
		3006 => '0',
		3007 => '0',
		3008 => '0',
		3009 => '0',
		3010 => '0',
		3011 => '0',
		3012 => '0',
		3013 => '0',
		3014 => '0',
		3015 => '0',
		3016 => '0',
		3017 => '0',
		3018 => '0',
		3019 => '0',
		3020 => '0',
		3021 => '0',
		3022 => '0',
		3023 => '0',
		3024 => '0',
		3025 => '0',
		3026 => '0',
		3027 => '0',
		3028 => '0',
		3029 => '0',
		3030 => '0',
		3031 => '0',
		3032 => '0',
		3033 => '0',
		3034 => '0',
		3035 => '0',
		3036 => '0',
		3037 => '0',
		3038 => '0',
		3039 => '0',
		3040 => '0',
		3041 => '0',
		3042 => '0',
		3043 => '0',
		3044 => '0',
		3045 => '0',
		3046 => '0',
		3047 => '0',
		3048 => '0',
		3049 => '0',
		3050 => '0',
		3051 => '0',
		3052 => '0',
		3053 => '0',
		3054 => '0',
		3055 => '0',
		3056 => '0',
		3057 => '0',
		3058 => '0',
		3059 => '0',
		3060 => '0',
		3061 => '0',
		3062 => '0',
		3063 => '0',
		3072 => '1',
		3073 => '1',
		3074 => '1',
		3075 => '1',
		3076 => '1',
		3077 => '1',
		3078 => '1',
		3079 => '1',
		3080 => '1',
		3081 => '1',
		3082 => '1',
		3083 => '1',
		3084 => '1',
		3085 => '0',
		3086 => '0',
		3087 => '1',
		3088 => '1',
		3089 => '1',
		3090 => '1',
		3091 => '1',
		3092 => '1',
		3093 => '1',
		3094 => '1',
		3095 => '0',
		3096 => '0',
		3097 => '1',
		3098 => '1',
		3099 => '1',
		3100 => '1',
		3101 => '1',
		3102 => '1',
		3103 => '1',
		3104 => '1',
		3105 => '1',
		3106 => '1',
		3107 => '1',
		3108 => '1',
		3109 => '1',
		3110 => '0',
		3111 => '0',
		3112 => '1',
		3113 => '1',
		3114 => '1',
		3115 => '1',
		3116 => '1',
		3117 => '1',
		3118 => '1',
		3119 => '1',
		3120 => '1',
		3121 => '1',
		3122 => '1',
		3123 => '1',
		3124 => '1',
		3125 => '0',
		3126 => '0',
		3127 => '1',
		3128 => '1',
		3129 => '1',
		3130 => '1',
		3131 => '1',
		3132 => '1',
		3133 => '1',
		3134 => '1',
		3135 => '1',
		3136 => '1',
		3137 => '1',
		3138 => '1',
		3139 => '1',
		3140 => '0',
		3141 => '0',
		3142 => '1',
		3143 => '1',
		3144 => '1',
		3145 => '1',
		3146 => '1',
		3147 => '1',
		3148 => '1',
		3149 => '1',
		3150 => '0',
		3151 => '0',
		3152 => '1',
		3153 => '1',
		3154 => '1',
		3155 => '1',
		3156 => '1',
		3157 => '1',
		3158 => '1',
		3159 => '1',
		3160 => '1',
		3161 => '1',
		3162 => '1',
		3163 => '1',
		3164 => '1',
		3165 => '0',
		3166 => '0',
		3167 => '1',
		3168 => '1',
		3169 => '1',
		3170 => '1',
		3171 => '1',
		3172 => '1',
		3173 => '1',
		3174 => '1',
		3175 => '1',
		3176 => '1',
		3177 => '1',
		3178 => '1',
		3179 => '1',
		3180 => '0',
		3181 => '0',
		3182 => '1',
		3183 => '1',
		3184 => '1',
		3185 => '1',
		3186 => '1',
		3187 => '1',
		3188 => '1',
		3189 => '1',
		3190 => '0',
		3191 => '0',
		3200 => '1',
		3201 => '1',
		3202 => '1',
		3203 => '1',
		3204 => '1',
		3205 => '1',
		3206 => '1',
		3207 => '1',
		3208 => '1',
		3209 => '1',
		3210 => '1',
		3211 => '1',
		3212 => '1',
		3213 => '0',
		3214 => '0',
		3215 => '1',
		3216 => '1',
		3217 => '1',
		3218 => '1',
		3219 => '1',
		3220 => '1',
		3221 => '1',
		3222 => '1',
		3223 => '0',
		3224 => '0',
		3225 => '1',
		3226 => '1',
		3227 => '1',
		3228 => '1',
		3229 => '1',
		3230 => '1',
		3231 => '1',
		3232 => '1',
		3233 => '1',
		3234 => '1',
		3235 => '1',
		3236 => '1',
		3237 => '1',
		3238 => '0',
		3239 => '0',
		3240 => '1',
		3241 => '1',
		3242 => '1',
		3243 => '1',
		3244 => '1',
		3245 => '1',
		3246 => '1',
		3247 => '1',
		3248 => '1',
		3249 => '1',
		3250 => '1',
		3251 => '1',
		3252 => '1',
		3253 => '0',
		3254 => '0',
		3255 => '1',
		3256 => '1',
		3257 => '1',
		3258 => '1',
		3259 => '1',
		3260 => '1',
		3261 => '1',
		3262 => '1',
		3263 => '1',
		3264 => '1',
		3265 => '1',
		3266 => '1',
		3267 => '1',
		3268 => '0',
		3269 => '0',
		3270 => '1',
		3271 => '1',
		3272 => '1',
		3273 => '1',
		3274 => '1',
		3275 => '1',
		3276 => '1',
		3277 => '1',
		3278 => '0',
		3279 => '0',
		3280 => '1',
		3281 => '1',
		3282 => '1',
		3283 => '1',
		3284 => '1',
		3285 => '1',
		3286 => '1',
		3287 => '1',
		3288 => '1',
		3289 => '1',
		3290 => '1',
		3291 => '1',
		3292 => '1',
		3293 => '0',
		3294 => '0',
		3295 => '1',
		3296 => '1',
		3297 => '1',
		3298 => '1',
		3299 => '1',
		3300 => '1',
		3301 => '1',
		3302 => '1',
		3303 => '1',
		3304 => '1',
		3305 => '1',
		3306 => '1',
		3307 => '1',
		3308 => '0',
		3309 => '0',
		3310 => '1',
		3311 => '1',
		3312 => '1',
		3313 => '1',
		3314 => '1',
		3315 => '1',
		3316 => '1',
		3317 => '1',
		3318 => '0',
		3319 => '0',
		3328 => '1',
		3329 => '1',
		3330 => '1',
		3331 => '1',
		3332 => '1',
		3333 => '1',
		3334 => '1',
		3335 => '1',
		3336 => '1',
		3337 => '1',
		3338 => '1',
		3339 => '1',
		3340 => '1',
		3341 => '0',
		3342 => '0',
		3343 => '1',
		3344 => '1',
		3345 => '1',
		3346 => '1',
		3347 => '1',
		3348 => '1',
		3349 => '1',
		3350 => '1',
		3351 => '0',
		3352 => '0',
		3353 => '1',
		3354 => '1',
		3355 => '1',
		3356 => '1',
		3357 => '1',
		3358 => '1',
		3359 => '1',
		3360 => '1',
		3361 => '1',
		3362 => '1',
		3363 => '1',
		3364 => '1',
		3365 => '1',
		3366 => '0',
		3367 => '0',
		3368 => '1',
		3369 => '1',
		3370 => '1',
		3371 => '1',
		3372 => '1',
		3373 => '1',
		3374 => '1',
		3375 => '1',
		3376 => '1',
		3377 => '1',
		3378 => '1',
		3379 => '1',
		3380 => '1',
		3381 => '0',
		3382 => '0',
		3383 => '1',
		3384 => '1',
		3385 => '1',
		3386 => '1',
		3387 => '1',
		3388 => '1',
		3389 => '1',
		3390 => '1',
		3391 => '1',
		3392 => '1',
		3393 => '1',
		3394 => '1',
		3395 => '1',
		3396 => '0',
		3397 => '0',
		3398 => '1',
		3399 => '1',
		3400 => '1',
		3401 => '1',
		3402 => '1',
		3403 => '1',
		3404 => '1',
		3405 => '1',
		3406 => '0',
		3407 => '0',
		3408 => '1',
		3409 => '1',
		3410 => '1',
		3411 => '1',
		3412 => '1',
		3413 => '1',
		3414 => '1',
		3415 => '1',
		3416 => '1',
		3417 => '1',
		3418 => '1',
		3419 => '1',
		3420 => '1',
		3421 => '0',
		3422 => '0',
		3423 => '1',
		3424 => '1',
		3425 => '1',
		3426 => '1',
		3427 => '1',
		3428 => '1',
		3429 => '1',
		3430 => '1',
		3431 => '1',
		3432 => '1',
		3433 => '1',
		3434 => '1',
		3435 => '1',
		3436 => '0',
		3437 => '0',
		3438 => '1',
		3439 => '1',
		3440 => '1',
		3441 => '1',
		3442 => '1',
		3443 => '1',
		3444 => '1',
		3445 => '1',
		3446 => '0',
		3447 => '0',
		3456 => '1',
		3457 => '1',
		3458 => '1',
		3459 => '0',
		3460 => '0',
		3461 => '1',
		3462 => '1',
		3463 => '1',
		3464 => '0',
		3465 => '0',
		3466 => '1',
		3467 => '1',
		3468 => '1',
		3469 => '0',
		3470 => '0',
		3471 => '1',
		3472 => '1',
		3473 => '1',
		3474 => '0',
		3475 => '0',
		3476 => '1',
		3477 => '1',
		3478 => '1',
		3479 => '0',
		3480 => '0',
		3481 => '1',
		3482 => '1',
		3483 => '1',
		3484 => '0',
		3485 => '0',
		3486 => '0',
		3487 => '0',
		3488 => '0',
		3489 => '0',
		3490 => '0',
		3491 => '1',
		3492 => '1',
		3493 => '1',
		3494 => '0',
		3495 => '0',
		3496 => '1',
		3497 => '1',
		3498 => '1',
		3499 => '0',
		3500 => '0',
		3501 => '0',
		3502 => '0',
		3503 => '0',
		3504 => '0',
		3505 => '0',
		3506 => '1',
		3507 => '1',
		3508 => '1',
		3509 => '0',
		3510 => '0',
		3511 => '1',
		3512 => '1',
		3513 => '1',
		3514 => '0',
		3515 => '0',
		3516 => '0',
		3517 => '0',
		3518 => '0',
		3519 => '0',
		3520 => '0',
		3521 => '1',
		3522 => '1',
		3523 => '1',
		3524 => '0',
		3525 => '0',
		3526 => '1',
		3527 => '1',
		3528 => '1',
		3529 => '0',
		3530 => '0',
		3531 => '1',
		3532 => '1',
		3533 => '1',
		3534 => '0',
		3535 => '0',
		3536 => '1',
		3537 => '1',
		3538 => '1',
		3539 => '0',
		3540 => '0',
		3541 => '0',
		3542 => '0',
		3543 => '0',
		3544 => '0',
		3545 => '0',
		3546 => '1',
		3547 => '1',
		3548 => '1',
		3549 => '0',
		3550 => '0',
		3551 => '1',
		3552 => '1',
		3553 => '1',
		3554 => '0',
		3555 => '0',
		3556 => '0',
		3557 => '0',
		3558 => '0',
		3559 => '0',
		3560 => '0',
		3561 => '1',
		3562 => '1',
		3563 => '1',
		3564 => '0',
		3565 => '0',
		3566 => '1',
		3567 => '1',
		3568 => '1',
		3569 => '0',
		3570 => '0',
		3571 => '1',
		3572 => '1',
		3573 => '1',
		3574 => '0',
		3575 => '0',
		3584 => '1',
		3585 => '1',
		3586 => '1',
		3587 => '0',
		3588 => '0',
		3589 => '1',
		3590 => '1',
		3591 => '1',
		3592 => '0',
		3593 => '0',
		3594 => '1',
		3595 => '1',
		3596 => '1',
		3597 => '0',
		3598 => '0',
		3599 => '1',
		3600 => '1',
		3601 => '1',
		3602 => '0',
		3603 => '0',
		3604 => '1',
		3605 => '1',
		3606 => '1',
		3607 => '0',
		3608 => '0',
		3609 => '1',
		3610 => '1',
		3611 => '1',
		3612 => '0',
		3613 => '0',
		3614 => '0',
		3615 => '0',
		3616 => '0',
		3617 => '0',
		3618 => '0',
		3619 => '1',
		3620 => '1',
		3621 => '1',
		3622 => '0',
		3623 => '0',
		3624 => '1',
		3625 => '1',
		3626 => '1',
		3627 => '0',
		3628 => '0',
		3629 => '0',
		3630 => '0',
		3631 => '0',
		3632 => '0',
		3633 => '0',
		3634 => '1',
		3635 => '1',
		3636 => '1',
		3637 => '0',
		3638 => '0',
		3639 => '1',
		3640 => '1',
		3641 => '1',
		3642 => '0',
		3643 => '0',
		3644 => '0',
		3645 => '0',
		3646 => '0',
		3647 => '0',
		3648 => '0',
		3649 => '1',
		3650 => '1',
		3651 => '1',
		3652 => '0',
		3653 => '0',
		3654 => '1',
		3655 => '1',
		3656 => '1',
		3657 => '0',
		3658 => '0',
		3659 => '1',
		3660 => '1',
		3661 => '1',
		3662 => '0',
		3663 => '0',
		3664 => '1',
		3665 => '1',
		3666 => '1',
		3667 => '0',
		3668 => '0',
		3669 => '0',
		3670 => '0',
		3671 => '0',
		3672 => '0',
		3673 => '0',
		3674 => '1',
		3675 => '1',
		3676 => '1',
		3677 => '0',
		3678 => '0',
		3679 => '1',
		3680 => '1',
		3681 => '1',
		3682 => '0',
		3683 => '0',
		3684 => '0',
		3685 => '0',
		3686 => '0',
		3687 => '0',
		3688 => '0',
		3689 => '1',
		3690 => '1',
		3691 => '1',
		3692 => '0',
		3693 => '0',
		3694 => '1',
		3695 => '1',
		3696 => '1',
		3697 => '0',
		3698 => '0',
		3699 => '1',
		3700 => '1',
		3701 => '1',
		3702 => '0',
		3703 => '0',
		3712 => '1',
		3713 => '1',
		3714 => '1',
		3715 => '0',
		3716 => '0',
		3717 => '1',
		3718 => '1',
		3719 => '1',
		3720 => '0',
		3721 => '0',
		3722 => '1',
		3723 => '1',
		3724 => '1',
		3725 => '0',
		3726 => '0',
		3727 => '1',
		3728 => '1',
		3729 => '1',
		3730 => '0',
		3731 => '0',
		3732 => '1',
		3733 => '1',
		3734 => '1',
		3735 => '0',
		3736 => '0',
		3737 => '1',
		3738 => '1',
		3739 => '1',
		3740 => '0',
		3741 => '0',
		3742 => '0',
		3743 => '0',
		3744 => '0',
		3745 => '0',
		3746 => '0',
		3747 => '1',
		3748 => '1',
		3749 => '1',
		3750 => '0',
		3751 => '0',
		3752 => '1',
		3753 => '1',
		3754 => '1',
		3755 => '1',
		3756 => '1',
		3757 => '1',
		3758 => '0',
		3759 => '1',
		3760 => '1',
		3761 => '1',
		3762 => '1',
		3763 => '1',
		3764 => '1',
		3765 => '0',
		3766 => '0',
		3767 => '1',
		3768 => '1',
		3769 => '1',
		3770 => '0',
		3771 => '0',
		3772 => '0',
		3773 => '0',
		3774 => '0',
		3775 => '0',
		3776 => '0',
		3777 => '1',
		3778 => '1',
		3779 => '1',
		3780 => '0',
		3781 => '0',
		3782 => '1',
		3783 => '1',
		3784 => '1',
		3785 => '0',
		3786 => '0',
		3787 => '1',
		3788 => '1',
		3789 => '1',
		3790 => '0',
		3791 => '0',
		3792 => '1',
		3793 => '1',
		3794 => '1',
		3795 => '0',
		3796 => '0',
		3797 => '1',
		3798 => '1',
		3799 => '1',
		3800 => '0',
		3801 => '0',
		3802 => '1',
		3803 => '1',
		3804 => '1',
		3805 => '0',
		3806 => '0',
		3807 => '1',
		3808 => '1',
		3809 => '1',
		3810 => '0',
		3811 => '0',
		3812 => '1',
		3813 => '1',
		3814 => '1',
		3815 => '1',
		3816 => '1',
		3817 => '1',
		3818 => '1',
		3819 => '1',
		3820 => '0',
		3821 => '0',
		3822 => '1',
		3823 => '1',
		3824 => '1',
		3825 => '0',
		3826 => '0',
		3827 => '1',
		3828 => '1',
		3829 => '1',
		3830 => '0',
		3831 => '0',
		3840 => '1',
		3841 => '1',
		3842 => '1',
		3843 => '0',
		3844 => '0',
		3845 => '1',
		3846 => '1',
		3847 => '1',
		3848 => '0',
		3849 => '0',
		3850 => '1',
		3851 => '1',
		3852 => '1',
		3853 => '0',
		3854 => '0',
		3855 => '1',
		3856 => '1',
		3857 => '1',
		3858 => '0',
		3859 => '0',
		3860 => '1',
		3861 => '1',
		3862 => '1',
		3863 => '0',
		3864 => '0',
		3865 => '1',
		3866 => '1',
		3867 => '1',
		3868 => '0',
		3869 => '0',
		3870 => '1',
		3871 => '1',
		3872 => '1',
		3873 => '0',
		3874 => '0',
		3875 => '1',
		3876 => '1',
		3877 => '1',
		3878 => '0',
		3879 => '0',
		3880 => '1',
		3881 => '1',
		3882 => '1',
		3883 => '1',
		3884 => '1',
		3885 => '1',
		3886 => '0',
		3887 => '1',
		3888 => '1',
		3889 => '1',
		3890 => '1',
		3891 => '1',
		3892 => '1',
		3893 => '0',
		3894 => '0',
		3895 => '1',
		3896 => '1',
		3897 => '1',
		3898 => '0',
		3899 => '0',
		3900 => '1',
		3901 => '1',
		3902 => '1',
		3903 => '0',
		3904 => '0',
		3905 => '1',
		3906 => '1',
		3907 => '1',
		3908 => '0',
		3909 => '0',
		3910 => '1',
		3911 => '1',
		3912 => '1',
		3913 => '0',
		3914 => '0',
		3915 => '1',
		3916 => '1',
		3917 => '1',
		3918 => '0',
		3919 => '0',
		3920 => '1',
		3921 => '1',
		3922 => '1',
		3923 => '0',
		3924 => '0',
		3925 => '1',
		3926 => '1',
		3927 => '1',
		3928 => '0',
		3929 => '0',
		3930 => '1',
		3931 => '1',
		3932 => '1',
		3933 => '0',
		3934 => '0',
		3935 => '1',
		3936 => '1',
		3937 => '1',
		3938 => '0',
		3939 => '0',
		3940 => '1',
		3941 => '1',
		3942 => '1',
		3943 => '1',
		3944 => '1',
		3945 => '1',
		3946 => '1',
		3947 => '1',
		3948 => '0',
		3949 => '0',
		3950 => '1',
		3951 => '1',
		3952 => '1',
		3953 => '0',
		3954 => '0',
		3955 => '1',
		3956 => '1',
		3957 => '1',
		3958 => '0',
		3959 => '0',
		3968 => '1',
		3969 => '1',
		3970 => '1',
		3971 => '0',
		3972 => '0',
		3973 => '1',
		3974 => '1',
		3975 => '1',
		3976 => '0',
		3977 => '0',
		3978 => '1',
		3979 => '1',
		3980 => '1',
		3981 => '0',
		3982 => '0',
		3983 => '1',
		3984 => '1',
		3985 => '1',
		3986 => '0',
		3987 => '0',
		3988 => '1',
		3989 => '1',
		3990 => '1',
		3991 => '0',
		3992 => '0',
		3993 => '1',
		3994 => '1',
		3995 => '1',
		3996 => '0',
		3997 => '0',
		3998 => '1',
		3999 => '1',
		4000 => '1',
		4001 => '0',
		4002 => '0',
		4003 => '1',
		4004 => '1',
		4005 => '1',
		4006 => '0',
		4007 => '0',
		4008 => '1',
		4009 => '1',
		4010 => '1',
		4011 => '1',
		4012 => '1',
		4013 => '1',
		4014 => '0',
		4015 => '1',
		4016 => '1',
		4017 => '1',
		4018 => '1',
		4019 => '1',
		4020 => '1',
		4021 => '0',
		4022 => '0',
		4023 => '1',
		4024 => '1',
		4025 => '1',
		4026 => '0',
		4027 => '0',
		4028 => '1',
		4029 => '1',
		4030 => '1',
		4031 => '0',
		4032 => '0',
		4033 => '1',
		4034 => '1',
		4035 => '1',
		4036 => '0',
		4037 => '0',
		4038 => '1',
		4039 => '1',
		4040 => '1',
		4041 => '0',
		4042 => '0',
		4043 => '1',
		4044 => '1',
		4045 => '1',
		4046 => '0',
		4047 => '0',
		4048 => '1',
		4049 => '1',
		4050 => '1',
		4051 => '0',
		4052 => '0',
		4053 => '1',
		4054 => '1',
		4055 => '1',
		4056 => '0',
		4057 => '0',
		4058 => '1',
		4059 => '1',
		4060 => '1',
		4061 => '0',
		4062 => '0',
		4063 => '1',
		4064 => '1',
		4065 => '1',
		4066 => '0',
		4067 => '0',
		4068 => '1',
		4069 => '1',
		4070 => '1',
		4071 => '1',
		4072 => '1',
		4073 => '1',
		4074 => '1',
		4075 => '1',
		4076 => '0',
		4077 => '0',
		4078 => '1',
		4079 => '1',
		4080 => '1',
		4081 => '0',
		4082 => '0',
		4083 => '1',
		4084 => '1',
		4085 => '1',
		4086 => '0',
		4087 => '0',
		4096 => '1',
		4097 => '1',
		4098 => '1',
		4099 => '0',
		4100 => '0',
		4101 => '1',
		4102 => '1',
		4103 => '1',
		4104 => '0',
		4105 => '0',
		4106 => '1',
		4107 => '1',
		4108 => '1',
		4109 => '0',
		4110 => '0',
		4111 => '1',
		4112 => '1',
		4113 => '1',
		4114 => '0',
		4115 => '0',
		4116 => '1',
		4117 => '1',
		4118 => '1',
		4119 => '0',
		4120 => '0',
		4121 => '1',
		4122 => '1',
		4123 => '1',
		4124 => '0',
		4125 => '0',
		4126 => '1',
		4127 => '1',
		4128 => '1',
		4129 => '1',
		4130 => '1',
		4131 => '1',
		4132 => '1',
		4133 => '1',
		4134 => '0',
		4135 => '0',
		4136 => '0',
		4137 => '0',
		4138 => '0',
		4139 => '1',
		4140 => '1',
		4141 => '1',
		4142 => '0',
		4143 => '1',
		4144 => '1',
		4145 => '1',
		4146 => '0',
		4147 => '0',
		4148 => '0',
		4149 => '0',
		4150 => '0',
		4151 => '1',
		4152 => '1',
		4153 => '1',
		4154 => '0',
		4155 => '0',
		4156 => '1',
		4157 => '1',
		4158 => '1',
		4159 => '0',
		4160 => '0',
		4161 => '1',
		4162 => '1',
		4163 => '1',
		4164 => '0',
		4165 => '0',
		4166 => '1',
		4167 => '1',
		4168 => '1',
		4169 => '0',
		4170 => '0',
		4171 => '1',
		4172 => '1',
		4173 => '1',
		4174 => '0',
		4175 => '0',
		4176 => '1',
		4177 => '1',
		4178 => '1',
		4179 => '0',
		4180 => '0',
		4181 => '0',
		4182 => '0',
		4183 => '0',
		4184 => '1',
		4185 => '1',
		4186 => '1',
		4187 => '1',
		4188 => '1',
		4189 => '0',
		4190 => '0',
		4191 => '1',
		4192 => '1',
		4193 => '1',
		4194 => '0',
		4195 => '0',
		4196 => '0',
		4197 => '0',
		4198 => '0',
		4199 => '0',
		4200 => '0',
		4201 => '1',
		4202 => '1',
		4203 => '1',
		4204 => '0',
		4205 => '0',
		4206 => '1',
		4207 => '1',
		4208 => '1',
		4209 => '0',
		4210 => '0',
		4211 => '1',
		4212 => '1',
		4213 => '1',
		4214 => '0',
		4215 => '0',
		4224 => '1',
		4225 => '1',
		4226 => '1',
		4227 => '0',
		4228 => '0',
		4229 => '1',
		4230 => '1',
		4231 => '1',
		4232 => '0',
		4233 => '0',
		4234 => '1',
		4235 => '1',
		4236 => '1',
		4237 => '0',
		4238 => '0',
		4239 => '1',
		4240 => '1',
		4241 => '1',
		4242 => '0',
		4243 => '0',
		4244 => '1',
		4245 => '1',
		4246 => '1',
		4247 => '0',
		4248 => '0',
		4249 => '1',
		4250 => '1',
		4251 => '1',
		4252 => '0',
		4253 => '0',
		4254 => '1',
		4255 => '1',
		4256 => '1',
		4257 => '1',
		4258 => '1',
		4259 => '1',
		4260 => '1',
		4261 => '1',
		4262 => '0',
		4263 => '0',
		4264 => '0',
		4265 => '0',
		4266 => '0',
		4267 => '1',
		4268 => '1',
		4269 => '1',
		4270 => '0',
		4271 => '1',
		4272 => '1',
		4273 => '1',
		4274 => '0',
		4275 => '0',
		4276 => '0',
		4277 => '0',
		4278 => '0',
		4279 => '1',
		4280 => '1',
		4281 => '1',
		4282 => '0',
		4283 => '0',
		4284 => '1',
		4285 => '1',
		4286 => '1',
		4287 => '0',
		4288 => '0',
		4289 => '1',
		4290 => '1',
		4291 => '1',
		4292 => '0',
		4293 => '0',
		4294 => '1',
		4295 => '1',
		4296 => '1',
		4297 => '0',
		4298 => '0',
		4299 => '1',
		4300 => '1',
		4301 => '1',
		4302 => '0',
		4303 => '0',
		4304 => '1',
		4305 => '1',
		4306 => '1',
		4307 => '0',
		4308 => '0',
		4309 => '0',
		4310 => '0',
		4311 => '0',
		4312 => '1',
		4313 => '1',
		4314 => '1',
		4315 => '1',
		4316 => '1',
		4317 => '0',
		4318 => '0',
		4319 => '1',
		4320 => '1',
		4321 => '1',
		4322 => '0',
		4323 => '0',
		4324 => '0',
		4325 => '0',
		4326 => '0',
		4327 => '0',
		4328 => '0',
		4329 => '1',
		4330 => '1',
		4331 => '1',
		4332 => '0',
		4333 => '0',
		4334 => '1',
		4335 => '1',
		4336 => '1',
		4337 => '0',
		4338 => '0',
		4339 => '1',
		4340 => '1',
		4341 => '1',
		4342 => '0',
		4343 => '0',
		4352 => '1',
		4353 => '1',
		4354 => '1',
		4355 => '0',
		4356 => '0',
		4357 => '1',
		4358 => '1',
		4359 => '1',
		4360 => '0',
		4361 => '0',
		4362 => '1',
		4363 => '1',
		4364 => '1',
		4365 => '0',
		4366 => '0',
		4367 => '1',
		4368 => '1',
		4369 => '1',
		4370 => '0',
		4371 => '0',
		4372 => '1',
		4373 => '1',
		4374 => '1',
		4375 => '0',
		4376 => '0',
		4377 => '1',
		4378 => '1',
		4379 => '1',
		4380 => '0',
		4381 => '0',
		4382 => '1',
		4383 => '1',
		4384 => '1',
		4385 => '1',
		4386 => '1',
		4387 => '1',
		4388 => '1',
		4389 => '1',
		4390 => '0',
		4391 => '0',
		4392 => '0',
		4393 => '0',
		4394 => '0',
		4395 => '1',
		4396 => '1',
		4397 => '1',
		4398 => '0',
		4399 => '1',
		4400 => '1',
		4401 => '1',
		4402 => '0',
		4403 => '0',
		4404 => '0',
		4405 => '0',
		4406 => '0',
		4407 => '1',
		4408 => '1',
		4409 => '1',
		4410 => '0',
		4411 => '0',
		4412 => '1',
		4413 => '1',
		4414 => '1',
		4415 => '0',
		4416 => '0',
		4417 => '1',
		4418 => '1',
		4419 => '1',
		4420 => '0',
		4421 => '0',
		4422 => '1',
		4423 => '1',
		4424 => '1',
		4425 => '0',
		4426 => '0',
		4427 => '1',
		4428 => '1',
		4429 => '1',
		4430 => '0',
		4431 => '0',
		4432 => '1',
		4433 => '1',
		4434 => '1',
		4435 => '0',
		4436 => '0',
		4437 => '1',
		4438 => '1',
		4439 => '1',
		4440 => '1',
		4441 => '1',
		4442 => '1',
		4443 => '1',
		4444 => '1',
		4445 => '0',
		4446 => '0',
		4447 => '1',
		4448 => '1',
		4449 => '1',
		4450 => '0',
		4451 => '0',
		4452 => '1',
		4453 => '1',
		4454 => '1',
		4455 => '1',
		4456 => '1',
		4457 => '1',
		4458 => '1',
		4459 => '1',
		4460 => '0',
		4461 => '0',
		4462 => '1',
		4463 => '1',
		4464 => '1',
		4465 => '1',
		4466 => '1',
		4467 => '1',
		4468 => '1',
		4469 => '1',
		4470 => '0',
		4471 => '0',
		4480 => '1',
		4481 => '1',
		4482 => '1',
		4483 => '0',
		4484 => '0',
		4485 => '1',
		4486 => '1',
		4487 => '1',
		4488 => '0',
		4489 => '0',
		4490 => '1',
		4491 => '1',
		4492 => '1',
		4493 => '0',
		4494 => '0',
		4495 => '1',
		4496 => '1',
		4497 => '1',
		4498 => '0',
		4499 => '0',
		4500 => '1',
		4501 => '1',
		4502 => '1',
		4503 => '0',
		4504 => '0',
		4505 => '1',
		4506 => '1',
		4507 => '1',
		4508 => '0',
		4509 => '0',
		4510 => '1',
		4511 => '1',
		4512 => '1',
		4513 => '0',
		4514 => '0',
		4515 => '1',
		4516 => '1',
		4517 => '1',
		4518 => '0',
		4519 => '0',
		4520 => '0',
		4521 => '0',
		4522 => '0',
		4523 => '1',
		4524 => '1',
		4525 => '1',
		4526 => '0',
		4527 => '1',
		4528 => '1',
		4529 => '1',
		4530 => '0',
		4531 => '0',
		4532 => '0',
		4533 => '0',
		4534 => '0',
		4535 => '1',
		4536 => '1',
		4537 => '1',
		4538 => '0',
		4539 => '0',
		4540 => '1',
		4541 => '1',
		4542 => '1',
		4543 => '0',
		4544 => '0',
		4545 => '1',
		4546 => '1',
		4547 => '1',
		4548 => '0',
		4549 => '0',
		4550 => '1',
		4551 => '1',
		4552 => '1',
		4553 => '0',
		4554 => '0',
		4555 => '1',
		4556 => '1',
		4557 => '1',
		4558 => '0',
		4559 => '0',
		4560 => '1',
		4561 => '1',
		4562 => '1',
		4563 => '0',
		4564 => '0',
		4565 => '1',
		4566 => '1',
		4567 => '1',
		4568 => '0',
		4569 => '0',
		4570 => '1',
		4571 => '1',
		4572 => '1',
		4573 => '0',
		4574 => '0',
		4575 => '1',
		4576 => '1',
		4577 => '1',
		4578 => '0',
		4579 => '0',
		4580 => '1',
		4581 => '1',
		4582 => '1',
		4583 => '1',
		4584 => '1',
		4585 => '1',
		4586 => '1',
		4587 => '1',
		4588 => '0',
		4589 => '0',
		4590 => '1',
		4591 => '1',
		4592 => '1',
		4593 => '1',
		4594 => '1',
		4595 => '1',
		4596 => '1',
		4597 => '1',
		4598 => '0',
		4599 => '0',
		4608 => '1',
		4609 => '1',
		4610 => '1',
		4611 => '0',
		4612 => '0',
		4613 => '1',
		4614 => '1',
		4615 => '1',
		4616 => '0',
		4617 => '0',
		4618 => '1',
		4619 => '1',
		4620 => '1',
		4621 => '0',
		4622 => '0',
		4623 => '1',
		4624 => '1',
		4625 => '1',
		4626 => '0',
		4627 => '0',
		4628 => '1',
		4629 => '1',
		4630 => '1',
		4631 => '0',
		4632 => '0',
		4633 => '1',
		4634 => '1',
		4635 => '1',
		4636 => '0',
		4637 => '0',
		4638 => '1',
		4639 => '1',
		4640 => '1',
		4641 => '0',
		4642 => '0',
		4643 => '1',
		4644 => '1',
		4645 => '1',
		4646 => '0',
		4647 => '0',
		4648 => '0',
		4649 => '0',
		4650 => '0',
		4651 => '1',
		4652 => '1',
		4653 => '1',
		4654 => '0',
		4655 => '1',
		4656 => '1',
		4657 => '1',
		4658 => '0',
		4659 => '0',
		4660 => '0',
		4661 => '0',
		4662 => '0',
		4663 => '1',
		4664 => '1',
		4665 => '1',
		4666 => '0',
		4667 => '0',
		4668 => '1',
		4669 => '1',
		4670 => '1',
		4671 => '0',
		4672 => '0',
		4673 => '1',
		4674 => '1',
		4675 => '1',
		4676 => '0',
		4677 => '0',
		4678 => '1',
		4679 => '1',
		4680 => '1',
		4681 => '0',
		4682 => '0',
		4683 => '1',
		4684 => '1',
		4685 => '1',
		4686 => '0',
		4687 => '0',
		4688 => '1',
		4689 => '1',
		4690 => '1',
		4691 => '0',
		4692 => '0',
		4693 => '1',
		4694 => '1',
		4695 => '1',
		4696 => '0',
		4697 => '0',
		4698 => '1',
		4699 => '1',
		4700 => '1',
		4701 => '0',
		4702 => '0',
		4703 => '1',
		4704 => '1',
		4705 => '1',
		4706 => '0',
		4707 => '0',
		4708 => '1',
		4709 => '1',
		4710 => '1',
		4711 => '1',
		4712 => '1',
		4713 => '1',
		4714 => '1',
		4715 => '1',
		4716 => '0',
		4717 => '0',
		4718 => '1',
		4719 => '1',
		4720 => '1',
		4721 => '1',
		4722 => '1',
		4723 => '1',
		4724 => '1',
		4725 => '1',
		4726 => '0',
		4727 => '0',
		4736 => '1',
		4737 => '1',
		4738 => '1',
		4739 => '1',
		4740 => '1',
		4741 => '0',
		4742 => '0',
		4743 => '0',
		4744 => '1',
		4745 => '1',
		4746 => '1',
		4747 => '1',
		4748 => '1',
		4749 => '0',
		4750 => '0',
		4751 => '1',
		4752 => '1',
		4753 => '1',
		4754 => '0',
		4755 => '0',
		4756 => '1',
		4757 => '1',
		4758 => '1',
		4759 => '0',
		4760 => '0',
		4761 => '1',
		4762 => '1',
		4763 => '1',
		4764 => '0',
		4765 => '0',
		4766 => '0',
		4767 => '0',
		4768 => '0',
		4769 => '0',
		4770 => '0',
		4771 => '1',
		4772 => '1',
		4773 => '1',
		4774 => '0',
		4775 => '0',
		4776 => '0',
		4777 => '0',
		4778 => '0',
		4779 => '1',
		4780 => '1',
		4781 => '1',
		4782 => '0',
		4783 => '1',
		4784 => '1',
		4785 => '1',
		4786 => '0',
		4787 => '0',
		4788 => '0',
		4789 => '0',
		4790 => '0',
		4791 => '1',
		4792 => '1',
		4793 => '1',
		4794 => '0',
		4795 => '0',
		4796 => '0',
		4797 => '0',
		4798 => '0',
		4799 => '0',
		4800 => '0',
		4801 => '1',
		4802 => '1',
		4803 => '1',
		4804 => '0',
		4805 => '0',
		4806 => '1',
		4807 => '1',
		4808 => '1',
		4809 => '0',
		4810 => '0',
		4811 => '1',
		4812 => '1',
		4813 => '1',
		4814 => '0',
		4815 => '0',
		4816 => '1',
		4817 => '1',
		4818 => '1',
		4819 => '0',
		4820 => '0',
		4821 => '1',
		4822 => '1',
		4823 => '1',
		4824 => '0',
		4825 => '0',
		4826 => '1',
		4827 => '1',
		4828 => '1',
		4829 => '0',
		4830 => '0',
		4831 => '1',
		4832 => '1',
		4833 => '1',
		4834 => '0',
		4835 => '0',
		4836 => '0',
		4837 => '0',
		4838 => '0',
		4839 => '0',
		4840 => '0',
		4841 => '1',
		4842 => '1',
		4843 => '1',
		4844 => '0',
		4845 => '0',
		4846 => '1',
		4847 => '1',
		4848 => '1',
		4849 => '0',
		4850 => '0',
		4851 => '1',
		4852 => '1',
		4853 => '1',
		4854 => '0',
		4855 => '0',
		4864 => '1',
		4865 => '1',
		4866 => '1',
		4867 => '1',
		4868 => '1',
		4869 => '0',
		4870 => '0',
		4871 => '0',
		4872 => '1',
		4873 => '1',
		4874 => '1',
		4875 => '1',
		4876 => '1',
		4877 => '0',
		4878 => '0',
		4879 => '1',
		4880 => '1',
		4881 => '1',
		4882 => '0',
		4883 => '0',
		4884 => '1',
		4885 => '1',
		4886 => '1',
		4887 => '0',
		4888 => '0',
		4889 => '1',
		4890 => '1',
		4891 => '1',
		4892 => '0',
		4893 => '0',
		4894 => '0',
		4895 => '0',
		4896 => '0',
		4897 => '0',
		4898 => '0',
		4899 => '1',
		4900 => '1',
		4901 => '1',
		4902 => '0',
		4903 => '0',
		4904 => '0',
		4905 => '0',
		4906 => '0',
		4907 => '1',
		4908 => '1',
		4909 => '1',
		4910 => '0',
		4911 => '1',
		4912 => '1',
		4913 => '1',
		4914 => '0',
		4915 => '0',
		4916 => '0',
		4917 => '0',
		4918 => '0',
		4919 => '1',
		4920 => '1',
		4921 => '1',
		4922 => '0',
		4923 => '0',
		4924 => '0',
		4925 => '0',
		4926 => '0',
		4927 => '0',
		4928 => '0',
		4929 => '1',
		4930 => '1',
		4931 => '1',
		4932 => '0',
		4933 => '0',
		4934 => '1',
		4935 => '1',
		4936 => '1',
		4937 => '0',
		4938 => '0',
		4939 => '1',
		4940 => '1',
		4941 => '1',
		4942 => '0',
		4943 => '0',
		4944 => '1',
		4945 => '1',
		4946 => '1',
		4947 => '0',
		4948 => '0',
		4949 => '1',
		4950 => '1',
		4951 => '1',
		4952 => '0',
		4953 => '0',
		4954 => '1',
		4955 => '1',
		4956 => '1',
		4957 => '0',
		4958 => '0',
		4959 => '1',
		4960 => '1',
		4961 => '1',
		4962 => '0',
		4963 => '0',
		4964 => '0',
		4965 => '0',
		4966 => '0',
		4967 => '0',
		4968 => '0',
		4969 => '1',
		4970 => '1',
		4971 => '1',
		4972 => '0',
		4973 => '0',
		4974 => '1',
		4975 => '1',
		4976 => '1',
		4977 => '0',
		4978 => '0',
		4979 => '1',
		4980 => '1',
		4981 => '1',
		4982 => '0',
		4983 => '0',
		4992 => '0',
		4993 => '0',
		4994 => '0',
		4995 => '1',
		4996 => '1',
		4997 => '1',
		4998 => '1',
		4999 => '1',
		5000 => '1',
		5001 => '1',
		5002 => '0',
		5003 => '0',
		5004 => '0',
		5005 => '0',
		5006 => '0',
		5007 => '1',
		5008 => '1',
		5009 => '1',
		5010 => '1',
		5011 => '1',
		5012 => '1',
		5013 => '1',
		5014 => '1',
		5015 => '0',
		5016 => '0',
		5017 => '1',
		5018 => '1',
		5019 => '1',
		5020 => '1',
		5021 => '1',
		5022 => '1',
		5023 => '1',
		5024 => '1',
		5025 => '1',
		5026 => '1',
		5027 => '1',
		5028 => '1',
		5029 => '1',
		5030 => '0',
		5031 => '0',
		5032 => '0',
		5033 => '0',
		5034 => '0',
		5035 => '1',
		5036 => '1',
		5037 => '1',
		5038 => '1',
		5039 => '1',
		5040 => '1',
		5041 => '1',
		5042 => '0',
		5043 => '0',
		5044 => '0',
		5045 => '0',
		5046 => '0',
		5047 => '1',
		5048 => '1',
		5049 => '1',
		5050 => '1',
		5051 => '1',
		5052 => '1',
		5053 => '1',
		5054 => '1',
		5055 => '1',
		5056 => '1',
		5057 => '1',
		5058 => '1',
		5059 => '1',
		5060 => '0',
		5061 => '0',
		5062 => '1',
		5063 => '1',
		5064 => '1',
		5065 => '1',
		5066 => '1',
		5067 => '1',
		5068 => '1',
		5069 => '1',
		5070 => '0',
		5071 => '0',
		5072 => '1',
		5073 => '1',
		5074 => '1',
		5075 => '1',
		5076 => '1',
		5077 => '1',
		5078 => '1',
		5079 => '1',
		5080 => '1',
		5081 => '1',
		5082 => '1',
		5083 => '1',
		5084 => '1',
		5085 => '0',
		5086 => '0',
		5087 => '1',
		5088 => '1',
		5089 => '1',
		5090 => '1',
		5091 => '1',
		5092 => '1',
		5093 => '1',
		5094 => '1',
		5095 => '1',
		5096 => '1',
		5097 => '1',
		5098 => '1',
		5099 => '1',
		5100 => '0',
		5101 => '0',
		5102 => '1',
		5103 => '1',
		5104 => '1',
		5105 => '1',
		5106 => '1',
		5107 => '1',
		5108 => '1',
		5109 => '1',
		5110 => '0',
		5111 => '0',
		5120 => '0',
		5121 => '0',
		5122 => '0',
		5123 => '1',
		5124 => '1',
		5125 => '1',
		5126 => '1',
		5127 => '1',
		5128 => '1',
		5129 => '1',
		5130 => '0',
		5131 => '0',
		5132 => '0',
		5133 => '0',
		5134 => '0',
		5135 => '1',
		5136 => '1',
		5137 => '1',
		5138 => '1',
		5139 => '1',
		5140 => '1',
		5141 => '1',
		5142 => '1',
		5143 => '0',
		5144 => '0',
		5145 => '1',
		5146 => '1',
		5147 => '1',
		5148 => '1',
		5149 => '1',
		5150 => '1',
		5151 => '1',
		5152 => '1',
		5153 => '1',
		5154 => '1',
		5155 => '1',
		5156 => '1',
		5157 => '1',
		5158 => '0',
		5159 => '0',
		5160 => '0',
		5161 => '0',
		5162 => '0',
		5163 => '1',
		5164 => '1',
		5165 => '1',
		5166 => '1',
		5167 => '1',
		5168 => '1',
		5169 => '1',
		5170 => '0',
		5171 => '0',
		5172 => '0',
		5173 => '0',
		5174 => '0',
		5175 => '1',
		5176 => '1',
		5177 => '1',
		5178 => '1',
		5179 => '1',
		5180 => '1',
		5181 => '1',
		5182 => '1',
		5183 => '1',
		5184 => '1',
		5185 => '1',
		5186 => '1',
		5187 => '1',
		5188 => '0',
		5189 => '0',
		5190 => '1',
		5191 => '1',
		5192 => '1',
		5193 => '1',
		5194 => '1',
		5195 => '1',
		5196 => '1',
		5197 => '1',
		5198 => '0',
		5199 => '0',
		5200 => '1',
		5201 => '1',
		5202 => '1',
		5203 => '1',
		5204 => '1',
		5205 => '1',
		5206 => '1',
		5207 => '1',
		5208 => '1',
		5209 => '1',
		5210 => '1',
		5211 => '1',
		5212 => '1',
		5213 => '0',
		5214 => '0',
		5215 => '1',
		5216 => '1',
		5217 => '1',
		5218 => '1',
		5219 => '1',
		5220 => '1',
		5221 => '1',
		5222 => '1',
		5223 => '1',
		5224 => '1',
		5225 => '1',
		5226 => '1',
		5227 => '1',
		5228 => '0',
		5229 => '0',
		5230 => '1',
		5231 => '1',
		5232 => '1',
		5233 => '1',
		5234 => '1',
		5235 => '1',
		5236 => '1',
		5237 => '1',
		5238 => '0',
		5239 => '0',
		5248 => '0',
		5249 => '0',
		5250 => '0',
		5251 => '1',
		5252 => '1',
		5253 => '1',
		5254 => '1',
		5255 => '1',
		5256 => '1',
		5257 => '1',
		5258 => '0',
		5259 => '0',
		5260 => '0',
		5261 => '0',
		5262 => '0',
		5263 => '1',
		5264 => '1',
		5265 => '1',
		5266 => '1',
		5267 => '1',
		5268 => '1',
		5269 => '1',
		5270 => '1',
		5271 => '0',
		5272 => '0',
		5273 => '1',
		5274 => '1',
		5275 => '1',
		5276 => '1',
		5277 => '1',
		5278 => '1',
		5279 => '1',
		5280 => '1',
		5281 => '1',
		5282 => '1',
		5283 => '1',
		5284 => '1',
		5285 => '1',
		5286 => '0',
		5287 => '0',
		5288 => '0',
		5289 => '0',
		5290 => '0',
		5291 => '1',
		5292 => '1',
		5293 => '1',
		5294 => '1',
		5295 => '1',
		5296 => '1',
		5297 => '1',
		5298 => '0',
		5299 => '0',
		5300 => '0',
		5301 => '0',
		5302 => '0',
		5303 => '1',
		5304 => '1',
		5305 => '1',
		5306 => '1',
		5307 => '1',
		5308 => '1',
		5309 => '1',
		5310 => '1',
		5311 => '1',
		5312 => '1',
		5313 => '1',
		5314 => '1',
		5315 => '1',
		5316 => '0',
		5317 => '0',
		5318 => '1',
		5319 => '1',
		5320 => '1',
		5321 => '1',
		5322 => '1',
		5323 => '1',
		5324 => '1',
		5325 => '1',
		5326 => '0',
		5327 => '0',
		5328 => '1',
		5329 => '1',
		5330 => '1',
		5331 => '1',
		5332 => '1',
		5333 => '1',
		5334 => '1',
		5335 => '1',
		5336 => '1',
		5337 => '1',
		5338 => '1',
		5339 => '1',
		5340 => '1',
		5341 => '0',
		5342 => '0',
		5343 => '1',
		5344 => '1',
		5345 => '1',
		5346 => '1',
		5347 => '1',
		5348 => '1',
		5349 => '1',
		5350 => '1',
		5351 => '1',
		5352 => '1',
		5353 => '1',
		5354 => '1',
		5355 => '1',
		5356 => '0',
		5357 => '0',
		5358 => '1',
		5359 => '1',
		5360 => '1',
		5361 => '1',
		5362 => '1',
		5363 => '1',
		5364 => '1',
		5365 => '1',
		5366 => '0',
		5367 => '0',
		5376 => '0',
		5377 => '0',
		5378 => '0',
		5379 => '0',
		5380 => '0',
		5381 => '0',
		5382 => '0',
		5383 => '0',
		5384 => '0',
		5385 => '0',
		5386 => '0',
		5387 => '0',
		5388 => '0',
		5389 => '0',
		5390 => '0',
		5391 => '0',
		5392 => '0',
		5393 => '0',
		5394 => '0',
		5395 => '0',
		5396 => '0',
		5397 => '0',
		5398 => '0',
		5399 => '0',
		5400 => '0',
		5401 => '0',
		5402 => '0',
		5403 => '0',
		5404 => '0',
		5405 => '0',
		5406 => '0',
		5407 => '0',
		5408 => '0',
		5409 => '0',
		5410 => '0',
		5411 => '0',
		5412 => '0',
		5413 => '0',
		5414 => '0',
		5415 => '0',
		5416 => '0',
		5417 => '0',
		5418 => '0',
		5419 => '0',
		5420 => '0',
		5421 => '0',
		5422 => '0',
		5423 => '0',
		5424 => '0',
		5425 => '0',
		5426 => '0',
		5427 => '0',
		5428 => '0',
		5429 => '0',
		5430 => '0',
		5431 => '0',
		5432 => '0',
		5433 => '0',
		5434 => '0',
		5435 => '0',
		5436 => '0',
		5437 => '0',
		5438 => '0',
		5439 => '0',
		5440 => '0',
		5441 => '0',
		5442 => '0',
		5443 => '0',
		5444 => '0',
		5445 => '0',
		5446 => '0',
		5447 => '0',
		5448 => '0',
		5449 => '0',
		5450 => '0',
		5451 => '0',
		5452 => '0',
		5453 => '0',
		5454 => '0',
		5455 => '0',
		5456 => '0',
		5457 => '0',
		5458 => '0',
		5459 => '0',
		5460 => '0',
		5461 => '0',
		5462 => '0',
		5463 => '0',
		5464 => '0',
		5465 => '0',
		5466 => '0',
		5467 => '0',
		5468 => '0',
		5469 => '0',
		5470 => '0',
		5471 => '0',
		5472 => '0',
		5473 => '0',
		5474 => '0',
		5475 => '0',
		5476 => '0',
		5477 => '0',
		5478 => '0',
		5479 => '0',
		5480 => '0',
		5481 => '0',
		5482 => '0',
		5483 => '0',
		5484 => '0',
		5485 => '0',
		5486 => '0',
		5487 => '0',
		5488 => '0',
		5489 => '0',
		5490 => '0',
		5491 => '0',
		5492 => '0',
		5493 => '0',
		5494 => '0',
		5495 => '0',
		5504 => '0',
		5505 => '0',
		5506 => '0',
		5507 => '0',
		5508 => '0',
		5509 => '0',
		5510 => '0',
		5511 => '0',
		5512 => '0',
		5513 => '0',
		5514 => '0',
		5515 => '0',
		5516 => '0',
		5517 => '0',
		5518 => '0',
		5519 => '0',
		5520 => '0',
		5521 => '0',
		5522 => '0',
		5523 => '0',
		5524 => '0',
		5525 => '0',
		5526 => '0',
		5527 => '0',
		5528 => '0',
		5529 => '0',
		5530 => '0',
		5531 => '0',
		5532 => '0',
		5533 => '0',
		5534 => '0',
		5535 => '0',
		5536 => '0',
		5537 => '0',
		5538 => '0',
		5539 => '0',
		5540 => '0',
		5541 => '0',
		5542 => '0',
		5543 => '0',
		5544 => '0',
		5545 => '0',
		5546 => '0',
		5547 => '0',
		5548 => '0',
		5549 => '0',
		5550 => '0',
		5551 => '0',
		5552 => '0',
		5553 => '0',
		5554 => '0',
		5555 => '0',
		5556 => '0',
		5557 => '0',
		5558 => '0',
		5559 => '0',
		5560 => '0',
		5561 => '0',
		5562 => '0',
		5563 => '0',
		5564 => '0',
		5565 => '0',
		5566 => '0',
		5567 => '0',
		5568 => '0',
		5569 => '0',
		5570 => '0',
		5571 => '0',
		5572 => '0',
		5573 => '0',
		5574 => '0',
		5575 => '0',
		5576 => '0',
		5577 => '0',
		5578 => '0',
		5579 => '0',
		5580 => '0',
		5581 => '0',
		5582 => '0',
		5583 => '0',
		5584 => '0',
		5585 => '0',
		5586 => '0',
		5587 => '0',
		5588 => '0',
		5589 => '0',
		5590 => '0',
		5591 => '0',
		5592 => '0',
		5593 => '0',
		5594 => '0',
		5595 => '0',
		5596 => '0',
		5597 => '0',
		5598 => '0',
		5599 => '0',
		5600 => '0',
		5601 => '0',
		5602 => '0',
		5603 => '0',
		5604 => '0',
		5605 => '0',
		5606 => '0',
		5607 => '0',
		5608 => '0',
		5609 => '0',
		5610 => '0',
		5611 => '0',
		5612 => '0',
		5613 => '0',
		5614 => '0',
		5615 => '0',
		5616 => '0',
		5617 => '0',
		5618 => '0',
		5619 => '0',
		5620 => '0',
		5621 => '0',
		5622 => '0',
		5623 => '0',
		5632 => '0',
		5633 => '0',
		5634 => '0',
		5635 => '0',
		5636 => '0',
		5637 => '0',
		5638 => '0',
		5639 => '0',
		5640 => '0',
		5641 => '0',
		5642 => '0',
		5643 => '0',
		5644 => '0',
		5645 => '0',
		5646 => '0',
		5647 => '0',
		5648 => '0',
		5649 => '0',
		5650 => '0',
		5651 => '0',
		5652 => '0',
		5653 => '0',
		5654 => '0',
		5655 => '0',
		5656 => '0',
		5657 => '0',
		5658 => '0',
		5659 => '0',
		5660 => '0',
		5661 => '0',
		5662 => '0',
		5663 => '0',
		5664 => '0',
		5665 => '0',
		5666 => '0',
		5667 => '0',
		5668 => '0',
		5669 => '0',
		5670 => '0',
		5671 => '0',
		5672 => '0',
		5673 => '0',
		5674 => '0',
		5675 => '0',
		5676 => '0',
		5677 => '0',
		5678 => '0',
		5679 => '0',
		5680 => '0',
		5681 => '0',
		5682 => '0',
		5683 => '0',
		5684 => '0',
		5685 => '0',
		5686 => '0',
		5687 => '0',
		5688 => '0',
		5689 => '0',
		5690 => '0',
		5691 => '0',
		5692 => '0',
		5693 => '0',
		5694 => '0',
		5695 => '0',
		5696 => '0',
		5697 => '0',
		5698 => '0',
		5699 => '0',
		5700 => '0',
		5701 => '0',
		5702 => '0',
		5703 => '0',
		5704 => '0',
		5705 => '0',
		5706 => '0',
		5707 => '0',
		5708 => '0',
		5709 => '0',
		5710 => '0',
		5711 => '0',
		5712 => '0',
		5713 => '0',
		5714 => '0',
		5715 => '0',
		5716 => '0',
		5717 => '0',
		5718 => '0',
		5719 => '0',
		5720 => '0',
		5721 => '0',
		5722 => '0',
		5723 => '0',
		5724 => '0',
		5725 => '0',
		5726 => '0',
		5727 => '0',
		5728 => '0',
		5729 => '0',
		5730 => '0',
		5731 => '0',
		5732 => '0',
		5733 => '0',
		5734 => '0',
		5735 => '0',
		5736 => '0',
		5737 => '0',
		5738 => '0',
		5739 => '0',
		5740 => '0',
		5741 => '0',
		5742 => '0',
		5743 => '0',
		5744 => '0',
		5745 => '0',
		5746 => '0',
		5747 => '0',
		5748 => '0',
		5749 => '0',
		5750 => '0',
		5751 => '0',
		5760 => '0',
		5761 => '0',
		5762 => '0',
		5763 => '0',
		5764 => '0',
		5765 => '0',
		5766 => '0',
		5767 => '0',
		5768 => '0',
		5769 => '0',
		5770 => '0',
		5771 => '0',
		5772 => '0',
		5773 => '0',
		5774 => '0',
		5775 => '0',
		5776 => '0',
		5777 => '0',
		5778 => '0',
		5779 => '0',
		5780 => '0',
		5781 => '0',
		5782 => '0',
		5783 => '0',
		5784 => '0',
		5785 => '0',
		5786 => '0',
		5787 => '0',
		5788 => '0',
		5789 => '0',
		5790 => '0',
		5791 => '0',
		5792 => '0',
		5793 => '0',
		5794 => '0',
		5795 => '0',
		5796 => '0',
		5797 => '0',
		5798 => '0',
		5799 => '0',
		5800 => '0',
		5801 => '0',
		5802 => '0',
		5803 => '0',
		5804 => '0',
		5805 => '0',
		5806 => '0',
		5807 => '0',
		5808 => '0',
		5809 => '0',
		5810 => '0',
		5811 => '0',
		5812 => '0',
		5813 => '0',
		5814 => '0',
		5815 => '0',
		5816 => '0',
		5817 => '0',
		5818 => '0',
		5819 => '0',
		5820 => '0',
		5821 => '0',
		5822 => '0',
		5823 => '0',
		5824 => '0',
		5825 => '0',
		5826 => '0',
		5827 => '0',
		5828 => '0',
		5829 => '0',
		5830 => '0',
		5831 => '0',
		5832 => '0',
		5833 => '0',
		5834 => '0',
		5835 => '0',
		5836 => '0',
		5837 => '0',
		5838 => '0',
		5839 => '0',
		5840 => '0',
		5841 => '0',
		5842 => '0',
		5843 => '0',
		5844 => '0',
		5845 => '0',
		5846 => '0',
		5847 => '0',
		5848 => '0',
		5849 => '0',
		5850 => '0',
		5851 => '0',
		5852 => '0',
		5853 => '0',
		5854 => '0',
		5855 => '0',
		5856 => '0',
		5857 => '0',
		5858 => '0',
		5859 => '0',
		5860 => '0',
		5861 => '0',
		5862 => '0',
		5863 => '0',
		5864 => '0',
		5865 => '0',
		5866 => '0',
		5867 => '0',
		5868 => '0',
		5869 => '0',
		5870 => '0',
		5871 => '0',
		5872 => '0',
		5873 => '0',
		5874 => '0',
		5875 => '0',
		5876 => '0',
		5877 => '0',
		5878 => '0',
		5879 => '0',
		5888 => '0',
		5889 => '0',
		5890 => '0',
		5891 => '0',
		5892 => '0',
		5893 => '0',
		5894 => '0',
		5895 => '0',
		5896 => '0',
		5897 => '0',
		5898 => '0',
		5899 => '0',
		5900 => '0',
		5901 => '0',
		5902 => '0',
		5903 => '0',
		5904 => '0',
		5905 => '0',
		5906 => '0',
		5907 => '0',
		5908 => '0',
		5909 => '0',
		5910 => '0',
		5911 => '0',
		5912 => '0',
		5913 => '0',
		5914 => '0',
		5915 => '0',
		5916 => '0',
		5917 => '0',
		5918 => '0',
		5919 => '0',
		5920 => '0',
		5921 => '0',
		5922 => '0',
		5923 => '0',
		5924 => '0',
		5925 => '0',
		5926 => '0',
		5927 => '0',
		5928 => '0',
		5929 => '0',
		5930 => '0',
		5931 => '0',
		5932 => '0',
		5933 => '0',
		5934 => '0',
		5935 => '0',
		5936 => '0',
		5937 => '0',
		5938 => '0',
		5939 => '0',
		5940 => '0',
		5941 => '0',
		5942 => '0',
		5943 => '0',
		5944 => '0',
		5945 => '0',
		5946 => '0',
		5947 => '0',
		5948 => '0',
		5949 => '0',
		5950 => '0',
		5951 => '0',
		5952 => '0',
		5953 => '0',
		5954 => '0',
		5955 => '0',
		5956 => '0',
		5957 => '0',
		5958 => '0',
		5959 => '0',
		5960 => '0',
		5961 => '0',
		5962 => '0',
		5963 => '0',
		5964 => '0',
		5965 => '0',
		5966 => '0',
		5967 => '0',
		5968 => '0',
		5969 => '0',
		5970 => '0',
		5971 => '0',
		5972 => '0',
		5973 => '0',
		5974 => '0',
		5975 => '0',
		5976 => '0',
		5977 => '0',
		5978 => '0',
		5979 => '0',
		5980 => '0',
		5981 => '0',
		5982 => '0',
		5983 => '0',
		5984 => '0',
		5985 => '0',
		5986 => '0',
		5987 => '0',
		5988 => '0',
		5989 => '0',
		5990 => '0',
		5991 => '0',
		5992 => '0',
		5993 => '0',
		5994 => '0',
		5995 => '0',
		5996 => '0',
		5997 => '0',
		5998 => '0',
		5999 => '0',
		6000 => '0',
		6001 => '0',
		6002 => '0',
		6003 => '0',
		6004 => '0',
		6005 => '0',
		6006 => '0',
		6007 => '0',
		6016 => '0',
		6017 => '0',
		6018 => '0',
		6019 => '0',
		6020 => '0',
		6021 => '0',
		6022 => '0',
		6023 => '0',
		6024 => '0',
		6025 => '0',
		6026 => '0',
		6027 => '0',
		6028 => '0',
		6029 => '0',
		6030 => '0',
		6031 => '0',
		6032 => '0',
		6033 => '0',
		6034 => '0',
		6035 => '0',
		6036 => '0',
		6037 => '0',
		6038 => '0',
		6039 => '0',
		6040 => '0',
		6041 => '0',
		6042 => '0',
		6043 => '0',
		6044 => '0',
		6045 => '0',
		6046 => '0',
		6047 => '0',
		6048 => '0',
		6049 => '0',
		6050 => '0',
		6051 => '0',
		6052 => '0',
		6053 => '0',
		6054 => '0',
		6055 => '0',
		6056 => '0',
		6057 => '0',
		6058 => '0',
		6059 => '0',
		6060 => '0',
		6061 => '0',
		6062 => '0',
		6063 => '0',
		6064 => '0',
		6065 => '0',
		6066 => '0',
		6067 => '0',
		6068 => '0',
		6069 => '0',
		6070 => '0',
		6071 => '0',
		6072 => '0',
		6073 => '0',
		6074 => '0',
		6075 => '0',
		6076 => '0',
		6077 => '0',
		6078 => '0',
		6079 => '0',
		6080 => '0',
		6081 => '0',
		6082 => '0',
		6083 => '0',
		6084 => '0',
		6085 => '0',
		6086 => '0',
		6087 => '0',
		6088 => '0',
		6089 => '0',
		6090 => '0',
		6091 => '0',
		6092 => '0',
		6093 => '0',
		6094 => '0',
		6095 => '0',
		6096 => '0',
		6097 => '0',
		6098 => '0',
		6099 => '0',
		6100 => '0',
		6101 => '0',
		6102 => '0',
		6103 => '0',
		6104 => '0',
		6105 => '0',
		6106 => '0',
		6107 => '0',
		6108 => '0',
		6109 => '0',
		6110 => '0',
		6111 => '0',
		6112 => '0',
		6113 => '0',
		6114 => '0',
		6115 => '0',
		6116 => '0',
		6117 => '0',
		6118 => '0',
		6119 => '0',
		6120 => '0',
		6121 => '0',
		6122 => '0',
		6123 => '0',
		6124 => '0',
		6125 => '0',
		6126 => '0',
		6127 => '0',
		6128 => '0',
		6129 => '0',
		6130 => '0',
		6131 => '0',
		6132 => '0',
		6133 => '0',
		6134 => '0',
		6135 => '0',
		6144 => '1',
		6145 => '1',
		6146 => '1',
		6147 => '1',
		6148 => '1',
		6149 => '1',
		6150 => '1',
		6151 => '1',
		6152 => '1',
		6153 => '1',
		6154 => '1',
		6155 => '1',
		6156 => '1',
		6157 => '0',
		6158 => '0',
		6159 => '1',
		6160 => '1',
		6161 => '1',
		6162 => '1',
		6163 => '1',
		6164 => '1',
		6165 => '1',
		6166 => '1',
		6167 => '0',
		6168 => '0',
		6169 => '1',
		6170 => '1',
		6171 => '1',
		6172 => '1',
		6173 => '1',
		6174 => '1',
		6175 => '1',
		6176 => '1',
		6177 => '1',
		6178 => '1',
		6179 => '1',
		6180 => '1',
		6181 => '1',
		6182 => '0',
		6183 => '0',
		6184 => '1',
		6185 => '1',
		6186 => '1',
		6187 => '1',
		6188 => '1',
		6189 => '1',
		6190 => '1',
		6191 => '1',
		6192 => '1',
		6193 => '1',
		6194 => '1',
		6195 => '1',
		6196 => '1',
		6197 => '0',
		6198 => '0',
		6199 => '1',
		6200 => '1',
		6201 => '1',
		6202 => '1',
		6203 => '1',
		6204 => '1',
		6205 => '1',
		6206 => '1',
		6207 => '1',
		6208 => '1',
		6209 => '1',
		6210 => '1',
		6211 => '1',
		6212 => '0',
		6213 => '0',
		6214 => '1',
		6215 => '1',
		6216 => '1',
		6217 => '1',
		6218 => '1',
		6219 => '1',
		6220 => '1',
		6221 => '1',
		6222 => '0',
		6223 => '0',
		6224 => '1',
		6225 => '1',
		6226 => '1',
		6227 => '1',
		6228 => '1',
		6229 => '1',
		6230 => '1',
		6231 => '1',
		6232 => '1',
		6233 => '1',
		6234 => '1',
		6235 => '1',
		6236 => '1',
		6237 => '0',
		6238 => '0',
		6239 => '1',
		6240 => '1',
		6241 => '1',
		6242 => '1',
		6243 => '1',
		6244 => '1',
		6245 => '1',
		6246 => '1',
		6247 => '1',
		6248 => '1',
		6249 => '1',
		6250 => '1',
		6251 => '1',
		6252 => '0',
		6253 => '0',
		6254 => '1',
		6255 => '1',
		6256 => '1',
		6257 => '1',
		6258 => '1',
		6259 => '1',
		6260 => '1',
		6261 => '1',
		6262 => '0',
		6263 => '0',
		6272 => '1',
		6273 => '1',
		6274 => '1',
		6275 => '1',
		6276 => '1',
		6277 => '1',
		6278 => '1',
		6279 => '1',
		6280 => '1',
		6281 => '1',
		6282 => '1',
		6283 => '1',
		6284 => '1',
		6285 => '0',
		6286 => '0',
		6287 => '1',
		6288 => '1',
		6289 => '1',
		6290 => '1',
		6291 => '1',
		6292 => '1',
		6293 => '1',
		6294 => '1',
		6295 => '0',
		6296 => '0',
		6297 => '1',
		6298 => '1',
		6299 => '1',
		6300 => '1',
		6301 => '1',
		6302 => '1',
		6303 => '1',
		6304 => '1',
		6305 => '1',
		6306 => '1',
		6307 => '1',
		6308 => '1',
		6309 => '1',
		6310 => '0',
		6311 => '0',
		6312 => '1',
		6313 => '1',
		6314 => '1',
		6315 => '1',
		6316 => '1',
		6317 => '1',
		6318 => '1',
		6319 => '1',
		6320 => '1',
		6321 => '1',
		6322 => '1',
		6323 => '1',
		6324 => '1',
		6325 => '0',
		6326 => '0',
		6327 => '1',
		6328 => '1',
		6329 => '1',
		6330 => '1',
		6331 => '1',
		6332 => '1',
		6333 => '1',
		6334 => '1',
		6335 => '1',
		6336 => '1',
		6337 => '1',
		6338 => '1',
		6339 => '1',
		6340 => '0',
		6341 => '0',
		6342 => '1',
		6343 => '1',
		6344 => '1',
		6345 => '1',
		6346 => '1',
		6347 => '1',
		6348 => '1',
		6349 => '1',
		6350 => '0',
		6351 => '0',
		6352 => '1',
		6353 => '1',
		6354 => '1',
		6355 => '1',
		6356 => '1',
		6357 => '1',
		6358 => '1',
		6359 => '1',
		6360 => '1',
		6361 => '1',
		6362 => '1',
		6363 => '1',
		6364 => '1',
		6365 => '0',
		6366 => '0',
		6367 => '1',
		6368 => '1',
		6369 => '1',
		6370 => '1',
		6371 => '1',
		6372 => '1',
		6373 => '1',
		6374 => '1',
		6375 => '1',
		6376 => '1',
		6377 => '1',
		6378 => '1',
		6379 => '1',
		6380 => '0',
		6381 => '0',
		6382 => '1',
		6383 => '1',
		6384 => '1',
		6385 => '1',
		6386 => '1',
		6387 => '1',
		6388 => '1',
		6389 => '1',
		6390 => '0',
		6391 => '0',
		6400 => '1',
		6401 => '1',
		6402 => '1',
		6403 => '1',
		6404 => '1',
		6405 => '1',
		6406 => '1',
		6407 => '1',
		6408 => '1',
		6409 => '1',
		6410 => '1',
		6411 => '1',
		6412 => '1',
		6413 => '0',
		6414 => '0',
		6415 => '1',
		6416 => '1',
		6417 => '1',
		6418 => '1',
		6419 => '1',
		6420 => '1',
		6421 => '1',
		6422 => '1',
		6423 => '0',
		6424 => '0',
		6425 => '1',
		6426 => '1',
		6427 => '1',
		6428 => '1',
		6429 => '1',
		6430 => '1',
		6431 => '1',
		6432 => '1',
		6433 => '1',
		6434 => '1',
		6435 => '1',
		6436 => '1',
		6437 => '1',
		6438 => '0',
		6439 => '0',
		6440 => '1',
		6441 => '1',
		6442 => '1',
		6443 => '1',
		6444 => '1',
		6445 => '1',
		6446 => '1',
		6447 => '1',
		6448 => '1',
		6449 => '1',
		6450 => '1',
		6451 => '1',
		6452 => '1',
		6453 => '0',
		6454 => '0',
		6455 => '1',
		6456 => '1',
		6457 => '1',
		6458 => '1',
		6459 => '1',
		6460 => '1',
		6461 => '1',
		6462 => '1',
		6463 => '1',
		6464 => '1',
		6465 => '1',
		6466 => '1',
		6467 => '1',
		6468 => '0',
		6469 => '0',
		6470 => '1',
		6471 => '1',
		6472 => '1',
		6473 => '1',
		6474 => '1',
		6475 => '1',
		6476 => '1',
		6477 => '1',
		6478 => '0',
		6479 => '0',
		6480 => '1',
		6481 => '1',
		6482 => '1',
		6483 => '1',
		6484 => '1',
		6485 => '1',
		6486 => '1',
		6487 => '1',
		6488 => '1',
		6489 => '1',
		6490 => '1',
		6491 => '1',
		6492 => '1',
		6493 => '0',
		6494 => '0',
		6495 => '1',
		6496 => '1',
		6497 => '1',
		6498 => '1',
		6499 => '1',
		6500 => '1',
		6501 => '1',
		6502 => '1',
		6503 => '1',
		6504 => '1',
		6505 => '1',
		6506 => '1',
		6507 => '1',
		6508 => '0',
		6509 => '0',
		6510 => '1',
		6511 => '1',
		6512 => '1',
		6513 => '1',
		6514 => '1',
		6515 => '1',
		6516 => '1',
		6517 => '1',
		6518 => '0',
		6519 => '0',
		6528 => '1',
		6529 => '1',
		6530 => '1',
		6531 => '0',
		6532 => '0',
		6533 => '1',
		6534 => '1',
		6535 => '1',
		6536 => '0',
		6537 => '0',
		6538 => '1',
		6539 => '1',
		6540 => '1',
		6541 => '0',
		6542 => '0',
		6543 => '1',
		6544 => '1',
		6545 => '1',
		6546 => '0',
		6547 => '0',
		6548 => '1',
		6549 => '1',
		6550 => '1',
		6551 => '0',
		6552 => '0',
		6553 => '1',
		6554 => '1',
		6555 => '1',
		6556 => '0',
		6557 => '0',
		6558 => '0',
		6559 => '0',
		6560 => '0',
		6561 => '0',
		6562 => '0',
		6563 => '1',
		6564 => '1',
		6565 => '1',
		6566 => '0',
		6567 => '0',
		6568 => '1',
		6569 => '1',
		6570 => '1',
		6571 => '0',
		6572 => '0',
		6573 => '0',
		6574 => '0',
		6575 => '0',
		6576 => '0',
		6577 => '0',
		6578 => '1',
		6579 => '1',
		6580 => '1',
		6581 => '0',
		6582 => '0',
		6583 => '1',
		6584 => '1',
		6585 => '1',
		6586 => '0',
		6587 => '0',
		6588 => '0',
		6589 => '0',
		6590 => '0',
		6591 => '0',
		6592 => '0',
		6593 => '1',
		6594 => '1',
		6595 => '1',
		6596 => '0',
		6597 => '0',
		6598 => '1',
		6599 => '1',
		6600 => '1',
		6601 => '0',
		6602 => '0',
		6603 => '1',
		6604 => '1',
		6605 => '1',
		6606 => '0',
		6607 => '0',
		6608 => '1',
		6609 => '1',
		6610 => '1',
		6611 => '0',
		6612 => '0',
		6613 => '0',
		6614 => '0',
		6615 => '0',
		6616 => '0',
		6617 => '0',
		6618 => '1',
		6619 => '1',
		6620 => '1',
		6621 => '0',
		6622 => '0',
		6623 => '1',
		6624 => '1',
		6625 => '1',
		6626 => '0',
		6627 => '0',
		6628 => '0',
		6629 => '0',
		6630 => '0',
		6631 => '0',
		6632 => '0',
		6633 => '1',
		6634 => '1',
		6635 => '1',
		6636 => '0',
		6637 => '0',
		6638 => '1',
		6639 => '1',
		6640 => '1',
		6641 => '0',
		6642 => '0',
		6643 => '1',
		6644 => '1',
		6645 => '1',
		6646 => '0',
		6647 => '0',
		6656 => '1',
		6657 => '1',
		6658 => '1',
		6659 => '0',
		6660 => '0',
		6661 => '1',
		6662 => '1',
		6663 => '1',
		6664 => '0',
		6665 => '0',
		6666 => '1',
		6667 => '1',
		6668 => '1',
		6669 => '0',
		6670 => '0',
		6671 => '1',
		6672 => '1',
		6673 => '1',
		6674 => '0',
		6675 => '0',
		6676 => '1',
		6677 => '1',
		6678 => '1',
		6679 => '0',
		6680 => '0',
		6681 => '1',
		6682 => '1',
		6683 => '1',
		6684 => '0',
		6685 => '0',
		6686 => '0',
		6687 => '0',
		6688 => '0',
		6689 => '0',
		6690 => '0',
		6691 => '1',
		6692 => '1',
		6693 => '1',
		6694 => '0',
		6695 => '0',
		6696 => '1',
		6697 => '1',
		6698 => '1',
		6699 => '0',
		6700 => '0',
		6701 => '0',
		6702 => '0',
		6703 => '0',
		6704 => '0',
		6705 => '0',
		6706 => '1',
		6707 => '1',
		6708 => '1',
		6709 => '0',
		6710 => '0',
		6711 => '1',
		6712 => '1',
		6713 => '1',
		6714 => '0',
		6715 => '0',
		6716 => '0',
		6717 => '0',
		6718 => '0',
		6719 => '0',
		6720 => '0',
		6721 => '1',
		6722 => '1',
		6723 => '1',
		6724 => '0',
		6725 => '0',
		6726 => '1',
		6727 => '1',
		6728 => '1',
		6729 => '0',
		6730 => '0',
		6731 => '1',
		6732 => '1',
		6733 => '1',
		6734 => '0',
		6735 => '0',
		6736 => '1',
		6737 => '1',
		6738 => '1',
		6739 => '0',
		6740 => '0',
		6741 => '0',
		6742 => '0',
		6743 => '0',
		6744 => '0',
		6745 => '0',
		6746 => '1',
		6747 => '1',
		6748 => '1',
		6749 => '0',
		6750 => '0',
		6751 => '1',
		6752 => '1',
		6753 => '1',
		6754 => '0',
		6755 => '0',
		6756 => '0',
		6757 => '0',
		6758 => '0',
		6759 => '0',
		6760 => '0',
		6761 => '1',
		6762 => '1',
		6763 => '1',
		6764 => '0',
		6765 => '0',
		6766 => '1',
		6767 => '1',
		6768 => '1',
		6769 => '0',
		6770 => '0',
		6771 => '1',
		6772 => '1',
		6773 => '1',
		6774 => '0',
		6775 => '0',
		6784 => '1',
		6785 => '1',
		6786 => '1',
		6787 => '0',
		6788 => '0',
		6789 => '1',
		6790 => '1',
		6791 => '1',
		6792 => '0',
		6793 => '0',
		6794 => '1',
		6795 => '1',
		6796 => '1',
		6797 => '0',
		6798 => '0',
		6799 => '1',
		6800 => '1',
		6801 => '1',
		6802 => '0',
		6803 => '0',
		6804 => '1',
		6805 => '1',
		6806 => '1',
		6807 => '0',
		6808 => '0',
		6809 => '1',
		6810 => '1',
		6811 => '1',
		6812 => '0',
		6813 => '0',
		6814 => '0',
		6815 => '0',
		6816 => '0',
		6817 => '0',
		6818 => '0',
		6819 => '1',
		6820 => '1',
		6821 => '1',
		6822 => '0',
		6823 => '0',
		6824 => '1',
		6825 => '1',
		6826 => '1',
		6827 => '1',
		6828 => '1',
		6829 => '1',
		6830 => '0',
		6831 => '1',
		6832 => '1',
		6833 => '1',
		6834 => '1',
		6835 => '1',
		6836 => '1',
		6837 => '0',
		6838 => '0',
		6839 => '1',
		6840 => '1',
		6841 => '1',
		6842 => '0',
		6843 => '0',
		6844 => '0',
		6845 => '0',
		6846 => '0',
		6847 => '0',
		6848 => '0',
		6849 => '1',
		6850 => '1',
		6851 => '1',
		6852 => '0',
		6853 => '0',
		6854 => '1',
		6855 => '1',
		6856 => '1',
		6857 => '0',
		6858 => '0',
		6859 => '1',
		6860 => '1',
		6861 => '1',
		6862 => '0',
		6863 => '0',
		6864 => '1',
		6865 => '1',
		6866 => '1',
		6867 => '0',
		6868 => '0',
		6869 => '1',
		6870 => '1',
		6871 => '1',
		6872 => '0',
		6873 => '0',
		6874 => '1',
		6875 => '1',
		6876 => '1',
		6877 => '0',
		6878 => '0',
		6879 => '1',
		6880 => '1',
		6881 => '1',
		6882 => '0',
		6883 => '0',
		6884 => '1',
		6885 => '1',
		6886 => '1',
		6887 => '1',
		6888 => '1',
		6889 => '1',
		6890 => '1',
		6891 => '1',
		6892 => '0',
		6893 => '0',
		6894 => '1',
		6895 => '1',
		6896 => '1',
		6897 => '0',
		6898 => '0',
		6899 => '1',
		6900 => '1',
		6901 => '1',
		6902 => '0',
		6903 => '0',
		6912 => '1',
		6913 => '1',
		6914 => '1',
		6915 => '0',
		6916 => '0',
		6917 => '1',
		6918 => '1',
		6919 => '1',
		6920 => '0',
		6921 => '0',
		6922 => '1',
		6923 => '1',
		6924 => '1',
		6925 => '0',
		6926 => '0',
		6927 => '1',
		6928 => '1',
		6929 => '1',
		6930 => '0',
		6931 => '0',
		6932 => '1',
		6933 => '1',
		6934 => '1',
		6935 => '0',
		6936 => '0',
		6937 => '1',
		6938 => '1',
		6939 => '1',
		6940 => '0',
		6941 => '0',
		6942 => '1',
		6943 => '1',
		6944 => '1',
		6945 => '0',
		6946 => '0',
		6947 => '1',
		6948 => '1',
		6949 => '1',
		6950 => '0',
		6951 => '0',
		6952 => '1',
		6953 => '1',
		6954 => '1',
		6955 => '1',
		6956 => '1',
		6957 => '1',
		6958 => '0',
		6959 => '1',
		6960 => '1',
		6961 => '1',
		6962 => '1',
		6963 => '1',
		6964 => '1',
		6965 => '0',
		6966 => '0',
		6967 => '1',
		6968 => '1',
		6969 => '1',
		6970 => '0',
		6971 => '0',
		6972 => '1',
		6973 => '1',
		6974 => '1',
		6975 => '0',
		6976 => '0',
		6977 => '1',
		6978 => '1',
		6979 => '1',
		6980 => '0',
		6981 => '0',
		6982 => '1',
		6983 => '1',
		6984 => '1',
		6985 => '0',
		6986 => '0',
		6987 => '1',
		6988 => '1',
		6989 => '1',
		6990 => '0',
		6991 => '0',
		6992 => '1',
		6993 => '1',
		6994 => '1',
		6995 => '0',
		6996 => '0',
		6997 => '1',
		6998 => '1',
		6999 => '1',
		7000 => '0',
		7001 => '0',
		7002 => '1',
		7003 => '1',
		7004 => '1',
		7005 => '0',
		7006 => '0',
		7007 => '1',
		7008 => '1',
		7009 => '1',
		7010 => '0',
		7011 => '0',
		7012 => '1',
		7013 => '1',
		7014 => '1',
		7015 => '1',
		7016 => '1',
		7017 => '1',
		7018 => '1',
		7019 => '1',
		7020 => '0',
		7021 => '0',
		7022 => '1',
		7023 => '1',
		7024 => '1',
		7025 => '0',
		7026 => '0',
		7027 => '1',
		7028 => '1',
		7029 => '1',
		7030 => '0',
		7031 => '0',
		7040 => '1',
		7041 => '1',
		7042 => '1',
		7043 => '0',
		7044 => '0',
		7045 => '1',
		7046 => '1',
		7047 => '1',
		7048 => '0',
		7049 => '0',
		7050 => '1',
		7051 => '1',
		7052 => '1',
		7053 => '0',
		7054 => '0',
		7055 => '1',
		7056 => '1',
		7057 => '1',
		7058 => '0',
		7059 => '0',
		7060 => '1',
		7061 => '1',
		7062 => '1',
		7063 => '0',
		7064 => '0',
		7065 => '1',
		7066 => '1',
		7067 => '1',
		7068 => '0',
		7069 => '0',
		7070 => '1',
		7071 => '1',
		7072 => '1',
		7073 => '0',
		7074 => '0',
		7075 => '1',
		7076 => '1',
		7077 => '1',
		7078 => '0',
		7079 => '0',
		7080 => '1',
		7081 => '1',
		7082 => '1',
		7083 => '1',
		7084 => '1',
		7085 => '1',
		7086 => '0',
		7087 => '1',
		7088 => '1',
		7089 => '1',
		7090 => '1',
		7091 => '1',
		7092 => '1',
		7093 => '0',
		7094 => '0',
		7095 => '1',
		7096 => '1',
		7097 => '1',
		7098 => '0',
		7099 => '0',
		7100 => '1',
		7101 => '1',
		7102 => '1',
		7103 => '0',
		7104 => '0',
		7105 => '1',
		7106 => '1',
		7107 => '1',
		7108 => '0',
		7109 => '0',
		7110 => '1',
		7111 => '1',
		7112 => '1',
		7113 => '0',
		7114 => '0',
		7115 => '1',
		7116 => '1',
		7117 => '1',
		7118 => '0',
		7119 => '0',
		7120 => '1',
		7121 => '1',
		7122 => '1',
		7123 => '0',
		7124 => '0',
		7125 => '1',
		7126 => '1',
		7127 => '1',
		7128 => '0',
		7129 => '0',
		7130 => '1',
		7131 => '1',
		7132 => '1',
		7133 => '0',
		7134 => '0',
		7135 => '1',
		7136 => '1',
		7137 => '1',
		7138 => '0',
		7139 => '0',
		7140 => '1',
		7141 => '1',
		7142 => '1',
		7143 => '1',
		7144 => '1',
		7145 => '1',
		7146 => '1',
		7147 => '1',
		7148 => '0',
		7149 => '0',
		7150 => '1',
		7151 => '1',
		7152 => '1',
		7153 => '0',
		7154 => '0',
		7155 => '1',
		7156 => '1',
		7157 => '1',
		7158 => '0',
		7159 => '0',
		7168 => '1',
		7169 => '1',
		7170 => '1',
		7171 => '0',
		7172 => '0',
		7173 => '1',
		7174 => '1',
		7175 => '1',
		7176 => '0',
		7177 => '0',
		7178 => '1',
		7179 => '1',
		7180 => '1',
		7181 => '0',
		7182 => '0',
		7183 => '1',
		7184 => '1',
		7185 => '1',
		7186 => '0',
		7187 => '0',
		7188 => '1',
		7189 => '1',
		7190 => '1',
		7191 => '0',
		7192 => '0',
		7193 => '1',
		7194 => '1',
		7195 => '1',
		7196 => '0',
		7197 => '0',
		7198 => '1',
		7199 => '1',
		7200 => '1',
		7201 => '1',
		7202 => '1',
		7203 => '1',
		7204 => '1',
		7205 => '1',
		7206 => '0',
		7207 => '0',
		7208 => '0',
		7209 => '0',
		7210 => '0',
		7211 => '1',
		7212 => '1',
		7213 => '1',
		7214 => '0',
		7215 => '1',
		7216 => '1',
		7217 => '1',
		7218 => '0',
		7219 => '0',
		7220 => '0',
		7221 => '0',
		7222 => '0',
		7223 => '1',
		7224 => '1',
		7225 => '1',
		7226 => '0',
		7227 => '0',
		7228 => '1',
		7229 => '1',
		7230 => '1',
		7231 => '0',
		7232 => '0',
		7233 => '1',
		7234 => '1',
		7235 => '1',
		7236 => '0',
		7237 => '0',
		7238 => '1',
		7239 => '1',
		7240 => '1',
		7241 => '0',
		7242 => '0',
		7243 => '1',
		7244 => '1',
		7245 => '1',
		7246 => '0',
		7247 => '0',
		7248 => '1',
		7249 => '1',
		7250 => '1',
		7251 => '0',
		7252 => '0',
		7253 => '0',
		7254 => '0',
		7255 => '0',
		7256 => '1',
		7257 => '1',
		7258 => '1',
		7259 => '1',
		7260 => '1',
		7261 => '0',
		7262 => '0',
		7263 => '1',
		7264 => '1',
		7265 => '1',
		7266 => '0',
		7267 => '0',
		7268 => '0',
		7269 => '0',
		7270 => '0',
		7271 => '0',
		7272 => '0',
		7273 => '1',
		7274 => '1',
		7275 => '1',
		7276 => '0',
		7277 => '0',
		7278 => '1',
		7279 => '1',
		7280 => '1',
		7281 => '0',
		7282 => '0',
		7283 => '1',
		7284 => '1',
		7285 => '1',
		7286 => '0',
		7287 => '0',
		7296 => '1',
		7297 => '1',
		7298 => '1',
		7299 => '0',
		7300 => '0',
		7301 => '1',
		7302 => '1',
		7303 => '1',
		7304 => '0',
		7305 => '0',
		7306 => '1',
		7307 => '1',
		7308 => '1',
		7309 => '0',
		7310 => '0',
		7311 => '1',
		7312 => '1',
		7313 => '1',
		7314 => '0',
		7315 => '0',
		7316 => '1',
		7317 => '1',
		7318 => '1',
		7319 => '0',
		7320 => '0',
		7321 => '1',
		7322 => '1',
		7323 => '1',
		7324 => '0',
		7325 => '0',
		7326 => '1',
		7327 => '1',
		7328 => '1',
		7329 => '1',
		7330 => '1',
		7331 => '1',
		7332 => '1',
		7333 => '1',
		7334 => '0',
		7335 => '0',
		7336 => '0',
		7337 => '0',
		7338 => '0',
		7339 => '1',
		7340 => '1',
		7341 => '1',
		7342 => '0',
		7343 => '1',
		7344 => '1',
		7345 => '1',
		7346 => '0',
		7347 => '0',
		7348 => '0',
		7349 => '0',
		7350 => '0',
		7351 => '1',
		7352 => '1',
		7353 => '1',
		7354 => '0',
		7355 => '0',
		7356 => '1',
		7357 => '1',
		7358 => '1',
		7359 => '0',
		7360 => '0',
		7361 => '1',
		7362 => '1',
		7363 => '1',
		7364 => '0',
		7365 => '0',
		7366 => '1',
		7367 => '1',
		7368 => '1',
		7369 => '0',
		7370 => '0',
		7371 => '1',
		7372 => '1',
		7373 => '1',
		7374 => '0',
		7375 => '0',
		7376 => '1',
		7377 => '1',
		7378 => '1',
		7379 => '0',
		7380 => '0',
		7381 => '0',
		7382 => '0',
		7383 => '0',
		7384 => '1',
		7385 => '1',
		7386 => '1',
		7387 => '1',
		7388 => '1',
		7389 => '0',
		7390 => '0',
		7391 => '1',
		7392 => '1',
		7393 => '1',
		7394 => '0',
		7395 => '0',
		7396 => '0',
		7397 => '0',
		7398 => '0',
		7399 => '0',
		7400 => '0',
		7401 => '1',
		7402 => '1',
		7403 => '1',
		7404 => '0',
		7405 => '0',
		7406 => '1',
		7407 => '1',
		7408 => '1',
		7409 => '0',
		7410 => '0',
		7411 => '1',
		7412 => '1',
		7413 => '1',
		7414 => '0',
		7415 => '0',
		7424 => '1',
		7425 => '1',
		7426 => '1',
		7427 => '0',
		7428 => '0',
		7429 => '1',
		7430 => '1',
		7431 => '1',
		7432 => '0',
		7433 => '0',
		7434 => '1',
		7435 => '1',
		7436 => '1',
		7437 => '0',
		7438 => '0',
		7439 => '1',
		7440 => '1',
		7441 => '1',
		7442 => '0',
		7443 => '0',
		7444 => '1',
		7445 => '1',
		7446 => '1',
		7447 => '0',
		7448 => '0',
		7449 => '1',
		7450 => '1',
		7451 => '1',
		7452 => '0',
		7453 => '0',
		7454 => '1',
		7455 => '1',
		7456 => '1',
		7457 => '1',
		7458 => '1',
		7459 => '1',
		7460 => '1',
		7461 => '1',
		7462 => '0',
		7463 => '0',
		7464 => '0',
		7465 => '0',
		7466 => '0',
		7467 => '1',
		7468 => '1',
		7469 => '1',
		7470 => '0',
		7471 => '1',
		7472 => '1',
		7473 => '1',
		7474 => '0',
		7475 => '0',
		7476 => '0',
		7477 => '0',
		7478 => '0',
		7479 => '1',
		7480 => '1',
		7481 => '1',
		7482 => '0',
		7483 => '0',
		7484 => '1',
		7485 => '1',
		7486 => '1',
		7487 => '0',
		7488 => '0',
		7489 => '1',
		7490 => '1',
		7491 => '1',
		7492 => '0',
		7493 => '0',
		7494 => '1',
		7495 => '1',
		7496 => '1',
		7497 => '0',
		7498 => '0',
		7499 => '1',
		7500 => '1',
		7501 => '1',
		7502 => '0',
		7503 => '0',
		7504 => '1',
		7505 => '1',
		7506 => '1',
		7507 => '0',
		7508 => '0',
		7509 => '1',
		7510 => '1',
		7511 => '1',
		7512 => '1',
		7513 => '1',
		7514 => '1',
		7515 => '1',
		7516 => '1',
		7517 => '0',
		7518 => '0',
		7519 => '1',
		7520 => '1',
		7521 => '1',
		7522 => '0',
		7523 => '0',
		7524 => '1',
		7525 => '1',
		7526 => '1',
		7527 => '1',
		7528 => '1',
		7529 => '1',
		7530 => '1',
		7531 => '1',
		7532 => '0',
		7533 => '0',
		7534 => '1',
		7535 => '1',
		7536 => '1',
		7537 => '1',
		7538 => '1',
		7539 => '1',
		7540 => '1',
		7541 => '1',
		7542 => '0',
		7543 => '0',
		7552 => '1',
		7553 => '1',
		7554 => '1',
		7555 => '0',
		7556 => '0',
		7557 => '1',
		7558 => '1',
		7559 => '1',
		7560 => '0',
		7561 => '0',
		7562 => '1',
		7563 => '1',
		7564 => '1',
		7565 => '0',
		7566 => '0',
		7567 => '1',
		7568 => '1',
		7569 => '1',
		7570 => '0',
		7571 => '0',
		7572 => '1',
		7573 => '1',
		7574 => '1',
		7575 => '0',
		7576 => '0',
		7577 => '1',
		7578 => '1',
		7579 => '1',
		7580 => '0',
		7581 => '0',
		7582 => '1',
		7583 => '1',
		7584 => '1',
		7585 => '0',
		7586 => '0',
		7587 => '1',
		7588 => '1',
		7589 => '1',
		7590 => '0',
		7591 => '0',
		7592 => '0',
		7593 => '0',
		7594 => '0',
		7595 => '1',
		7596 => '1',
		7597 => '1',
		7598 => '0',
		7599 => '1',
		7600 => '1',
		7601 => '1',
		7602 => '0',
		7603 => '0',
		7604 => '0',
		7605 => '0',
		7606 => '0',
		7607 => '1',
		7608 => '1',
		7609 => '1',
		7610 => '0',
		7611 => '0',
		7612 => '1',
		7613 => '1',
		7614 => '1',
		7615 => '0',
		7616 => '0',
		7617 => '1',
		7618 => '1',
		7619 => '1',
		7620 => '0',
		7621 => '0',
		7622 => '1',
		7623 => '1',
		7624 => '1',
		7625 => '0',
		7626 => '0',
		7627 => '1',
		7628 => '1',
		7629 => '1',
		7630 => '0',
		7631 => '0',
		7632 => '1',
		7633 => '1',
		7634 => '1',
		7635 => '0',
		7636 => '0',
		7637 => '1',
		7638 => '1',
		7639 => '1',
		7640 => '0',
		7641 => '0',
		7642 => '1',
		7643 => '1',
		7644 => '1',
		7645 => '0',
		7646 => '0',
		7647 => '1',
		7648 => '1',
		7649 => '1',
		7650 => '0',
		7651 => '0',
		7652 => '1',
		7653 => '1',
		7654 => '1',
		7655 => '1',
		7656 => '1',
		7657 => '1',
		7658 => '1',
		7659 => '1',
		7660 => '0',
		7661 => '0',
		7662 => '1',
		7663 => '1',
		7664 => '1',
		7665 => '1',
		7666 => '1',
		7667 => '1',
		7668 => '1',
		7669 => '1',
		7670 => '0',
		7671 => '0',
		7680 => '1',
		7681 => '1',
		7682 => '1',
		7683 => '0',
		7684 => '0',
		7685 => '1',
		7686 => '1',
		7687 => '1',
		7688 => '0',
		7689 => '0',
		7690 => '1',
		7691 => '1',
		7692 => '1',
		7693 => '0',
		7694 => '0',
		7695 => '1',
		7696 => '1',
		7697 => '1',
		7698 => '0',
		7699 => '0',
		7700 => '1',
		7701 => '1',
		7702 => '1',
		7703 => '0',
		7704 => '0',
		7705 => '1',
		7706 => '1',
		7707 => '1',
		7708 => '0',
		7709 => '0',
		7710 => '1',
		7711 => '1',
		7712 => '1',
		7713 => '0',
		7714 => '0',
		7715 => '1',
		7716 => '1',
		7717 => '1',
		7718 => '0',
		7719 => '0',
		7720 => '0',
		7721 => '0',
		7722 => '0',
		7723 => '1',
		7724 => '1',
		7725 => '1',
		7726 => '0',
		7727 => '1',
		7728 => '1',
		7729 => '1',
		7730 => '0',
		7731 => '0',
		7732 => '0',
		7733 => '0',
		7734 => '0',
		7735 => '1',
		7736 => '1',
		7737 => '1',
		7738 => '0',
		7739 => '0',
		7740 => '1',
		7741 => '1',
		7742 => '1',
		7743 => '0',
		7744 => '0',
		7745 => '1',
		7746 => '1',
		7747 => '1',
		7748 => '0',
		7749 => '0',
		7750 => '1',
		7751 => '1',
		7752 => '1',
		7753 => '0',
		7754 => '0',
		7755 => '1',
		7756 => '1',
		7757 => '1',
		7758 => '0',
		7759 => '0',
		7760 => '1',
		7761 => '1',
		7762 => '1',
		7763 => '0',
		7764 => '0',
		7765 => '1',
		7766 => '1',
		7767 => '1',
		7768 => '0',
		7769 => '0',
		7770 => '1',
		7771 => '1',
		7772 => '1',
		7773 => '0',
		7774 => '0',
		7775 => '1',
		7776 => '1',
		7777 => '1',
		7778 => '0',
		7779 => '0',
		7780 => '1',
		7781 => '1',
		7782 => '1',
		7783 => '1',
		7784 => '1',
		7785 => '1',
		7786 => '1',
		7787 => '1',
		7788 => '0',
		7789 => '0',
		7790 => '1',
		7791 => '1',
		7792 => '1',
		7793 => '1',
		7794 => '1',
		7795 => '1',
		7796 => '1',
		7797 => '1',
		7798 => '0',
		7799 => '0',
		7808 => '1',
		7809 => '1',
		7810 => '1',
		7811 => '1',
		7812 => '1',
		7813 => '0',
		7814 => '0',
		7815 => '0',
		7816 => '1',
		7817 => '1',
		7818 => '1',
		7819 => '1',
		7820 => '1',
		7821 => '0',
		7822 => '0',
		7823 => '1',
		7824 => '1',
		7825 => '1',
		7826 => '0',
		7827 => '0',
		7828 => '1',
		7829 => '1',
		7830 => '1',
		7831 => '0',
		7832 => '0',
		7833 => '1',
		7834 => '1',
		7835 => '1',
		7836 => '0',
		7837 => '0',
		7838 => '0',
		7839 => '0',
		7840 => '0',
		7841 => '0',
		7842 => '0',
		7843 => '1',
		7844 => '1',
		7845 => '1',
		7846 => '0',
		7847 => '0',
		7848 => '0',
		7849 => '0',
		7850 => '0',
		7851 => '1',
		7852 => '1',
		7853 => '1',
		7854 => '0',
		7855 => '1',
		7856 => '1',
		7857 => '1',
		7858 => '0',
		7859 => '0',
		7860 => '0',
		7861 => '0',
		7862 => '0',
		7863 => '1',
		7864 => '1',
		7865 => '1',
		7866 => '0',
		7867 => '0',
		7868 => '0',
		7869 => '0',
		7870 => '0',
		7871 => '0',
		7872 => '0',
		7873 => '1',
		7874 => '1',
		7875 => '1',
		7876 => '0',
		7877 => '0',
		7878 => '1',
		7879 => '1',
		7880 => '1',
		7881 => '0',
		7882 => '0',
		7883 => '1',
		7884 => '1',
		7885 => '1',
		7886 => '0',
		7887 => '0',
		7888 => '1',
		7889 => '1',
		7890 => '1',
		7891 => '0',
		7892 => '0',
		7893 => '1',
		7894 => '1',
		7895 => '1',
		7896 => '0',
		7897 => '0',
		7898 => '1',
		7899 => '1',
		7900 => '1',
		7901 => '0',
		7902 => '0',
		7903 => '1',
		7904 => '1',
		7905 => '1',
		7906 => '0',
		7907 => '0',
		7908 => '0',
		7909 => '0',
		7910 => '0',
		7911 => '0',
		7912 => '0',
		7913 => '1',
		7914 => '1',
		7915 => '1',
		7916 => '0',
		7917 => '0',
		7918 => '1',
		7919 => '1',
		7920 => '1',
		7921 => '0',
		7922 => '0',
		7923 => '1',
		7924 => '1',
		7925 => '1',
		7926 => '0',
		7927 => '0',
		7936 => '1',
		7937 => '1',
		7938 => '1',
		7939 => '1',
		7940 => '1',
		7941 => '0',
		7942 => '0',
		7943 => '0',
		7944 => '1',
		7945 => '1',
		7946 => '1',
		7947 => '1',
		7948 => '1',
		7949 => '0',
		7950 => '0',
		7951 => '1',
		7952 => '1',
		7953 => '1',
		7954 => '0',
		7955 => '0',
		7956 => '1',
		7957 => '1',
		7958 => '1',
		7959 => '0',
		7960 => '0',
		7961 => '1',
		7962 => '1',
		7963 => '1',
		7964 => '0',
		7965 => '0',
		7966 => '0',
		7967 => '0',
		7968 => '0',
		7969 => '0',
		7970 => '0',
		7971 => '1',
		7972 => '1',
		7973 => '1',
		7974 => '0',
		7975 => '0',
		7976 => '0',
		7977 => '0',
		7978 => '0',
		7979 => '1',
		7980 => '1',
		7981 => '1',
		7982 => '0',
		7983 => '1',
		7984 => '1',
		7985 => '1',
		7986 => '0',
		7987 => '0',
		7988 => '0',
		7989 => '0',
		7990 => '0',
		7991 => '1',
		7992 => '1',
		7993 => '1',
		7994 => '0',
		7995 => '0',
		7996 => '0',
		7997 => '0',
		7998 => '0',
		7999 => '0',
		8000 => '0',
		8001 => '1',
		8002 => '1',
		8003 => '1',
		8004 => '0',
		8005 => '0',
		8006 => '1',
		8007 => '1',
		8008 => '1',
		8009 => '0',
		8010 => '0',
		8011 => '1',
		8012 => '1',
		8013 => '1',
		8014 => '0',
		8015 => '0',
		8016 => '1',
		8017 => '1',
		8018 => '1',
		8019 => '0',
		8020 => '0',
		8021 => '1',
		8022 => '1',
		8023 => '1',
		8024 => '0',
		8025 => '0',
		8026 => '1',
		8027 => '1',
		8028 => '1',
		8029 => '0',
		8030 => '0',
		8031 => '1',
		8032 => '1',
		8033 => '1',
		8034 => '0',
		8035 => '0',
		8036 => '0',
		8037 => '0',
		8038 => '0',
		8039 => '0',
		8040 => '0',
		8041 => '1',
		8042 => '1',
		8043 => '1',
		8044 => '0',
		8045 => '0',
		8046 => '1',
		8047 => '1',
		8048 => '1',
		8049 => '0',
		8050 => '0',
		8051 => '1',
		8052 => '1',
		8053 => '1',
		8054 => '0',
		8055 => '0',
		8064 => '0',
		8065 => '0',
		8066 => '0',
		8067 => '1',
		8068 => '1',
		8069 => '1',
		8070 => '1',
		8071 => '1',
		8072 => '1',
		8073 => '1',
		8074 => '0',
		8075 => '0',
		8076 => '0',
		8077 => '0',
		8078 => '0',
		8079 => '1',
		8080 => '1',
		8081 => '1',
		8082 => '1',
		8083 => '1',
		8084 => '1',
		8085 => '1',
		8086 => '1',
		8087 => '0',
		8088 => '0',
		8089 => '1',
		8090 => '1',
		8091 => '1',
		8092 => '1',
		8093 => '1',
		8094 => '1',
		8095 => '1',
		8096 => '1',
		8097 => '1',
		8098 => '1',
		8099 => '1',
		8100 => '1',
		8101 => '1',
		8102 => '0',
		8103 => '0',
		8104 => '0',
		8105 => '0',
		8106 => '0',
		8107 => '1',
		8108 => '1',
		8109 => '1',
		8110 => '1',
		8111 => '1',
		8112 => '1',
		8113 => '1',
		8114 => '0',
		8115 => '0',
		8116 => '0',
		8117 => '0',
		8118 => '0',
		8119 => '1',
		8120 => '1',
		8121 => '1',
		8122 => '1',
		8123 => '1',
		8124 => '1',
		8125 => '1',
		8126 => '1',
		8127 => '1',
		8128 => '1',
		8129 => '1',
		8130 => '1',
		8131 => '1',
		8132 => '0',
		8133 => '0',
		8134 => '1',
		8135 => '1',
		8136 => '1',
		8137 => '1',
		8138 => '1',
		8139 => '1',
		8140 => '1',
		8141 => '1',
		8142 => '0',
		8143 => '0',
		8144 => '1',
		8145 => '1',
		8146 => '1',
		8147 => '1',
		8148 => '1',
		8149 => '1',
		8150 => '1',
		8151 => '1',
		8152 => '1',
		8153 => '1',
		8154 => '1',
		8155 => '1',
		8156 => '1',
		8157 => '0',
		8158 => '0',
		8159 => '1',
		8160 => '1',
		8161 => '1',
		8162 => '1',
		8163 => '1',
		8164 => '1',
		8165 => '1',
		8166 => '1',
		8167 => '1',
		8168 => '1',
		8169 => '1',
		8170 => '1',
		8171 => '1',
		8172 => '0',
		8173 => '0',
		8174 => '1',
		8175 => '1',
		8176 => '1',
		8177 => '1',
		8178 => '1',
		8179 => '1',
		8180 => '1',
		8181 => '1',
		8182 => '0',
		8183 => '0',
		8192 => '0',
		8193 => '0',
		8194 => '0',
		8195 => '1',
		8196 => '1',
		8197 => '1',
		8198 => '1',
		8199 => '1',
		8200 => '1',
		8201 => '1',
		8202 => '0',
		8203 => '0',
		8204 => '0',
		8205 => '0',
		8206 => '0',
		8207 => '1',
		8208 => '1',
		8209 => '1',
		8210 => '1',
		8211 => '1',
		8212 => '1',
		8213 => '1',
		8214 => '1',
		8215 => '0',
		8216 => '0',
		8217 => '1',
		8218 => '1',
		8219 => '1',
		8220 => '1',
		8221 => '1',
		8222 => '1',
		8223 => '1',
		8224 => '1',
		8225 => '1',
		8226 => '1',
		8227 => '1',
		8228 => '1',
		8229 => '1',
		8230 => '0',
		8231 => '0',
		8232 => '0',
		8233 => '0',
		8234 => '0',
		8235 => '1',
		8236 => '1',
		8237 => '1',
		8238 => '1',
		8239 => '1',
		8240 => '1',
		8241 => '1',
		8242 => '0',
		8243 => '0',
		8244 => '0',
		8245 => '0',
		8246 => '0',
		8247 => '1',
		8248 => '1',
		8249 => '1',
		8250 => '1',
		8251 => '1',
		8252 => '1',
		8253 => '1',
		8254 => '1',
		8255 => '1',
		8256 => '1',
		8257 => '1',
		8258 => '1',
		8259 => '1',
		8260 => '0',
		8261 => '0',
		8262 => '1',
		8263 => '1',
		8264 => '1',
		8265 => '1',
		8266 => '1',
		8267 => '1',
		8268 => '1',
		8269 => '1',
		8270 => '0',
		8271 => '0',
		8272 => '1',
		8273 => '1',
		8274 => '1',
		8275 => '1',
		8276 => '1',
		8277 => '1',
		8278 => '1',
		8279 => '1',
		8280 => '1',
		8281 => '1',
		8282 => '1',
		8283 => '1',
		8284 => '1',
		8285 => '0',
		8286 => '0',
		8287 => '1',
		8288 => '1',
		8289 => '1',
		8290 => '1',
		8291 => '1',
		8292 => '1',
		8293 => '1',
		8294 => '1',
		8295 => '1',
		8296 => '1',
		8297 => '1',
		8298 => '1',
		8299 => '1',
		8300 => '0',
		8301 => '0',
		8302 => '1',
		8303 => '1',
		8304 => '1',
		8305 => '1',
		8306 => '1',
		8307 => '1',
		8308 => '1',
		8309 => '1',
		8310 => '0',
		8311 => '0',
		8320 => '0',
		8321 => '0',
		8322 => '0',
		8323 => '1',
		8324 => '1',
		8325 => '1',
		8326 => '1',
		8327 => '1',
		8328 => '1',
		8329 => '1',
		8330 => '0',
		8331 => '0',
		8332 => '0',
		8333 => '0',
		8334 => '0',
		8335 => '1',
		8336 => '1',
		8337 => '1',
		8338 => '1',
		8339 => '1',
		8340 => '1',
		8341 => '1',
		8342 => '1',
		8343 => '0',
		8344 => '0',
		8345 => '1',
		8346 => '1',
		8347 => '1',
		8348 => '1',
		8349 => '1',
		8350 => '1',
		8351 => '1',
		8352 => '1',
		8353 => '1',
		8354 => '1',
		8355 => '1',
		8356 => '1',
		8357 => '1',
		8358 => '0',
		8359 => '0',
		8360 => '0',
		8361 => '0',
		8362 => '0',
		8363 => '1',
		8364 => '1',
		8365 => '1',
		8366 => '1',
		8367 => '1',
		8368 => '1',
		8369 => '1',
		8370 => '0',
		8371 => '0',
		8372 => '0',
		8373 => '0',
		8374 => '0',
		8375 => '1',
		8376 => '1',
		8377 => '1',
		8378 => '1',
		8379 => '1',
		8380 => '1',
		8381 => '1',
		8382 => '1',
		8383 => '1',
		8384 => '1',
		8385 => '1',
		8386 => '1',
		8387 => '1',
		8388 => '0',
		8389 => '0',
		8390 => '1',
		8391 => '1',
		8392 => '1',
		8393 => '1',
		8394 => '1',
		8395 => '1',
		8396 => '1',
		8397 => '1',
		8398 => '0',
		8399 => '0',
		8400 => '1',
		8401 => '1',
		8402 => '1',
		8403 => '1',
		8404 => '1',
		8405 => '1',
		8406 => '1',
		8407 => '1',
		8408 => '1',
		8409 => '1',
		8410 => '1',
		8411 => '1',
		8412 => '1',
		8413 => '0',
		8414 => '0',
		8415 => '1',
		8416 => '1',
		8417 => '1',
		8418 => '1',
		8419 => '1',
		8420 => '1',
		8421 => '1',
		8422 => '1',
		8423 => '1',
		8424 => '1',
		8425 => '1',
		8426 => '1',
		8427 => '1',
		8428 => '0',
		8429 => '0',
		8430 => '1',
		8431 => '1',
		8432 => '1',
		8433 => '1',
		8434 => '1',
		8435 => '1',
		8436 => '1',
		8437 => '1',
		8438 => '0',
		8439 => '0',
		8448 => '0',
		8449 => '0',
		8450 => '0',
		8451 => '0',
		8452 => '0',
		8453 => '0',
		8454 => '0',
		8455 => '0',
		8456 => '0',
		8457 => '0',
		8458 => '0',
		8459 => '0',
		8460 => '0',
		8461 => '0',
		8462 => '0',
		8463 => '0',
		8464 => '0',
		8465 => '0',
		8466 => '0',
		8467 => '0',
		8468 => '0',
		8469 => '0',
		8470 => '0',
		8471 => '0',
		8472 => '0',
		8473 => '0',
		8474 => '0',
		8475 => '0',
		8476 => '0',
		8477 => '0',
		8478 => '0',
		8479 => '0',
		8480 => '0',
		8481 => '0',
		8482 => '0',
		8483 => '0',
		8484 => '0',
		8485 => '0',
		8486 => '0',
		8487 => '0',
		8488 => '0',
		8489 => '0',
		8490 => '0',
		8491 => '0',
		8492 => '0',
		8493 => '0',
		8494 => '0',
		8495 => '0',
		8496 => '0',
		8497 => '0',
		8498 => '0',
		8499 => '0',
		8500 => '0',
		8501 => '0',
		8502 => '0',
		8503 => '0',
		8504 => '0',
		8505 => '0',
		8506 => '0',
		8507 => '0',
		8508 => '0',
		8509 => '0',
		8510 => '0',
		8511 => '0',
		8512 => '0',
		8513 => '0',
		8514 => '0',
		8515 => '0',
		8516 => '0',
		8517 => '0',
		8518 => '0',
		8519 => '0',
		8520 => '0',
		8521 => '0',
		8522 => '0',
		8523 => '0',
		8524 => '0',
		8525 => '0',
		8526 => '0',
		8527 => '0',
		8528 => '0',
		8529 => '0',
		8530 => '0',
		8531 => '0',
		8532 => '0',
		8533 => '0',
		8534 => '0',
		8535 => '0',
		8536 => '0',
		8537 => '0',
		8538 => '0',
		8539 => '0',
		8540 => '0',
		8541 => '0',
		8542 => '0',
		8543 => '0',
		8544 => '0',
		8545 => '0',
		8546 => '0',
		8547 => '0',
		8548 => '0',
		8549 => '0',
		8550 => '0',
		8551 => '0',
		8552 => '0',
		8553 => '0',
		8554 => '0',
		8555 => '0',
		8556 => '0',
		8557 => '0',
		8558 => '0',
		8559 => '0',
		8560 => '0',
		8561 => '0',
		8562 => '0',
		8563 => '0',
		8564 => '0',
		8565 => '0',
		8566 => '0',
		8567 => '0',
		8576 => '0',
		8577 => '0',
		8578 => '0',
		8579 => '0',
		8580 => '0',
		8581 => '0',
		8582 => '0',
		8583 => '0',
		8584 => '0',
		8585 => '0',
		8586 => '0',
		8587 => '0',
		8588 => '0',
		8589 => '0',
		8590 => '0',
		8591 => '0',
		8592 => '0',
		8593 => '0',
		8594 => '0',
		8595 => '0',
		8596 => '0',
		8597 => '0',
		8598 => '0',
		8599 => '0',
		8600 => '0',
		8601 => '0',
		8602 => '0',
		8603 => '0',
		8604 => '0',
		8605 => '0',
		8606 => '0',
		8607 => '0',
		8608 => '0',
		8609 => '0',
		8610 => '0',
		8611 => '0',
		8612 => '0',
		8613 => '0',
		8614 => '0',
		8615 => '0',
		8616 => '0',
		8617 => '0',
		8618 => '0',
		8619 => '0',
		8620 => '0',
		8621 => '0',
		8622 => '0',
		8623 => '0',
		8624 => '0',
		8625 => '0',
		8626 => '0',
		8627 => '0',
		8628 => '0',
		8629 => '0',
		8630 => '0',
		8631 => '0',
		8632 => '0',
		8633 => '0',
		8634 => '0',
		8635 => '0',
		8636 => '0',
		8637 => '0',
		8638 => '0',
		8639 => '0',
		8640 => '0',
		8641 => '0',
		8642 => '0',
		8643 => '0',
		8644 => '0',
		8645 => '0',
		8646 => '0',
		8647 => '0',
		8648 => '0',
		8649 => '0',
		8650 => '0',
		8651 => '0',
		8652 => '0',
		8653 => '0',
		8654 => '0',
		8655 => '0',
		8656 => '0',
		8657 => '0',
		8658 => '0',
		8659 => '0',
		8660 => '0',
		8661 => '0',
		8662 => '0',
		8663 => '0',
		8664 => '0',
		8665 => '0',
		8666 => '0',
		8667 => '0',
		8668 => '0',
		8669 => '0',
		8670 => '0',
		8671 => '0',
		8672 => '0',
		8673 => '0',
		8674 => '0',
		8675 => '0',
		8676 => '0',
		8677 => '0',
		8678 => '0',
		8679 => '0',
		8680 => '0',
		8681 => '0',
		8682 => '0',
		8683 => '0',
		8684 => '0',
		8685 => '0',
		8686 => '0',
		8687 => '0',
		8688 => '0',
		8689 => '0',
		8690 => '0',
		8691 => '0',
		8692 => '0',
		8693 => '0',
		8694 => '0',
		8695 => '0',
		8704 => '0',
		8705 => '0',
		8706 => '0',
		8707 => '0',
		8708 => '0',
		8709 => '0',
		8710 => '0',
		8711 => '0',
		8712 => '0',
		8713 => '0',
		8714 => '0',
		8715 => '0',
		8716 => '0',
		8717 => '0',
		8718 => '0',
		8719 => '0',
		8720 => '0',
		8721 => '0',
		8722 => '0',
		8723 => '0',
		8724 => '0',
		8725 => '0',
		8726 => '0',
		8727 => '0',
		8728 => '0',
		8729 => '0',
		8730 => '0',
		8731 => '0',
		8732 => '0',
		8733 => '0',
		8734 => '0',
		8735 => '0',
		8736 => '0',
		8737 => '0',
		8738 => '0',
		8739 => '0',
		8740 => '0',
		8741 => '0',
		8742 => '0',
		8743 => '0',
		8744 => '0',
		8745 => '0',
		8746 => '0',
		8747 => '0',
		8748 => '0',
		8749 => '0',
		8750 => '0',
		8751 => '0',
		8752 => '0',
		8753 => '0',
		8754 => '0',
		8755 => '0',
		8756 => '0',
		8757 => '0',
		8758 => '0',
		8759 => '0',
		8760 => '0',
		8761 => '0',
		8762 => '0',
		8763 => '0',
		8764 => '0',
		8765 => '0',
		8766 => '0',
		8767 => '0',
		8768 => '0',
		8769 => '0',
		8770 => '0',
		8771 => '0',
		8772 => '0',
		8773 => '0',
		8774 => '0',
		8775 => '0',
		8776 => '0',
		8777 => '0',
		8778 => '0',
		8779 => '0',
		8780 => '0',
		8781 => '0',
		8782 => '0',
		8783 => '0',
		8784 => '0',
		8785 => '0',
		8786 => '0',
		8787 => '0',
		8788 => '0',
		8789 => '0',
		8790 => '0',
		8791 => '0',
		8792 => '0',
		8793 => '0',
		8794 => '0',
		8795 => '0',
		8796 => '0',
		8797 => '0',
		8798 => '0',
		8799 => '0',
		8800 => '0',
		8801 => '0',
		8802 => '0',
		8803 => '0',
		8804 => '0',
		8805 => '0',
		8806 => '0',
		8807 => '0',
		8808 => '0',
		8809 => '0',
		8810 => '0',
		8811 => '0',
		8812 => '0',
		8813 => '0',
		8814 => '0',
		8815 => '0',
		8816 => '0',
		8817 => '0',
		8818 => '0',
		8819 => '0',
		8820 => '0',
		8821 => '0',
		8822 => '0',
		8823 => '0',
		8832 => '0',
		8833 => '0',
		8834 => '0',
		8835 => '0',
		8836 => '0',
		8837 => '0',
		8838 => '0',
		8839 => '0',
		8840 => '0',
		8841 => '0',
		8842 => '0',
		8843 => '0',
		8844 => '0',
		8845 => '0',
		8846 => '0',
		8847 => '0',
		8848 => '0',
		8849 => '0',
		8850 => '0',
		8851 => '0',
		8852 => '0',
		8853 => '0',
		8854 => '0',
		8855 => '0',
		8856 => '0',
		8857 => '0',
		8858 => '0',
		8859 => '0',
		8860 => '0',
		8861 => '0',
		8862 => '0',
		8863 => '0',
		8864 => '0',
		8865 => '0',
		8866 => '0',
		8867 => '0',
		8868 => '0',
		8869 => '0',
		8870 => '0',
		8871 => '0',
		8872 => '0',
		8873 => '0',
		8874 => '0',
		8875 => '0',
		8876 => '0',
		8877 => '0',
		8878 => '0',
		8879 => '0',
		8880 => '0',
		8881 => '0',
		8882 => '0',
		8883 => '0',
		8884 => '0',
		8885 => '0',
		8886 => '0',
		8887 => '0',
		8888 => '0',
		8889 => '0',
		8890 => '0',
		8891 => '0',
		8892 => '0',
		8893 => '0',
		8894 => '0',
		8895 => '0',
		8896 => '0',
		8897 => '0',
		8898 => '0',
		8899 => '0',
		8900 => '0',
		8901 => '0',
		8902 => '0',
		8903 => '0',
		8904 => '0',
		8905 => '0',
		8906 => '0',
		8907 => '0',
		8908 => '0',
		8909 => '0',
		8910 => '0',
		8911 => '0',
		8912 => '0',
		8913 => '0',
		8914 => '0',
		8915 => '0',
		8916 => '0',
		8917 => '0',
		8918 => '0',
		8919 => '0',
		8920 => '0',
		8921 => '0',
		8922 => '0',
		8923 => '0',
		8924 => '0',
		8925 => '0',
		8926 => '0',
		8927 => '0',
		8928 => '0',
		8929 => '0',
		8930 => '0',
		8931 => '0',
		8932 => '0',
		8933 => '0',
		8934 => '0',
		8935 => '0',
		8936 => '0',
		8937 => '0',
		8938 => '0',
		8939 => '0',
		8940 => '0',
		8941 => '0',
		8942 => '0',
		8943 => '0',
		8944 => '0',
		8945 => '0',
		8946 => '0',
		8947 => '0',
		8948 => '0',
		8949 => '0',
		8950 => '0',
		8951 => '0',
		8960 => '0',
		8961 => '0',
		8962 => '0',
		8963 => '0',
		8964 => '0',
		8965 => '0',
		8966 => '0',
		8967 => '0',
		8968 => '0',
		8969 => '0',
		8970 => '0',
		8971 => '0',
		8972 => '0',
		8973 => '0',
		8974 => '0',
		8975 => '0',
		8976 => '0',
		8977 => '0',
		8978 => '0',
		8979 => '0',
		8980 => '0',
		8981 => '0',
		8982 => '0',
		8983 => '0',
		8984 => '0',
		8985 => '0',
		8986 => '0',
		8987 => '0',
		8988 => '0',
		8989 => '0',
		8990 => '0',
		8991 => '0',
		8992 => '0',
		8993 => '0',
		8994 => '0',
		8995 => '0',
		8996 => '0',
		8997 => '0',
		8998 => '0',
		8999 => '0',
		9000 => '0',
		9001 => '0',
		9002 => '0',
		9003 => '0',
		9004 => '0',
		9005 => '0',
		9006 => '0',
		9007 => '0',
		9008 => '0',
		9009 => '0',
		9010 => '0',
		9011 => '0',
		9012 => '0',
		9013 => '0',
		9014 => '0',
		9015 => '0',
		9016 => '0',
		9017 => '0',
		9018 => '0',
		9019 => '0',
		9020 => '0',
		9021 => '0',
		9022 => '0',
		9023 => '0',
		9024 => '0',
		9025 => '0',
		9026 => '0',
		9027 => '0',
		9028 => '0',
		9029 => '0',
		9030 => '0',
		9031 => '0',
		9032 => '0',
		9033 => '0',
		9034 => '0',
		9035 => '0',
		9036 => '0',
		9037 => '0',
		9038 => '0',
		9039 => '0',
		9040 => '0',
		9041 => '0',
		9042 => '0',
		9043 => '0',
		9044 => '0',
		9045 => '0',
		9046 => '0',
		9047 => '0',
		9048 => '0',
		9049 => '0',
		9050 => '0',
		9051 => '0',
		9052 => '0',
		9053 => '0',
		9054 => '0',
		9055 => '0',
		9056 => '0',
		9057 => '0',
		9058 => '0',
		9059 => '0',
		9060 => '0',
		9061 => '0',
		9062 => '0',
		9063 => '0',
		9064 => '0',
		9065 => '0',
		9066 => '0',
		9067 => '0',
		9068 => '0',
		9069 => '0',
		9070 => '0',
		9071 => '0',
		9072 => '0',
		9073 => '0',
		9074 => '0',
		9075 => '0',
		9076 => '0',
		9077 => '0',
		9078 => '0',
		9079 => '0',
		9088 => '0',
		9089 => '0',
		9090 => '0',
		9091 => '0',
		9092 => '0',
		9093 => '0',
		9094 => '0',
		9095 => '0',
		9096 => '0',
		9097 => '0',
		9098 => '0',
		9099 => '0',
		9100 => '0',
		9101 => '0',
		9102 => '0',
		9103 => '0',
		9104 => '0',
		9105 => '0',
		9106 => '0',
		9107 => '0',
		9108 => '0',
		9109 => '0',
		9110 => '0',
		9111 => '0',
		9112 => '0',
		9113 => '0',
		9114 => '0',
		9115 => '0',
		9116 => '0',
		9117 => '0',
		9118 => '0',
		9119 => '0',
		9120 => '0',
		9121 => '0',
		9122 => '0',
		9123 => '0',
		9124 => '0',
		9125 => '0',
		9126 => '0',
		9127 => '0',
		9128 => '0',
		9129 => '0',
		9130 => '0',
		9131 => '0',
		9132 => '0',
		9133 => '0',
		9134 => '0',
		9135 => '0',
		9136 => '0',
		9137 => '0',
		9138 => '0',
		9139 => '0',
		9140 => '0',
		9141 => '0',
		9142 => '0',
		9143 => '0',
		9144 => '0',
		9145 => '0',
		9146 => '0',
		9147 => '0',
		9148 => '0',
		9149 => '0',
		9150 => '0',
		9151 => '0',
		9152 => '0',
		9153 => '0',
		9154 => '0',
		9155 => '0',
		9156 => '0',
		9157 => '0',
		9158 => '0',
		9159 => '0',
		9160 => '0',
		9161 => '0',
		9162 => '0',
		9163 => '0',
		9164 => '0',
		9165 => '0',
		9166 => '0',
		9167 => '0',
		9168 => '0',
		9169 => '0',
		9170 => '0',
		9171 => '0',
		9172 => '0',
		9173 => '0',
		9174 => '0',
		9175 => '0',
		9176 => '0',
		9177 => '0',
		9178 => '0',
		9179 => '0',
		9180 => '0',
		9181 => '0',
		9182 => '0',
		9183 => '0',
		9184 => '0',
		9185 => '0',
		9186 => '0',
		9187 => '0',
		9188 => '0',
		9189 => '0',
		9190 => '0',
		9191 => '0',
		9192 => '0',
		9193 => '0',
		9194 => '0',
		9195 => '0',
		9196 => '0',
		9197 => '0',
		9198 => '0',
		9199 => '0',
		9200 => '0',
		9201 => '0',
		9202 => '0',
		9203 => '0',
		9204 => '0',
		9205 => '0',
		9206 => '0',
		9207 => '0',
		9216 => '1',
		9217 => '1',
		9218 => '1',
		9219 => '1',
		9220 => '1',
		9221 => '1',
		9222 => '1',
		9223 => '1',
		9224 => '1',
		9225 => '1',
		9226 => '1',
		9227 => '1',
		9228 => '1',
		9229 => '0',
		9230 => '0',
		9231 => '1',
		9232 => '1',
		9233 => '1',
		9234 => '1',
		9235 => '1',
		9236 => '1',
		9237 => '1',
		9238 => '1',
		9239 => '0',
		9240 => '0',
		9241 => '1',
		9242 => '1',
		9243 => '1',
		9244 => '1',
		9245 => '1',
		9246 => '1',
		9247 => '1',
		9248 => '1',
		9249 => '1',
		9250 => '1',
		9251 => '1',
		9252 => '1',
		9253 => '1',
		9254 => '0',
		9255 => '0',
		9256 => '1',
		9257 => '1',
		9258 => '1',
		9259 => '1',
		9260 => '1',
		9261 => '1',
		9262 => '1',
		9263 => '1',
		9264 => '1',
		9265 => '1',
		9266 => '1',
		9267 => '1',
		9268 => '1',
		9269 => '0',
		9270 => '0',
		9271 => '1',
		9272 => '1',
		9273 => '1',
		9274 => '1',
		9275 => '1',
		9276 => '1',
		9277 => '1',
		9278 => '1',
		9279 => '1',
		9280 => '1',
		9281 => '1',
		9282 => '1',
		9283 => '1',
		9284 => '0',
		9285 => '0',
		9286 => '1',
		9287 => '1',
		9288 => '1',
		9289 => '1',
		9290 => '1',
		9291 => '1',
		9292 => '1',
		9293 => '1',
		9294 => '0',
		9295 => '0',
		9296 => '1',
		9297 => '1',
		9298 => '1',
		9299 => '1',
		9300 => '1',
		9301 => '1',
		9302 => '1',
		9303 => '1',
		9304 => '1',
		9305 => '1',
		9306 => '1',
		9307 => '1',
		9308 => '1',
		9309 => '0',
		9310 => '0',
		9311 => '1',
		9312 => '1',
		9313 => '1',
		9314 => '1',
		9315 => '1',
		9316 => '1',
		9317 => '1',
		9318 => '1',
		9319 => '1',
		9320 => '1',
		9321 => '1',
		9322 => '1',
		9323 => '1',
		9324 => '0',
		9325 => '0',
		9326 => '1',
		9327 => '1',
		9328 => '1',
		9329 => '1',
		9330 => '1',
		9331 => '1',
		9332 => '1',
		9333 => '1',
		9334 => '0',
		9335 => '0',
		9344 => '1',
		9345 => '1',
		9346 => '1',
		9347 => '1',
		9348 => '1',
		9349 => '1',
		9350 => '1',
		9351 => '1',
		9352 => '1',
		9353 => '1',
		9354 => '1',
		9355 => '1',
		9356 => '1',
		9357 => '0',
		9358 => '0',
		9359 => '1',
		9360 => '1',
		9361 => '1',
		9362 => '1',
		9363 => '1',
		9364 => '1',
		9365 => '1',
		9366 => '1',
		9367 => '0',
		9368 => '0',
		9369 => '1',
		9370 => '1',
		9371 => '1',
		9372 => '1',
		9373 => '1',
		9374 => '1',
		9375 => '1',
		9376 => '1',
		9377 => '1',
		9378 => '1',
		9379 => '1',
		9380 => '1',
		9381 => '1',
		9382 => '0',
		9383 => '0',
		9384 => '1',
		9385 => '1',
		9386 => '1',
		9387 => '1',
		9388 => '1',
		9389 => '1',
		9390 => '1',
		9391 => '1',
		9392 => '1',
		9393 => '1',
		9394 => '1',
		9395 => '1',
		9396 => '1',
		9397 => '0',
		9398 => '0',
		9399 => '1',
		9400 => '1',
		9401 => '1',
		9402 => '1',
		9403 => '1',
		9404 => '1',
		9405 => '1',
		9406 => '1',
		9407 => '1',
		9408 => '1',
		9409 => '1',
		9410 => '1',
		9411 => '1',
		9412 => '0',
		9413 => '0',
		9414 => '1',
		9415 => '1',
		9416 => '1',
		9417 => '1',
		9418 => '1',
		9419 => '1',
		9420 => '1',
		9421 => '1',
		9422 => '0',
		9423 => '0',
		9424 => '1',
		9425 => '1',
		9426 => '1',
		9427 => '1',
		9428 => '1',
		9429 => '1',
		9430 => '1',
		9431 => '1',
		9432 => '1',
		9433 => '1',
		9434 => '1',
		9435 => '1',
		9436 => '1',
		9437 => '0',
		9438 => '0',
		9439 => '1',
		9440 => '1',
		9441 => '1',
		9442 => '1',
		9443 => '1',
		9444 => '1',
		9445 => '1',
		9446 => '1',
		9447 => '1',
		9448 => '1',
		9449 => '1',
		9450 => '1',
		9451 => '1',
		9452 => '0',
		9453 => '0',
		9454 => '1',
		9455 => '1',
		9456 => '1',
		9457 => '1',
		9458 => '1',
		9459 => '1',
		9460 => '1',
		9461 => '1',
		9462 => '0',
		9463 => '0',
		9472 => '1',
		9473 => '1',
		9474 => '1',
		9475 => '1',
		9476 => '1',
		9477 => '1',
		9478 => '1',
		9479 => '1',
		9480 => '1',
		9481 => '1',
		9482 => '1',
		9483 => '1',
		9484 => '1',
		9485 => '0',
		9486 => '0',
		9487 => '1',
		9488 => '1',
		9489 => '1',
		9490 => '1',
		9491 => '1',
		9492 => '1',
		9493 => '1',
		9494 => '1',
		9495 => '0',
		9496 => '0',
		9497 => '1',
		9498 => '1',
		9499 => '1',
		9500 => '1',
		9501 => '1',
		9502 => '1',
		9503 => '1',
		9504 => '1',
		9505 => '1',
		9506 => '1',
		9507 => '1',
		9508 => '1',
		9509 => '1',
		9510 => '0',
		9511 => '0',
		9512 => '1',
		9513 => '1',
		9514 => '1',
		9515 => '1',
		9516 => '1',
		9517 => '1',
		9518 => '1',
		9519 => '1',
		9520 => '1',
		9521 => '1',
		9522 => '1',
		9523 => '1',
		9524 => '1',
		9525 => '0',
		9526 => '0',
		9527 => '1',
		9528 => '1',
		9529 => '1',
		9530 => '1',
		9531 => '1',
		9532 => '1',
		9533 => '1',
		9534 => '1',
		9535 => '1',
		9536 => '1',
		9537 => '1',
		9538 => '1',
		9539 => '1',
		9540 => '0',
		9541 => '0',
		9542 => '1',
		9543 => '1',
		9544 => '1',
		9545 => '1',
		9546 => '1',
		9547 => '1',
		9548 => '1',
		9549 => '1',
		9550 => '0',
		9551 => '0',
		9552 => '1',
		9553 => '1',
		9554 => '1',
		9555 => '1',
		9556 => '1',
		9557 => '1',
		9558 => '1',
		9559 => '1',
		9560 => '1',
		9561 => '1',
		9562 => '1',
		9563 => '1',
		9564 => '1',
		9565 => '0',
		9566 => '0',
		9567 => '1',
		9568 => '1',
		9569 => '1',
		9570 => '1',
		9571 => '1',
		9572 => '1',
		9573 => '1',
		9574 => '1',
		9575 => '1',
		9576 => '1',
		9577 => '1',
		9578 => '1',
		9579 => '1',
		9580 => '0',
		9581 => '0',
		9582 => '1',
		9583 => '1',
		9584 => '1',
		9585 => '1',
		9586 => '1',
		9587 => '1',
		9588 => '1',
		9589 => '1',
		9590 => '0',
		9591 => '0',
		9600 => '1',
		9601 => '1',
		9602 => '1',
		9603 => '0',
		9604 => '0',
		9605 => '1',
		9606 => '1',
		9607 => '1',
		9608 => '0',
		9609 => '0',
		9610 => '1',
		9611 => '1',
		9612 => '1',
		9613 => '0',
		9614 => '0',
		9615 => '1',
		9616 => '1',
		9617 => '1',
		9618 => '0',
		9619 => '0',
		9620 => '1',
		9621 => '1',
		9622 => '1',
		9623 => '0',
		9624 => '0',
		9625 => '1',
		9626 => '1',
		9627 => '1',
		9628 => '0',
		9629 => '0',
		9630 => '0',
		9631 => '0',
		9632 => '0',
		9633 => '0',
		9634 => '0',
		9635 => '1',
		9636 => '1',
		9637 => '1',
		9638 => '0',
		9639 => '0',
		9640 => '1',
		9641 => '1',
		9642 => '1',
		9643 => '0',
		9644 => '0',
		9645 => '0',
		9646 => '0',
		9647 => '0',
		9648 => '0',
		9649 => '0',
		9650 => '1',
		9651 => '1',
		9652 => '1',
		9653 => '0',
		9654 => '0',
		9655 => '1',
		9656 => '1',
		9657 => '1',
		9658 => '0',
		9659 => '0',
		9660 => '0',
		9661 => '0',
		9662 => '0',
		9663 => '0',
		9664 => '0',
		9665 => '1',
		9666 => '1',
		9667 => '1',
		9668 => '0',
		9669 => '0',
		9670 => '1',
		9671 => '1',
		9672 => '1',
		9673 => '0',
		9674 => '0',
		9675 => '1',
		9676 => '1',
		9677 => '1',
		9678 => '0',
		9679 => '0',
		9680 => '1',
		9681 => '1',
		9682 => '1',
		9683 => '0',
		9684 => '0',
		9685 => '0',
		9686 => '0',
		9687 => '0',
		9688 => '0',
		9689 => '0',
		9690 => '1',
		9691 => '1',
		9692 => '1',
		9693 => '0',
		9694 => '0',
		9695 => '1',
		9696 => '1',
		9697 => '1',
		9698 => '0',
		9699 => '0',
		9700 => '0',
		9701 => '0',
		9702 => '0',
		9703 => '0',
		9704 => '0',
		9705 => '1',
		9706 => '1',
		9707 => '1',
		9708 => '0',
		9709 => '0',
		9710 => '1',
		9711 => '1',
		9712 => '1',
		9713 => '0',
		9714 => '0',
		9715 => '1',
		9716 => '1',
		9717 => '1',
		9718 => '0',
		9719 => '0',
		9728 => '1',
		9729 => '1',
		9730 => '1',
		9731 => '0',
		9732 => '0',
		9733 => '1',
		9734 => '1',
		9735 => '1',
		9736 => '0',
		9737 => '0',
		9738 => '1',
		9739 => '1',
		9740 => '1',
		9741 => '0',
		9742 => '0',
		9743 => '1',
		9744 => '1',
		9745 => '1',
		9746 => '0',
		9747 => '0',
		9748 => '1',
		9749 => '1',
		9750 => '1',
		9751 => '0',
		9752 => '0',
		9753 => '1',
		9754 => '1',
		9755 => '1',
		9756 => '0',
		9757 => '0',
		9758 => '0',
		9759 => '0',
		9760 => '0',
		9761 => '0',
		9762 => '0',
		9763 => '1',
		9764 => '1',
		9765 => '1',
		9766 => '0',
		9767 => '0',
		9768 => '1',
		9769 => '1',
		9770 => '1',
		9771 => '0',
		9772 => '0',
		9773 => '0',
		9774 => '0',
		9775 => '0',
		9776 => '0',
		9777 => '0',
		9778 => '1',
		9779 => '1',
		9780 => '1',
		9781 => '0',
		9782 => '0',
		9783 => '1',
		9784 => '1',
		9785 => '1',
		9786 => '0',
		9787 => '0',
		9788 => '0',
		9789 => '0',
		9790 => '0',
		9791 => '0',
		9792 => '0',
		9793 => '1',
		9794 => '1',
		9795 => '1',
		9796 => '0',
		9797 => '0',
		9798 => '1',
		9799 => '1',
		9800 => '1',
		9801 => '0',
		9802 => '0',
		9803 => '1',
		9804 => '1',
		9805 => '1',
		9806 => '0',
		9807 => '0',
		9808 => '1',
		9809 => '1',
		9810 => '1',
		9811 => '0',
		9812 => '0',
		9813 => '0',
		9814 => '0',
		9815 => '0',
		9816 => '0',
		9817 => '0',
		9818 => '1',
		9819 => '1',
		9820 => '1',
		9821 => '0',
		9822 => '0',
		9823 => '1',
		9824 => '1',
		9825 => '1',
		9826 => '0',
		9827 => '0',
		9828 => '0',
		9829 => '0',
		9830 => '0',
		9831 => '0',
		9832 => '0',
		9833 => '1',
		9834 => '1',
		9835 => '1',
		9836 => '0',
		9837 => '0',
		9838 => '1',
		9839 => '1',
		9840 => '1',
		9841 => '0',
		9842 => '0',
		9843 => '1',
		9844 => '1',
		9845 => '1',
		9846 => '0',
		9847 => '0',
		9856 => '1',
		9857 => '1',
		9858 => '1',
		9859 => '0',
		9860 => '0',
		9861 => '1',
		9862 => '1',
		9863 => '1',
		9864 => '0',
		9865 => '0',
		9866 => '1',
		9867 => '1',
		9868 => '1',
		9869 => '0',
		9870 => '0',
		9871 => '1',
		9872 => '1',
		9873 => '1',
		9874 => '0',
		9875 => '0',
		9876 => '1',
		9877 => '1',
		9878 => '1',
		9879 => '0',
		9880 => '0',
		9881 => '1',
		9882 => '1',
		9883 => '1',
		9884 => '0',
		9885 => '0',
		9886 => '0',
		9887 => '0',
		9888 => '0',
		9889 => '0',
		9890 => '0',
		9891 => '1',
		9892 => '1',
		9893 => '1',
		9894 => '0',
		9895 => '0',
		9896 => '1',
		9897 => '1',
		9898 => '1',
		9899 => '1',
		9900 => '1',
		9901 => '1',
		9902 => '0',
		9903 => '1',
		9904 => '1',
		9905 => '1',
		9906 => '1',
		9907 => '1',
		9908 => '1',
		9909 => '0',
		9910 => '0',
		9911 => '1',
		9912 => '1',
		9913 => '1',
		9914 => '0',
		9915 => '0',
		9916 => '0',
		9917 => '0',
		9918 => '0',
		9919 => '0',
		9920 => '0',
		9921 => '1',
		9922 => '1',
		9923 => '1',
		9924 => '0',
		9925 => '0',
		9926 => '1',
		9927 => '1',
		9928 => '1',
		9929 => '0',
		9930 => '0',
		9931 => '1',
		9932 => '1',
		9933 => '1',
		9934 => '0',
		9935 => '0',
		9936 => '1',
		9937 => '1',
		9938 => '1',
		9939 => '0',
		9940 => '0',
		9941 => '1',
		9942 => '1',
		9943 => '1',
		9944 => '0',
		9945 => '0',
		9946 => '1',
		9947 => '1',
		9948 => '1',
		9949 => '0',
		9950 => '0',
		9951 => '1',
		9952 => '1',
		9953 => '1',
		9954 => '0',
		9955 => '0',
		9956 => '1',
		9957 => '1',
		9958 => '1',
		9959 => '1',
		9960 => '1',
		9961 => '1',
		9962 => '1',
		9963 => '1',
		9964 => '0',
		9965 => '0',
		9966 => '1',
		9967 => '1',
		9968 => '1',
		9969 => '0',
		9970 => '0',
		9971 => '1',
		9972 => '1',
		9973 => '1',
		9974 => '0',
		9975 => '0',
		9984 => '1',
		9985 => '1',
		9986 => '1',
		9987 => '0',
		9988 => '0',
		9989 => '1',
		9990 => '1',
		9991 => '1',
		9992 => '0',
		9993 => '0',
		9994 => '1',
		9995 => '1',
		9996 => '1',
		9997 => '0',
		9998 => '0',
		9999 => '1',
		10000 => '1',
		10001 => '1',
		10002 => '0',
		10003 => '0',
		10004 => '1',
		10005 => '1',
		10006 => '1',
		10007 => '0',
		10008 => '0',
		10009 => '1',
		10010 => '1',
		10011 => '1',
		10012 => '0',
		10013 => '0',
		10014 => '1',
		10015 => '1',
		10016 => '1',
		10017 => '0',
		10018 => '0',
		10019 => '1',
		10020 => '1',
		10021 => '1',
		10022 => '0',
		10023 => '0',
		10024 => '1',
		10025 => '1',
		10026 => '1',
		10027 => '1',
		10028 => '1',
		10029 => '1',
		10030 => '0',
		10031 => '1',
		10032 => '1',
		10033 => '1',
		10034 => '1',
		10035 => '1',
		10036 => '1',
		10037 => '0',
		10038 => '0',
		10039 => '1',
		10040 => '1',
		10041 => '1',
		10042 => '0',
		10043 => '0',
		10044 => '1',
		10045 => '1',
		10046 => '1',
		10047 => '0',
		10048 => '0',
		10049 => '1',
		10050 => '1',
		10051 => '1',
		10052 => '0',
		10053 => '0',
		10054 => '1',
		10055 => '1',
		10056 => '1',
		10057 => '0',
		10058 => '0',
		10059 => '1',
		10060 => '1',
		10061 => '1',
		10062 => '0',
		10063 => '0',
		10064 => '1',
		10065 => '1',
		10066 => '1',
		10067 => '0',
		10068 => '0',
		10069 => '1',
		10070 => '1',
		10071 => '1',
		10072 => '0',
		10073 => '0',
		10074 => '1',
		10075 => '1',
		10076 => '1',
		10077 => '0',
		10078 => '0',
		10079 => '1',
		10080 => '1',
		10081 => '1',
		10082 => '0',
		10083 => '0',
		10084 => '1',
		10085 => '1',
		10086 => '1',
		10087 => '1',
		10088 => '1',
		10089 => '1',
		10090 => '1',
		10091 => '1',
		10092 => '0',
		10093 => '0',
		10094 => '1',
		10095 => '1',
		10096 => '1',
		10097 => '0',
		10098 => '0',
		10099 => '1',
		10100 => '1',
		10101 => '1',
		10102 => '0',
		10103 => '0',
		10112 => '1',
		10113 => '1',
		10114 => '1',
		10115 => '0',
		10116 => '0',
		10117 => '1',
		10118 => '1',
		10119 => '1',
		10120 => '0',
		10121 => '0',
		10122 => '1',
		10123 => '1',
		10124 => '1',
		10125 => '0',
		10126 => '0',
		10127 => '1',
		10128 => '1',
		10129 => '1',
		10130 => '0',
		10131 => '0',
		10132 => '1',
		10133 => '1',
		10134 => '1',
		10135 => '0',
		10136 => '0',
		10137 => '1',
		10138 => '1',
		10139 => '1',
		10140 => '0',
		10141 => '0',
		10142 => '1',
		10143 => '1',
		10144 => '1',
		10145 => '0',
		10146 => '0',
		10147 => '1',
		10148 => '1',
		10149 => '1',
		10150 => '0',
		10151 => '0',
		10152 => '1',
		10153 => '1',
		10154 => '1',
		10155 => '1',
		10156 => '1',
		10157 => '1',
		10158 => '0',
		10159 => '1',
		10160 => '1',
		10161 => '1',
		10162 => '1',
		10163 => '1',
		10164 => '1',
		10165 => '0',
		10166 => '0',
		10167 => '1',
		10168 => '1',
		10169 => '1',
		10170 => '0',
		10171 => '0',
		10172 => '1',
		10173 => '1',
		10174 => '1',
		10175 => '0',
		10176 => '0',
		10177 => '1',
		10178 => '1',
		10179 => '1',
		10180 => '0',
		10181 => '0',
		10182 => '1',
		10183 => '1',
		10184 => '1',
		10185 => '0',
		10186 => '0',
		10187 => '1',
		10188 => '1',
		10189 => '1',
		10190 => '0',
		10191 => '0',
		10192 => '1',
		10193 => '1',
		10194 => '1',
		10195 => '0',
		10196 => '0',
		10197 => '1',
		10198 => '1',
		10199 => '1',
		10200 => '0',
		10201 => '0',
		10202 => '1',
		10203 => '1',
		10204 => '1',
		10205 => '0',
		10206 => '0',
		10207 => '1',
		10208 => '1',
		10209 => '1',
		10210 => '0',
		10211 => '0',
		10212 => '1',
		10213 => '1',
		10214 => '1',
		10215 => '1',
		10216 => '1',
		10217 => '1',
		10218 => '1',
		10219 => '1',
		10220 => '0',
		10221 => '0',
		10222 => '1',
		10223 => '1',
		10224 => '1',
		10225 => '0',
		10226 => '0',
		10227 => '1',
		10228 => '1',
		10229 => '1',
		10230 => '0',
		10231 => '0',
		10240 => '1',
		10241 => '1',
		10242 => '1',
		10243 => '0',
		10244 => '0',
		10245 => '1',
		10246 => '1',
		10247 => '1',
		10248 => '0',
		10249 => '0',
		10250 => '1',
		10251 => '1',
		10252 => '1',
		10253 => '0',
		10254 => '0',
		10255 => '1',
		10256 => '1',
		10257 => '1',
		10258 => '0',
		10259 => '0',
		10260 => '1',
		10261 => '1',
		10262 => '1',
		10263 => '0',
		10264 => '0',
		10265 => '1',
		10266 => '1',
		10267 => '1',
		10268 => '0',
		10269 => '0',
		10270 => '1',
		10271 => '1',
		10272 => '1',
		10273 => '1',
		10274 => '1',
		10275 => '1',
		10276 => '1',
		10277 => '1',
		10278 => '0',
		10279 => '0',
		10280 => '0',
		10281 => '0',
		10282 => '0',
		10283 => '1',
		10284 => '1',
		10285 => '1',
		10286 => '0',
		10287 => '1',
		10288 => '1',
		10289 => '1',
		10290 => '0',
		10291 => '0',
		10292 => '0',
		10293 => '0',
		10294 => '0',
		10295 => '1',
		10296 => '1',
		10297 => '1',
		10298 => '0',
		10299 => '0',
		10300 => '1',
		10301 => '1',
		10302 => '1',
		10303 => '0',
		10304 => '0',
		10305 => '1',
		10306 => '1',
		10307 => '1',
		10308 => '0',
		10309 => '0',
		10310 => '1',
		10311 => '1',
		10312 => '1',
		10313 => '0',
		10314 => '0',
		10315 => '1',
		10316 => '1',
		10317 => '1',
		10318 => '0',
		10319 => '0',
		10320 => '1',
		10321 => '1',
		10322 => '1',
		10323 => '0',
		10324 => '0',
		10325 => '0',
		10326 => '0',
		10327 => '0',
		10328 => '1',
		10329 => '1',
		10330 => '1',
		10331 => '1',
		10332 => '1',
		10333 => '0',
		10334 => '0',
		10335 => '1',
		10336 => '1',
		10337 => '1',
		10338 => '0',
		10339 => '0',
		10340 => '0',
		10341 => '0',
		10342 => '0',
		10343 => '0',
		10344 => '0',
		10345 => '1',
		10346 => '1',
		10347 => '1',
		10348 => '0',
		10349 => '0',
		10350 => '1',
		10351 => '1',
		10352 => '1',
		10353 => '0',
		10354 => '0',
		10355 => '1',
		10356 => '1',
		10357 => '1',
		10358 => '0',
		10359 => '0',
		10368 => '1',
		10369 => '1',
		10370 => '1',
		10371 => '0',
		10372 => '0',
		10373 => '1',
		10374 => '1',
		10375 => '1',
		10376 => '0',
		10377 => '0',
		10378 => '1',
		10379 => '1',
		10380 => '1',
		10381 => '0',
		10382 => '0',
		10383 => '1',
		10384 => '1',
		10385 => '1',
		10386 => '0',
		10387 => '0',
		10388 => '1',
		10389 => '1',
		10390 => '1',
		10391 => '0',
		10392 => '0',
		10393 => '1',
		10394 => '1',
		10395 => '1',
		10396 => '0',
		10397 => '0',
		10398 => '1',
		10399 => '1',
		10400 => '1',
		10401 => '1',
		10402 => '1',
		10403 => '1',
		10404 => '1',
		10405 => '1',
		10406 => '0',
		10407 => '0',
		10408 => '0',
		10409 => '0',
		10410 => '0',
		10411 => '1',
		10412 => '1',
		10413 => '1',
		10414 => '0',
		10415 => '1',
		10416 => '1',
		10417 => '1',
		10418 => '0',
		10419 => '0',
		10420 => '0',
		10421 => '0',
		10422 => '0',
		10423 => '1',
		10424 => '1',
		10425 => '1',
		10426 => '0',
		10427 => '0',
		10428 => '1',
		10429 => '1',
		10430 => '1',
		10431 => '0',
		10432 => '0',
		10433 => '1',
		10434 => '1',
		10435 => '1',
		10436 => '0',
		10437 => '0',
		10438 => '1',
		10439 => '1',
		10440 => '1',
		10441 => '0',
		10442 => '0',
		10443 => '1',
		10444 => '1',
		10445 => '1',
		10446 => '0',
		10447 => '0',
		10448 => '1',
		10449 => '1',
		10450 => '1',
		10451 => '0',
		10452 => '0',
		10453 => '0',
		10454 => '0',
		10455 => '0',
		10456 => '1',
		10457 => '1',
		10458 => '1',
		10459 => '1',
		10460 => '1',
		10461 => '0',
		10462 => '0',
		10463 => '1',
		10464 => '1',
		10465 => '1',
		10466 => '0',
		10467 => '0',
		10468 => '0',
		10469 => '0',
		10470 => '0',
		10471 => '0',
		10472 => '0',
		10473 => '1',
		10474 => '1',
		10475 => '1',
		10476 => '0',
		10477 => '0',
		10478 => '1',
		10479 => '1',
		10480 => '1',
		10481 => '0',
		10482 => '0',
		10483 => '1',
		10484 => '1',
		10485 => '1',
		10486 => '0',
		10487 => '0',
		10496 => '1',
		10497 => '1',
		10498 => '1',
		10499 => '0',
		10500 => '0',
		10501 => '1',
		10502 => '1',
		10503 => '1',
		10504 => '0',
		10505 => '0',
		10506 => '1',
		10507 => '1',
		10508 => '1',
		10509 => '0',
		10510 => '0',
		10511 => '1',
		10512 => '1',
		10513 => '1',
		10514 => '0',
		10515 => '0',
		10516 => '1',
		10517 => '1',
		10518 => '1',
		10519 => '0',
		10520 => '0',
		10521 => '1',
		10522 => '1',
		10523 => '1',
		10524 => '0',
		10525 => '0',
		10526 => '1',
		10527 => '1',
		10528 => '1',
		10529 => '1',
		10530 => '1',
		10531 => '1',
		10532 => '1',
		10533 => '1',
		10534 => '0',
		10535 => '0',
		10536 => '0',
		10537 => '0',
		10538 => '0',
		10539 => '1',
		10540 => '1',
		10541 => '1',
		10542 => '0',
		10543 => '1',
		10544 => '1',
		10545 => '1',
		10546 => '0',
		10547 => '0',
		10548 => '0',
		10549 => '0',
		10550 => '0',
		10551 => '1',
		10552 => '1',
		10553 => '1',
		10554 => '0',
		10555 => '0',
		10556 => '1',
		10557 => '1',
		10558 => '1',
		10559 => '0',
		10560 => '0',
		10561 => '1',
		10562 => '1',
		10563 => '1',
		10564 => '0',
		10565 => '0',
		10566 => '1',
		10567 => '1',
		10568 => '1',
		10569 => '0',
		10570 => '0',
		10571 => '1',
		10572 => '1',
		10573 => '1',
		10574 => '0',
		10575 => '0',
		10576 => '1',
		10577 => '1',
		10578 => '1',
		10579 => '0',
		10580 => '0',
		10581 => '1',
		10582 => '1',
		10583 => '1',
		10584 => '1',
		10585 => '1',
		10586 => '1',
		10587 => '1',
		10588 => '1',
		10589 => '0',
		10590 => '0',
		10591 => '1',
		10592 => '1',
		10593 => '1',
		10594 => '0',
		10595 => '0',
		10596 => '1',
		10597 => '1',
		10598 => '1',
		10599 => '1',
		10600 => '1',
		10601 => '1',
		10602 => '1',
		10603 => '1',
		10604 => '0',
		10605 => '0',
		10606 => '1',
		10607 => '1',
		10608 => '1',
		10609 => '1',
		10610 => '1',
		10611 => '1',
		10612 => '1',
		10613 => '1',
		10614 => '0',
		10615 => '0',
		10624 => '1',
		10625 => '1',
		10626 => '1',
		10627 => '0',
		10628 => '0',
		10629 => '1',
		10630 => '1',
		10631 => '1',
		10632 => '0',
		10633 => '0',
		10634 => '1',
		10635 => '1',
		10636 => '1',
		10637 => '0',
		10638 => '0',
		10639 => '1',
		10640 => '1',
		10641 => '1',
		10642 => '0',
		10643 => '0',
		10644 => '1',
		10645 => '1',
		10646 => '1',
		10647 => '0',
		10648 => '0',
		10649 => '1',
		10650 => '1',
		10651 => '1',
		10652 => '0',
		10653 => '0',
		10654 => '1',
		10655 => '1',
		10656 => '1',
		10657 => '0',
		10658 => '0',
		10659 => '1',
		10660 => '1',
		10661 => '1',
		10662 => '0',
		10663 => '0',
		10664 => '0',
		10665 => '0',
		10666 => '0',
		10667 => '1',
		10668 => '1',
		10669 => '1',
		10670 => '0',
		10671 => '1',
		10672 => '1',
		10673 => '1',
		10674 => '0',
		10675 => '0',
		10676 => '0',
		10677 => '0',
		10678 => '0',
		10679 => '1',
		10680 => '1',
		10681 => '1',
		10682 => '0',
		10683 => '0',
		10684 => '1',
		10685 => '1',
		10686 => '1',
		10687 => '0',
		10688 => '0',
		10689 => '1',
		10690 => '1',
		10691 => '1',
		10692 => '0',
		10693 => '0',
		10694 => '1',
		10695 => '1',
		10696 => '1',
		10697 => '0',
		10698 => '0',
		10699 => '1',
		10700 => '1',
		10701 => '1',
		10702 => '0',
		10703 => '0',
		10704 => '1',
		10705 => '1',
		10706 => '1',
		10707 => '0',
		10708 => '0',
		10709 => '1',
		10710 => '1',
		10711 => '1',
		10712 => '0',
		10713 => '0',
		10714 => '1',
		10715 => '1',
		10716 => '1',
		10717 => '0',
		10718 => '0',
		10719 => '1',
		10720 => '1',
		10721 => '1',
		10722 => '0',
		10723 => '0',
		10724 => '1',
		10725 => '1',
		10726 => '1',
		10727 => '1',
		10728 => '1',
		10729 => '1',
		10730 => '1',
		10731 => '1',
		10732 => '0',
		10733 => '0',
		10734 => '1',
		10735 => '1',
		10736 => '1',
		10737 => '1',
		10738 => '1',
		10739 => '1',
		10740 => '1',
		10741 => '1',
		10742 => '0',
		10743 => '0',
		10752 => '1',
		10753 => '1',
		10754 => '1',
		10755 => '0',
		10756 => '0',
		10757 => '1',
		10758 => '1',
		10759 => '1',
		10760 => '0',
		10761 => '0',
		10762 => '1',
		10763 => '1',
		10764 => '1',
		10765 => '0',
		10766 => '0',
		10767 => '1',
		10768 => '1',
		10769 => '1',
		10770 => '0',
		10771 => '0',
		10772 => '1',
		10773 => '1',
		10774 => '1',
		10775 => '0',
		10776 => '0',
		10777 => '1',
		10778 => '1',
		10779 => '1',
		10780 => '0',
		10781 => '0',
		10782 => '1',
		10783 => '1',
		10784 => '1',
		10785 => '0',
		10786 => '0',
		10787 => '1',
		10788 => '1',
		10789 => '1',
		10790 => '0',
		10791 => '0',
		10792 => '0',
		10793 => '0',
		10794 => '0',
		10795 => '1',
		10796 => '1',
		10797 => '1',
		10798 => '0',
		10799 => '1',
		10800 => '1',
		10801 => '1',
		10802 => '0',
		10803 => '0',
		10804 => '0',
		10805 => '0',
		10806 => '0',
		10807 => '1',
		10808 => '1',
		10809 => '1',
		10810 => '0',
		10811 => '0',
		10812 => '1',
		10813 => '1',
		10814 => '1',
		10815 => '0',
		10816 => '0',
		10817 => '1',
		10818 => '1',
		10819 => '1',
		10820 => '0',
		10821 => '0',
		10822 => '1',
		10823 => '1',
		10824 => '1',
		10825 => '0',
		10826 => '0',
		10827 => '1',
		10828 => '1',
		10829 => '1',
		10830 => '0',
		10831 => '0',
		10832 => '1',
		10833 => '1',
		10834 => '1',
		10835 => '0',
		10836 => '0',
		10837 => '1',
		10838 => '1',
		10839 => '1',
		10840 => '0',
		10841 => '0',
		10842 => '1',
		10843 => '1',
		10844 => '1',
		10845 => '0',
		10846 => '0',
		10847 => '1',
		10848 => '1',
		10849 => '1',
		10850 => '0',
		10851 => '0',
		10852 => '1',
		10853 => '1',
		10854 => '1',
		10855 => '1',
		10856 => '1',
		10857 => '1',
		10858 => '1',
		10859 => '1',
		10860 => '0',
		10861 => '0',
		10862 => '1',
		10863 => '1',
		10864 => '1',
		10865 => '1',
		10866 => '1',
		10867 => '1',
		10868 => '1',
		10869 => '1',
		10870 => '0',
		10871 => '0',
		10880 => '1',
		10881 => '1',
		10882 => '1',
		10883 => '1',
		10884 => '1',
		10885 => '0',
		10886 => '0',
		10887 => '0',
		10888 => '1',
		10889 => '1',
		10890 => '1',
		10891 => '1',
		10892 => '1',
		10893 => '0',
		10894 => '0',
		10895 => '1',
		10896 => '1',
		10897 => '1',
		10898 => '0',
		10899 => '0',
		10900 => '1',
		10901 => '1',
		10902 => '1',
		10903 => '0',
		10904 => '0',
		10905 => '1',
		10906 => '1',
		10907 => '1',
		10908 => '0',
		10909 => '0',
		10910 => '0',
		10911 => '0',
		10912 => '0',
		10913 => '0',
		10914 => '0',
		10915 => '1',
		10916 => '1',
		10917 => '1',
		10918 => '0',
		10919 => '0',
		10920 => '0',
		10921 => '0',
		10922 => '0',
		10923 => '1',
		10924 => '1',
		10925 => '1',
		10926 => '0',
		10927 => '1',
		10928 => '1',
		10929 => '1',
		10930 => '0',
		10931 => '0',
		10932 => '0',
		10933 => '0',
		10934 => '0',
		10935 => '1',
		10936 => '1',
		10937 => '1',
		10938 => '0',
		10939 => '0',
		10940 => '0',
		10941 => '0',
		10942 => '0',
		10943 => '0',
		10944 => '0',
		10945 => '1',
		10946 => '1',
		10947 => '1',
		10948 => '0',
		10949 => '0',
		10950 => '1',
		10951 => '1',
		10952 => '1',
		10953 => '0',
		10954 => '0',
		10955 => '1',
		10956 => '1',
		10957 => '1',
		10958 => '0',
		10959 => '0',
		10960 => '1',
		10961 => '1',
		10962 => '1',
		10963 => '0',
		10964 => '0',
		10965 => '1',
		10966 => '1',
		10967 => '1',
		10968 => '0',
		10969 => '0',
		10970 => '1',
		10971 => '1',
		10972 => '1',
		10973 => '0',
		10974 => '0',
		10975 => '1',
		10976 => '1',
		10977 => '1',
		10978 => '0',
		10979 => '0',
		10980 => '0',
		10981 => '0',
		10982 => '0',
		10983 => '0',
		10984 => '0',
		10985 => '1',
		10986 => '1',
		10987 => '1',
		10988 => '0',
		10989 => '0',
		10990 => '1',
		10991 => '1',
		10992 => '1',
		10993 => '0',
		10994 => '0',
		10995 => '1',
		10996 => '1',
		10997 => '1',
		10998 => '0',
		10999 => '0',
		11008 => '1',
		11009 => '1',
		11010 => '1',
		11011 => '1',
		11012 => '1',
		11013 => '0',
		11014 => '0',
		11015 => '0',
		11016 => '1',
		11017 => '1',
		11018 => '1',
		11019 => '1',
		11020 => '1',
		11021 => '0',
		11022 => '0',
		11023 => '1',
		11024 => '1',
		11025 => '1',
		11026 => '0',
		11027 => '0',
		11028 => '1',
		11029 => '1',
		11030 => '1',
		11031 => '0',
		11032 => '0',
		11033 => '1',
		11034 => '1',
		11035 => '1',
		11036 => '0',
		11037 => '0',
		11038 => '0',
		11039 => '0',
		11040 => '0',
		11041 => '0',
		11042 => '0',
		11043 => '1',
		11044 => '1',
		11045 => '1',
		11046 => '0',
		11047 => '0',
		11048 => '0',
		11049 => '0',
		11050 => '0',
		11051 => '1',
		11052 => '1',
		11053 => '1',
		11054 => '0',
		11055 => '1',
		11056 => '1',
		11057 => '1',
		11058 => '0',
		11059 => '0',
		11060 => '0',
		11061 => '0',
		11062 => '0',
		11063 => '1',
		11064 => '1',
		11065 => '1',
		11066 => '0',
		11067 => '0',
		11068 => '0',
		11069 => '0',
		11070 => '0',
		11071 => '0',
		11072 => '0',
		11073 => '1',
		11074 => '1',
		11075 => '1',
		11076 => '0',
		11077 => '0',
		11078 => '1',
		11079 => '1',
		11080 => '1',
		11081 => '0',
		11082 => '0',
		11083 => '1',
		11084 => '1',
		11085 => '1',
		11086 => '0',
		11087 => '0',
		11088 => '1',
		11089 => '1',
		11090 => '1',
		11091 => '0',
		11092 => '0',
		11093 => '1',
		11094 => '1',
		11095 => '1',
		11096 => '0',
		11097 => '0',
		11098 => '1',
		11099 => '1',
		11100 => '1',
		11101 => '0',
		11102 => '0',
		11103 => '1',
		11104 => '1',
		11105 => '1',
		11106 => '0',
		11107 => '0',
		11108 => '0',
		11109 => '0',
		11110 => '0',
		11111 => '0',
		11112 => '0',
		11113 => '1',
		11114 => '1',
		11115 => '1',
		11116 => '0',
		11117 => '0',
		11118 => '1',
		11119 => '1',
		11120 => '1',
		11121 => '0',
		11122 => '0',
		11123 => '1',
		11124 => '1',
		11125 => '1',
		11126 => '0',
		11127 => '0',
		11136 => '0',
		11137 => '0',
		11138 => '0',
		11139 => '1',
		11140 => '1',
		11141 => '1',
		11142 => '1',
		11143 => '1',
		11144 => '1',
		11145 => '1',
		11146 => '0',
		11147 => '0',
		11148 => '0',
		11149 => '0',
		11150 => '0',
		11151 => '1',
		11152 => '1',
		11153 => '1',
		11154 => '1',
		11155 => '1',
		11156 => '1',
		11157 => '1',
		11158 => '1',
		11159 => '0',
		11160 => '0',
		11161 => '1',
		11162 => '1',
		11163 => '1',
		11164 => '1',
		11165 => '1',
		11166 => '1',
		11167 => '1',
		11168 => '1',
		11169 => '1',
		11170 => '1',
		11171 => '1',
		11172 => '1',
		11173 => '1',
		11174 => '0',
		11175 => '0',
		11176 => '0',
		11177 => '0',
		11178 => '0',
		11179 => '1',
		11180 => '1',
		11181 => '1',
		11182 => '1',
		11183 => '1',
		11184 => '1',
		11185 => '1',
		11186 => '0',
		11187 => '0',
		11188 => '0',
		11189 => '0',
		11190 => '0',
		11191 => '1',
		11192 => '1',
		11193 => '1',
		11194 => '1',
		11195 => '1',
		11196 => '1',
		11197 => '1',
		11198 => '1',
		11199 => '1',
		11200 => '1',
		11201 => '1',
		11202 => '1',
		11203 => '1',
		11204 => '0',
		11205 => '0',
		11206 => '1',
		11207 => '1',
		11208 => '1',
		11209 => '1',
		11210 => '1',
		11211 => '1',
		11212 => '1',
		11213 => '1',
		11214 => '0',
		11215 => '0',
		11216 => '1',
		11217 => '1',
		11218 => '1',
		11219 => '1',
		11220 => '1',
		11221 => '1',
		11222 => '1',
		11223 => '1',
		11224 => '1',
		11225 => '1',
		11226 => '1',
		11227 => '1',
		11228 => '1',
		11229 => '0',
		11230 => '0',
		11231 => '1',
		11232 => '1',
		11233 => '1',
		11234 => '1',
		11235 => '1',
		11236 => '1',
		11237 => '1',
		11238 => '1',
		11239 => '1',
		11240 => '1',
		11241 => '1',
		11242 => '1',
		11243 => '1',
		11244 => '0',
		11245 => '0',
		11246 => '1',
		11247 => '1',
		11248 => '1',
		11249 => '1',
		11250 => '1',
		11251 => '1',
		11252 => '1',
		11253 => '1',
		11254 => '0',
		11255 => '0',
		11264 => '0',
		11265 => '0',
		11266 => '0',
		11267 => '1',
		11268 => '1',
		11269 => '1',
		11270 => '1',
		11271 => '1',
		11272 => '1',
		11273 => '1',
		11274 => '0',
		11275 => '0',
		11276 => '0',
		11277 => '0',
		11278 => '0',
		11279 => '1',
		11280 => '1',
		11281 => '1',
		11282 => '1',
		11283 => '1',
		11284 => '1',
		11285 => '1',
		11286 => '1',
		11287 => '0',
		11288 => '0',
		11289 => '1',
		11290 => '1',
		11291 => '1',
		11292 => '1',
		11293 => '1',
		11294 => '1',
		11295 => '1',
		11296 => '1',
		11297 => '1',
		11298 => '1',
		11299 => '1',
		11300 => '1',
		11301 => '1',
		11302 => '0',
		11303 => '0',
		11304 => '0',
		11305 => '0',
		11306 => '0',
		11307 => '1',
		11308 => '1',
		11309 => '1',
		11310 => '1',
		11311 => '1',
		11312 => '1',
		11313 => '1',
		11314 => '0',
		11315 => '0',
		11316 => '0',
		11317 => '0',
		11318 => '0',
		11319 => '1',
		11320 => '1',
		11321 => '1',
		11322 => '1',
		11323 => '1',
		11324 => '1',
		11325 => '1',
		11326 => '1',
		11327 => '1',
		11328 => '1',
		11329 => '1',
		11330 => '1',
		11331 => '1',
		11332 => '0',
		11333 => '0',
		11334 => '1',
		11335 => '1',
		11336 => '1',
		11337 => '1',
		11338 => '1',
		11339 => '1',
		11340 => '1',
		11341 => '1',
		11342 => '0',
		11343 => '0',
		11344 => '1',
		11345 => '1',
		11346 => '1',
		11347 => '1',
		11348 => '1',
		11349 => '1',
		11350 => '1',
		11351 => '1',
		11352 => '1',
		11353 => '1',
		11354 => '1',
		11355 => '1',
		11356 => '1',
		11357 => '0',
		11358 => '0',
		11359 => '1',
		11360 => '1',
		11361 => '1',
		11362 => '1',
		11363 => '1',
		11364 => '1',
		11365 => '1',
		11366 => '1',
		11367 => '1',
		11368 => '1',
		11369 => '1',
		11370 => '1',
		11371 => '1',
		11372 => '0',
		11373 => '0',
		11374 => '1',
		11375 => '1',
		11376 => '1',
		11377 => '1',
		11378 => '1',
		11379 => '1',
		11380 => '1',
		11381 => '1',
		11382 => '0',
		11383 => '0',
		11392 => '0',
		11393 => '0',
		11394 => '0',
		11395 => '1',
		11396 => '1',
		11397 => '1',
		11398 => '1',
		11399 => '1',
		11400 => '1',
		11401 => '1',
		11402 => '0',
		11403 => '0',
		11404 => '0',
		11405 => '0',
		11406 => '0',
		11407 => '1',
		11408 => '1',
		11409 => '1',
		11410 => '1',
		11411 => '1',
		11412 => '1',
		11413 => '1',
		11414 => '1',
		11415 => '0',
		11416 => '0',
		11417 => '1',
		11418 => '1',
		11419 => '1',
		11420 => '1',
		11421 => '1',
		11422 => '1',
		11423 => '1',
		11424 => '1',
		11425 => '1',
		11426 => '1',
		11427 => '1',
		11428 => '1',
		11429 => '1',
		11430 => '0',
		11431 => '0',
		11432 => '0',
		11433 => '0',
		11434 => '0',
		11435 => '1',
		11436 => '1',
		11437 => '1',
		11438 => '1',
		11439 => '1',
		11440 => '1',
		11441 => '1',
		11442 => '0',
		11443 => '0',
		11444 => '0',
		11445 => '0',
		11446 => '0',
		11447 => '1',
		11448 => '1',
		11449 => '1',
		11450 => '1',
		11451 => '1',
		11452 => '1',
		11453 => '1',
		11454 => '1',
		11455 => '1',
		11456 => '1',
		11457 => '1',
		11458 => '1',
		11459 => '1',
		11460 => '0',
		11461 => '0',
		11462 => '1',
		11463 => '1',
		11464 => '1',
		11465 => '1',
		11466 => '1',
		11467 => '1',
		11468 => '1',
		11469 => '1',
		11470 => '0',
		11471 => '0',
		11472 => '1',
		11473 => '1',
		11474 => '1',
		11475 => '1',
		11476 => '1',
		11477 => '1',
		11478 => '1',
		11479 => '1',
		11480 => '1',
		11481 => '1',
		11482 => '1',
		11483 => '1',
		11484 => '1',
		11485 => '0',
		11486 => '0',
		11487 => '1',
		11488 => '1',
		11489 => '1',
		11490 => '1',
		11491 => '1',
		11492 => '1',
		11493 => '1',
		11494 => '1',
		11495 => '1',
		11496 => '1',
		11497 => '1',
		11498 => '1',
		11499 => '1',
		11500 => '0',
		11501 => '0',
		11502 => '1',
		11503 => '1',
		11504 => '1',
		11505 => '1',
		11506 => '1',
		11507 => '1',
		11508 => '1',
		11509 => '1',
		11510 => '0',
		11511 => '0',
		11520 => '0',
		11521 => '0',
		11522 => '0',
		11523 => '0',
		11524 => '0',
		11525 => '0',
		11526 => '0',
		11527 => '0',
		11528 => '0',
		11529 => '0',
		11530 => '0',
		11531 => '0',
		11532 => '0',
		11533 => '0',
		11534 => '0',
		11535 => '0',
		11536 => '0',
		11537 => '0',
		11538 => '0',
		11539 => '0',
		11540 => '0',
		11541 => '0',
		11542 => '0',
		11543 => '0',
		11544 => '0',
		11545 => '0',
		11546 => '0',
		11547 => '0',
		11548 => '0',
		11549 => '0',
		11550 => '0',
		11551 => '0',
		11552 => '0',
		11553 => '0',
		11554 => '0',
		11555 => '0',
		11556 => '0',
		11557 => '0',
		11558 => '0',
		11559 => '0',
		11560 => '0',
		11561 => '0',
		11562 => '0',
		11563 => '0',
		11564 => '0',
		11565 => '0',
		11566 => '0',
		11567 => '0',
		11568 => '0',
		11569 => '0',
		11570 => '0',
		11571 => '0',
		11572 => '0',
		11573 => '0',
		11574 => '0',
		11575 => '0',
		11576 => '0',
		11577 => '0',
		11578 => '0',
		11579 => '0',
		11580 => '0',
		11581 => '0',
		11582 => '0',
		11583 => '0',
		11584 => '0',
		11585 => '0',
		11586 => '0',
		11587 => '0',
		11588 => '0',
		11589 => '0',
		11590 => '0',
		11591 => '0',
		11592 => '0',
		11593 => '0',
		11594 => '0',
		11595 => '0',
		11596 => '0',
		11597 => '0',
		11598 => '0',
		11599 => '0',
		11600 => '0',
		11601 => '0',
		11602 => '0',
		11603 => '0',
		11604 => '0',
		11605 => '0',
		11606 => '0',
		11607 => '0',
		11608 => '0',
		11609 => '0',
		11610 => '0',
		11611 => '0',
		11612 => '0',
		11613 => '0',
		11614 => '0',
		11615 => '0',
		11616 => '0',
		11617 => '0',
		11618 => '0',
		11619 => '0',
		11620 => '0',
		11621 => '0',
		11622 => '0',
		11623 => '0',
		11624 => '0',
		11625 => '0',
		11626 => '0',
		11627 => '0',
		11628 => '0',
		11629 => '0',
		11630 => '0',
		11631 => '0',
		11632 => '0',
		11633 => '0',
		11634 => '0',
		11635 => '0',
		11636 => '0',
		11637 => '0',
		11638 => '0',
		11639 => '0',
		11648 => '0',
		11649 => '0',
		11650 => '0',
		11651 => '0',
		11652 => '0',
		11653 => '0',
		11654 => '0',
		11655 => '0',
		11656 => '0',
		11657 => '0',
		11658 => '0',
		11659 => '0',
		11660 => '0',
		11661 => '0',
		11662 => '0',
		11663 => '0',
		11664 => '0',
		11665 => '0',
		11666 => '0',
		11667 => '0',
		11668 => '0',
		11669 => '0',
		11670 => '0',
		11671 => '0',
		11672 => '0',
		11673 => '0',
		11674 => '0',
		11675 => '0',
		11676 => '0',
		11677 => '0',
		11678 => '0',
		11679 => '0',
		11680 => '0',
		11681 => '0',
		11682 => '0',
		11683 => '0',
		11684 => '0',
		11685 => '0',
		11686 => '0',
		11687 => '0',
		11688 => '0',
		11689 => '0',
		11690 => '0',
		11691 => '0',
		11692 => '0',
		11693 => '0',
		11694 => '0',
		11695 => '0',
		11696 => '0',
		11697 => '0',
		11698 => '0',
		11699 => '0',
		11700 => '0',
		11701 => '0',
		11702 => '0',
		11703 => '0',
		11704 => '0',
		11705 => '0',
		11706 => '0',
		11707 => '0',
		11708 => '0',
		11709 => '0',
		11710 => '0',
		11711 => '0',
		11712 => '0',
		11713 => '0',
		11714 => '0',
		11715 => '0',
		11716 => '0',
		11717 => '0',
		11718 => '0',
		11719 => '0',
		11720 => '0',
		11721 => '0',
		11722 => '0',
		11723 => '0',
		11724 => '0',
		11725 => '0',
		11726 => '0',
		11727 => '0',
		11728 => '0',
		11729 => '0',
		11730 => '0',
		11731 => '0',
		11732 => '0',
		11733 => '0',
		11734 => '0',
		11735 => '0',
		11736 => '0',
		11737 => '0',
		11738 => '0',
		11739 => '0',
		11740 => '0',
		11741 => '0',
		11742 => '0',
		11743 => '0',
		11744 => '0',
		11745 => '0',
		11746 => '0',
		11747 => '0',
		11748 => '0',
		11749 => '0',
		11750 => '0',
		11751 => '0',
		11752 => '0',
		11753 => '0',
		11754 => '0',
		11755 => '0',
		11756 => '0',
		11757 => '0',
		11758 => '0',
		11759 => '0',
		11760 => '0',
		11761 => '0',
		11762 => '0',
		11763 => '0',
		11764 => '0',
		11765 => '0',
		11766 => '0',
		11767 => '0',
		11776 => '0',
		11777 => '0',
		11778 => '0',
		11779 => '0',
		11780 => '0',
		11781 => '0',
		11782 => '0',
		11783 => '0',
		11784 => '0',
		11785 => '0',
		11786 => '0',
		11787 => '0',
		11788 => '0',
		11789 => '0',
		11790 => '0',
		11791 => '0',
		11792 => '0',
		11793 => '0',
		11794 => '0',
		11795 => '0',
		11796 => '0',
		11797 => '0',
		11798 => '0',
		11799 => '0',
		11800 => '0',
		11801 => '0',
		11802 => '0',
		11803 => '0',
		11804 => '0',
		11805 => '0',
		11806 => '0',
		11807 => '0',
		11808 => '0',
		11809 => '0',
		11810 => '0',
		11811 => '0',
		11812 => '0',
		11813 => '0',
		11814 => '0',
		11815 => '0',
		11816 => '0',
		11817 => '0',
		11818 => '0',
		11819 => '0',
		11820 => '0',
		11821 => '0',
		11822 => '0',
		11823 => '0',
		11824 => '0',
		11825 => '0',
		11826 => '0',
		11827 => '0',
		11828 => '0',
		11829 => '0',
		11830 => '0',
		11831 => '0',
		11832 => '0',
		11833 => '0',
		11834 => '0',
		11835 => '0',
		11836 => '0',
		11837 => '0',
		11838 => '0',
		11839 => '0',
		11840 => '0',
		11841 => '0',
		11842 => '0',
		11843 => '0',
		11844 => '0',
		11845 => '0',
		11846 => '0',
		11847 => '0',
		11848 => '0',
		11849 => '0',
		11850 => '0',
		11851 => '0',
		11852 => '0',
		11853 => '0',
		11854 => '0',
		11855 => '0',
		11856 => '0',
		11857 => '0',
		11858 => '0',
		11859 => '0',
		11860 => '0',
		11861 => '0',
		11862 => '0',
		11863 => '0',
		11864 => '0',
		11865 => '0',
		11866 => '0',
		11867 => '0',
		11868 => '0',
		11869 => '0',
		11870 => '0',
		11871 => '0',
		11872 => '0',
		11873 => '0',
		11874 => '0',
		11875 => '0',
		11876 => '0',
		11877 => '0',
		11878 => '0',
		11879 => '0',
		11880 => '0',
		11881 => '0',
		11882 => '0',
		11883 => '0',
		11884 => '0',
		11885 => '0',
		11886 => '0',
		11887 => '0',
		11888 => '0',
		11889 => '0',
		11890 => '0',
		11891 => '0',
		11892 => '0',
		11893 => '0',
		11894 => '0',
		11895 => '0',
		11904 => '0',
		11905 => '0',
		11906 => '0',
		11907 => '0',
		11908 => '0',
		11909 => '0',
		11910 => '0',
		11911 => '0',
		11912 => '0',
		11913 => '0',
		11914 => '0',
		11915 => '0',
		11916 => '0',
		11917 => '0',
		11918 => '0',
		11919 => '0',
		11920 => '0',
		11921 => '0',
		11922 => '0',
		11923 => '0',
		11924 => '0',
		11925 => '0',
		11926 => '0',
		11927 => '0',
		11928 => '0',
		11929 => '0',
		11930 => '0',
		11931 => '0',
		11932 => '0',
		11933 => '0',
		11934 => '0',
		11935 => '0',
		11936 => '0',
		11937 => '0',
		11938 => '0',
		11939 => '0',
		11940 => '0',
		11941 => '0',
		11942 => '0',
		11943 => '0',
		11944 => '0',
		11945 => '0',
		11946 => '0',
		11947 => '0',
		11948 => '0',
		11949 => '0',
		11950 => '0',
		11951 => '0',
		11952 => '0',
		11953 => '0',
		11954 => '0',
		11955 => '0',
		11956 => '0',
		11957 => '0',
		11958 => '0',
		11959 => '0',
		11960 => '0',
		11961 => '0',
		11962 => '0',
		11963 => '0',
		11964 => '0',
		11965 => '0',
		11966 => '0',
		11967 => '0',
		11968 => '0',
		11969 => '0',
		11970 => '0',
		11971 => '0',
		11972 => '0',
		11973 => '0',
		11974 => '0',
		11975 => '0',
		11976 => '0',
		11977 => '0',
		11978 => '0',
		11979 => '0',
		11980 => '0',
		11981 => '0',
		11982 => '0',
		11983 => '0',
		11984 => '0',
		11985 => '0',
		11986 => '0',
		11987 => '0',
		11988 => '0',
		11989 => '0',
		11990 => '0',
		11991 => '0',
		11992 => '0',
		11993 => '0',
		11994 => '0',
		11995 => '0',
		11996 => '0',
		11997 => '0',
		11998 => '0',
		11999 => '0',
		12000 => '0',
		12001 => '0',
		12002 => '0',
		12003 => '0',
		12004 => '0',
		12005 => '0',
		12006 => '0',
		12007 => '0',
		12008 => '0',
		12009 => '0',
		12010 => '0',
		12011 => '0',
		12012 => '0',
		12013 => '0',
		12014 => '0',
		12015 => '0',
		12016 => '0',
		12017 => '0',
		12018 => '0',
		12019 => '0',
		12020 => '0',
		12021 => '0',
		12022 => '0',
		12023 => '0',
		12032 => '0',
		12033 => '0',
		12034 => '0',
		12035 => '0',
		12036 => '0',
		12037 => '0',
		12038 => '0',
		12039 => '0',
		12040 => '0',
		12041 => '0',
		12042 => '0',
		12043 => '0',
		12044 => '0',
		12045 => '0',
		12046 => '0',
		12047 => '0',
		12048 => '0',
		12049 => '0',
		12050 => '0',
		12051 => '0',
		12052 => '0',
		12053 => '0',
		12054 => '0',
		12055 => '0',
		12056 => '0',
		12057 => '0',
		12058 => '0',
		12059 => '0',
		12060 => '0',
		12061 => '0',
		12062 => '0',
		12063 => '0',
		12064 => '0',
		12065 => '0',
		12066 => '0',
		12067 => '0',
		12068 => '0',
		12069 => '0',
		12070 => '0',
		12071 => '0',
		12072 => '0',
		12073 => '0',
		12074 => '0',
		12075 => '0',
		12076 => '0',
		12077 => '0',
		12078 => '0',
		12079 => '0',
		12080 => '0',
		12081 => '0',
		12082 => '0',
		12083 => '0',
		12084 => '0',
		12085 => '0',
		12086 => '0',
		12087 => '0',
		12088 => '0',
		12089 => '0',
		12090 => '0',
		12091 => '0',
		12092 => '0',
		12093 => '0',
		12094 => '0',
		12095 => '0',
		12096 => '0',
		12097 => '0',
		12098 => '0',
		12099 => '0',
		12100 => '0',
		12101 => '0',
		12102 => '0',
		12103 => '0',
		12104 => '0',
		12105 => '0',
		12106 => '0',
		12107 => '0',
		12108 => '0',
		12109 => '0',
		12110 => '0',
		12111 => '0',
		12112 => '0',
		12113 => '0',
		12114 => '0',
		12115 => '0',
		12116 => '0',
		12117 => '0',
		12118 => '0',
		12119 => '0',
		12120 => '0',
		12121 => '0',
		12122 => '0',
		12123 => '0',
		12124 => '0',
		12125 => '0',
		12126 => '0',
		12127 => '0',
		12128 => '0',
		12129 => '0',
		12130 => '0',
		12131 => '0',
		12132 => '0',
		12133 => '0',
		12134 => '0',
		12135 => '0',
		12136 => '0',
		12137 => '0',
		12138 => '0',
		12139 => '0',
		12140 => '0',
		12141 => '0',
		12142 => '0',
		12143 => '0',
		12144 => '0',
		12145 => '0',
		12146 => '0',
		12147 => '0',
		12148 => '0',
		12149 => '0',
		12150 => '0',
		12151 => '0',
		12160 => '0',
		12161 => '0',
		12162 => '0',
		12163 => '0',
		12164 => '0',
		12165 => '0',
		12166 => '0',
		12167 => '0',
		12168 => '0',
		12169 => '0',
		12170 => '0',
		12171 => '0',
		12172 => '0',
		12173 => '0',
		12174 => '0',
		12175 => '0',
		12176 => '0',
		12177 => '0',
		12178 => '0',
		12179 => '0',
		12180 => '0',
		12181 => '0',
		12182 => '0',
		12183 => '0',
		12184 => '0',
		12185 => '0',
		12186 => '0',
		12187 => '0',
		12188 => '0',
		12189 => '0',
		12190 => '0',
		12191 => '0',
		12192 => '0',
		12193 => '0',
		12194 => '0',
		12195 => '0',
		12196 => '0',
		12197 => '0',
		12198 => '0',
		12199 => '0',
		12200 => '0',
		12201 => '0',
		12202 => '0',
		12203 => '0',
		12204 => '0',
		12205 => '0',
		12206 => '0',
		12207 => '0',
		12208 => '0',
		12209 => '0',
		12210 => '0',
		12211 => '0',
		12212 => '0',
		12213 => '0',
		12214 => '0',
		12215 => '0',
		12216 => '0',
		12217 => '0',
		12218 => '0',
		12219 => '0',
		12220 => '0',
		12221 => '0',
		12222 => '0',
		12223 => '0',
		12224 => '0',
		12225 => '0',
		12226 => '0',
		12227 => '0',
		12228 => '0',
		12229 => '0',
		12230 => '0',
		12231 => '0',
		12232 => '0',
		12233 => '0',
		12234 => '0',
		12235 => '0',
		12236 => '0',
		12237 => '0',
		12238 => '0',
		12239 => '0',
		12240 => '0',
		12241 => '0',
		12242 => '0',
		12243 => '0',
		12244 => '0',
		12245 => '0',
		12246 => '0',
		12247 => '0',
		12248 => '0',
		12249 => '0',
		12250 => '0',
		12251 => '0',
		12252 => '0',
		12253 => '0',
		12254 => '0',
		12255 => '0',
		12256 => '0',
		12257 => '0',
		12258 => '0',
		12259 => '0',
		12260 => '0',
		12261 => '0',
		12262 => '0',
		12263 => '0',
		12264 => '0',
		12265 => '0',
		12266 => '0',
		12267 => '0',
		12268 => '0',
		12269 => '0',
		12270 => '0',
		12271 => '0',
		12272 => '0',
		12273 => '0',
		12274 => '0',
		12275 => '0',
		12276 => '0',
		12277 => '0',
		12278 => '0',
		12279 => '0',
		12288 => '1',
		12289 => '1',
		12290 => '1',
		12291 => '1',
		12292 => '1',
		12293 => '1',
		12294 => '1',
		12295 => '1',
		12296 => '1',
		12297 => '1',
		12298 => '1',
		12299 => '1',
		12300 => '1',
		12301 => '0',
		12302 => '0',
		12303 => '1',
		12304 => '1',
		12305 => '1',
		12306 => '1',
		12307 => '1',
		12308 => '1',
		12309 => '1',
		12310 => '1',
		12311 => '0',
		12312 => '0',
		12313 => '1',
		12314 => '1',
		12315 => '1',
		12316 => '1',
		12317 => '1',
		12318 => '1',
		12319 => '1',
		12320 => '1',
		12321 => '1',
		12322 => '1',
		12323 => '1',
		12324 => '1',
		12325 => '1',
		12326 => '0',
		12327 => '0',
		12328 => '1',
		12329 => '1',
		12330 => '1',
		12331 => '1',
		12332 => '1',
		12333 => '1',
		12334 => '1',
		12335 => '1',
		12336 => '1',
		12337 => '1',
		12338 => '1',
		12339 => '1',
		12340 => '1',
		12341 => '0',
		12342 => '0',
		12343 => '1',
		12344 => '1',
		12345 => '1',
		12346 => '1',
		12347 => '1',
		12348 => '1',
		12349 => '1',
		12350 => '1',
		12351 => '1',
		12352 => '1',
		12353 => '1',
		12354 => '1',
		12355 => '1',
		12356 => '0',
		12357 => '0',
		12358 => '1',
		12359 => '1',
		12360 => '1',
		12361 => '1',
		12362 => '1',
		12363 => '1',
		12364 => '1',
		12365 => '1',
		12366 => '0',
		12367 => '0',
		12368 => '1',
		12369 => '1',
		12370 => '1',
		12371 => '1',
		12372 => '1',
		12373 => '1',
		12374 => '1',
		12375 => '1',
		12376 => '1',
		12377 => '1',
		12378 => '1',
		12379 => '1',
		12380 => '1',
		12381 => '0',
		12382 => '0',
		12383 => '1',
		12384 => '1',
		12385 => '1',
		12386 => '1',
		12387 => '1',
		12388 => '1',
		12389 => '1',
		12390 => '1',
		12391 => '1',
		12392 => '1',
		12393 => '1',
		12394 => '1',
		12395 => '1',
		12396 => '0',
		12397 => '0',
		12398 => '1',
		12399 => '1',
		12400 => '1',
		12401 => '1',
		12402 => '1',
		12403 => '1',
		12404 => '1',
		12405 => '1',
		12406 => '0',
		12407 => '0',
		12416 => '1',
		12417 => '1',
		12418 => '1',
		12419 => '1',
		12420 => '1',
		12421 => '1',
		12422 => '1',
		12423 => '1',
		12424 => '1',
		12425 => '1',
		12426 => '1',
		12427 => '1',
		12428 => '1',
		12429 => '0',
		12430 => '0',
		12431 => '1',
		12432 => '1',
		12433 => '1',
		12434 => '1',
		12435 => '1',
		12436 => '1',
		12437 => '1',
		12438 => '1',
		12439 => '0',
		12440 => '0',
		12441 => '1',
		12442 => '1',
		12443 => '1',
		12444 => '1',
		12445 => '1',
		12446 => '1',
		12447 => '1',
		12448 => '1',
		12449 => '1',
		12450 => '1',
		12451 => '1',
		12452 => '1',
		12453 => '1',
		12454 => '0',
		12455 => '0',
		12456 => '1',
		12457 => '1',
		12458 => '1',
		12459 => '1',
		12460 => '1',
		12461 => '1',
		12462 => '1',
		12463 => '1',
		12464 => '1',
		12465 => '1',
		12466 => '1',
		12467 => '1',
		12468 => '1',
		12469 => '0',
		12470 => '0',
		12471 => '1',
		12472 => '1',
		12473 => '1',
		12474 => '1',
		12475 => '1',
		12476 => '1',
		12477 => '1',
		12478 => '1',
		12479 => '1',
		12480 => '1',
		12481 => '1',
		12482 => '1',
		12483 => '1',
		12484 => '0',
		12485 => '0',
		12486 => '1',
		12487 => '1',
		12488 => '1',
		12489 => '1',
		12490 => '1',
		12491 => '1',
		12492 => '1',
		12493 => '1',
		12494 => '0',
		12495 => '0',
		12496 => '1',
		12497 => '1',
		12498 => '1',
		12499 => '1',
		12500 => '1',
		12501 => '1',
		12502 => '1',
		12503 => '1',
		12504 => '1',
		12505 => '1',
		12506 => '1',
		12507 => '1',
		12508 => '1',
		12509 => '0',
		12510 => '0',
		12511 => '1',
		12512 => '1',
		12513 => '1',
		12514 => '1',
		12515 => '1',
		12516 => '1',
		12517 => '1',
		12518 => '1',
		12519 => '1',
		12520 => '1',
		12521 => '1',
		12522 => '1',
		12523 => '1',
		12524 => '0',
		12525 => '0',
		12526 => '1',
		12527 => '1',
		12528 => '1',
		12529 => '1',
		12530 => '1',
		12531 => '1',
		12532 => '1',
		12533 => '1',
		12534 => '0',
		12535 => '0',
		12544 => '1',
		12545 => '1',
		12546 => '1',
		12547 => '1',
		12548 => '1',
		12549 => '1',
		12550 => '1',
		12551 => '1',
		12552 => '1',
		12553 => '1',
		12554 => '1',
		12555 => '1',
		12556 => '1',
		12557 => '0',
		12558 => '0',
		12559 => '1',
		12560 => '1',
		12561 => '1',
		12562 => '1',
		12563 => '1',
		12564 => '1',
		12565 => '1',
		12566 => '1',
		12567 => '0',
		12568 => '0',
		12569 => '1',
		12570 => '1',
		12571 => '1',
		12572 => '1',
		12573 => '1',
		12574 => '1',
		12575 => '1',
		12576 => '1',
		12577 => '1',
		12578 => '1',
		12579 => '1',
		12580 => '1',
		12581 => '1',
		12582 => '0',
		12583 => '0',
		12584 => '1',
		12585 => '1',
		12586 => '1',
		12587 => '1',
		12588 => '1',
		12589 => '1',
		12590 => '1',
		12591 => '1',
		12592 => '1',
		12593 => '1',
		12594 => '1',
		12595 => '1',
		12596 => '1',
		12597 => '0',
		12598 => '0',
		12599 => '1',
		12600 => '1',
		12601 => '1',
		12602 => '1',
		12603 => '1',
		12604 => '1',
		12605 => '1',
		12606 => '1',
		12607 => '1',
		12608 => '1',
		12609 => '1',
		12610 => '1',
		12611 => '1',
		12612 => '0',
		12613 => '0',
		12614 => '1',
		12615 => '1',
		12616 => '1',
		12617 => '1',
		12618 => '1',
		12619 => '1',
		12620 => '1',
		12621 => '1',
		12622 => '0',
		12623 => '0',
		12624 => '1',
		12625 => '1',
		12626 => '1',
		12627 => '1',
		12628 => '1',
		12629 => '1',
		12630 => '1',
		12631 => '1',
		12632 => '1',
		12633 => '1',
		12634 => '1',
		12635 => '1',
		12636 => '1',
		12637 => '0',
		12638 => '0',
		12639 => '1',
		12640 => '1',
		12641 => '1',
		12642 => '1',
		12643 => '1',
		12644 => '1',
		12645 => '1',
		12646 => '1',
		12647 => '1',
		12648 => '1',
		12649 => '1',
		12650 => '1',
		12651 => '1',
		12652 => '0',
		12653 => '0',
		12654 => '1',
		12655 => '1',
		12656 => '1',
		12657 => '1',
		12658 => '1',
		12659 => '1',
		12660 => '1',
		12661 => '1',
		12662 => '0',
		12663 => '0',
		12672 => '1',
		12673 => '1',
		12674 => '1',
		12675 => '0',
		12676 => '0',
		12677 => '1',
		12678 => '1',
		12679 => '1',
		12680 => '0',
		12681 => '0',
		12682 => '1',
		12683 => '1',
		12684 => '1',
		12685 => '0',
		12686 => '0',
		12687 => '1',
		12688 => '1',
		12689 => '1',
		12690 => '0',
		12691 => '0',
		12692 => '1',
		12693 => '1',
		12694 => '1',
		12695 => '0',
		12696 => '0',
		12697 => '1',
		12698 => '1',
		12699 => '1',
		12700 => '0',
		12701 => '0',
		12702 => '0',
		12703 => '0',
		12704 => '0',
		12705 => '0',
		12706 => '0',
		12707 => '1',
		12708 => '1',
		12709 => '1',
		12710 => '0',
		12711 => '0',
		12712 => '1',
		12713 => '1',
		12714 => '1',
		12715 => '0',
		12716 => '0',
		12717 => '0',
		12718 => '0',
		12719 => '0',
		12720 => '0',
		12721 => '0',
		12722 => '1',
		12723 => '1',
		12724 => '1',
		12725 => '0',
		12726 => '0',
		12727 => '1',
		12728 => '1',
		12729 => '1',
		12730 => '0',
		12731 => '0',
		12732 => '0',
		12733 => '0',
		12734 => '0',
		12735 => '0',
		12736 => '0',
		12737 => '1',
		12738 => '1',
		12739 => '1',
		12740 => '0',
		12741 => '0',
		12742 => '1',
		12743 => '1',
		12744 => '1',
		12745 => '0',
		12746 => '0',
		12747 => '1',
		12748 => '1',
		12749 => '1',
		12750 => '0',
		12751 => '0',
		12752 => '1',
		12753 => '1',
		12754 => '1',
		12755 => '0',
		12756 => '0',
		12757 => '0',
		12758 => '0',
		12759 => '0',
		12760 => '0',
		12761 => '0',
		12762 => '1',
		12763 => '1',
		12764 => '1',
		12765 => '0',
		12766 => '0',
		12767 => '1',
		12768 => '1',
		12769 => '1',
		12770 => '0',
		12771 => '0',
		12772 => '0',
		12773 => '0',
		12774 => '0',
		12775 => '0',
		12776 => '0',
		12777 => '1',
		12778 => '1',
		12779 => '1',
		12780 => '0',
		12781 => '0',
		12782 => '1',
		12783 => '1',
		12784 => '1',
		12785 => '0',
		12786 => '0',
		12787 => '1',
		12788 => '1',
		12789 => '1',
		12790 => '0',
		12791 => '0',
		12800 => '1',
		12801 => '1',
		12802 => '1',
		12803 => '0',
		12804 => '0',
		12805 => '1',
		12806 => '1',
		12807 => '1',
		12808 => '0',
		12809 => '0',
		12810 => '1',
		12811 => '1',
		12812 => '1',
		12813 => '0',
		12814 => '0',
		12815 => '1',
		12816 => '1',
		12817 => '1',
		12818 => '0',
		12819 => '0',
		12820 => '1',
		12821 => '1',
		12822 => '1',
		12823 => '0',
		12824 => '0',
		12825 => '1',
		12826 => '1',
		12827 => '1',
		12828 => '0',
		12829 => '0',
		12830 => '0',
		12831 => '0',
		12832 => '0',
		12833 => '0',
		12834 => '0',
		12835 => '1',
		12836 => '1',
		12837 => '1',
		12838 => '0',
		12839 => '0',
		12840 => '1',
		12841 => '1',
		12842 => '1',
		12843 => '0',
		12844 => '0',
		12845 => '0',
		12846 => '0',
		12847 => '0',
		12848 => '0',
		12849 => '0',
		12850 => '1',
		12851 => '1',
		12852 => '1',
		12853 => '0',
		12854 => '0',
		12855 => '1',
		12856 => '1',
		12857 => '1',
		12858 => '0',
		12859 => '0',
		12860 => '0',
		12861 => '0',
		12862 => '0',
		12863 => '0',
		12864 => '0',
		12865 => '1',
		12866 => '1',
		12867 => '1',
		12868 => '0',
		12869 => '0',
		12870 => '1',
		12871 => '1',
		12872 => '1',
		12873 => '0',
		12874 => '0',
		12875 => '1',
		12876 => '1',
		12877 => '1',
		12878 => '0',
		12879 => '0',
		12880 => '1',
		12881 => '1',
		12882 => '1',
		12883 => '0',
		12884 => '0',
		12885 => '0',
		12886 => '0',
		12887 => '0',
		12888 => '0',
		12889 => '0',
		12890 => '1',
		12891 => '1',
		12892 => '1',
		12893 => '0',
		12894 => '0',
		12895 => '1',
		12896 => '1',
		12897 => '1',
		12898 => '0',
		12899 => '0',
		12900 => '0',
		12901 => '0',
		12902 => '0',
		12903 => '0',
		12904 => '0',
		12905 => '1',
		12906 => '1',
		12907 => '1',
		12908 => '0',
		12909 => '0',
		12910 => '1',
		12911 => '1',
		12912 => '1',
		12913 => '0',
		12914 => '0',
		12915 => '1',
		12916 => '1',
		12917 => '1',
		12918 => '0',
		12919 => '0',
		12928 => '1',
		12929 => '1',
		12930 => '1',
		12931 => '0',
		12932 => '0',
		12933 => '1',
		12934 => '1',
		12935 => '1',
		12936 => '0',
		12937 => '0',
		12938 => '1',
		12939 => '1',
		12940 => '1',
		12941 => '0',
		12942 => '0',
		12943 => '1',
		12944 => '1',
		12945 => '1',
		12946 => '0',
		12947 => '0',
		12948 => '1',
		12949 => '1',
		12950 => '1',
		12951 => '0',
		12952 => '0',
		12953 => '1',
		12954 => '1',
		12955 => '1',
		12956 => '0',
		12957 => '0',
		12958 => '0',
		12959 => '0',
		12960 => '0',
		12961 => '0',
		12962 => '0',
		12963 => '1',
		12964 => '1',
		12965 => '1',
		12966 => '0',
		12967 => '0',
		12968 => '1',
		12969 => '1',
		12970 => '1',
		12971 => '1',
		12972 => '1',
		12973 => '1',
		12974 => '0',
		12975 => '1',
		12976 => '1',
		12977 => '1',
		12978 => '1',
		12979 => '1',
		12980 => '1',
		12981 => '0',
		12982 => '0',
		12983 => '1',
		12984 => '1',
		12985 => '1',
		12986 => '0',
		12987 => '0',
		12988 => '0',
		12989 => '0',
		12990 => '0',
		12991 => '0',
		12992 => '0',
		12993 => '1',
		12994 => '1',
		12995 => '1',
		12996 => '0',
		12997 => '0',
		12998 => '1',
		12999 => '1',
		13000 => '1',
		13001 => '0',
		13002 => '0',
		13003 => '1',
		13004 => '1',
		13005 => '1',
		13006 => '0',
		13007 => '0',
		13008 => '1',
		13009 => '1',
		13010 => '1',
		13011 => '0',
		13012 => '0',
		13013 => '1',
		13014 => '1',
		13015 => '1',
		13016 => '0',
		13017 => '0',
		13018 => '1',
		13019 => '1',
		13020 => '1',
		13021 => '0',
		13022 => '0',
		13023 => '1',
		13024 => '1',
		13025 => '1',
		13026 => '0',
		13027 => '0',
		13028 => '1',
		13029 => '1',
		13030 => '1',
		13031 => '1',
		13032 => '1',
		13033 => '1',
		13034 => '1',
		13035 => '1',
		13036 => '0',
		13037 => '0',
		13038 => '1',
		13039 => '1',
		13040 => '1',
		13041 => '0',
		13042 => '0',
		13043 => '1',
		13044 => '1',
		13045 => '1',
		13046 => '0',
		13047 => '0',
		13056 => '1',
		13057 => '1',
		13058 => '1',
		13059 => '0',
		13060 => '0',
		13061 => '1',
		13062 => '1',
		13063 => '1',
		13064 => '0',
		13065 => '0',
		13066 => '1',
		13067 => '1',
		13068 => '1',
		13069 => '0',
		13070 => '0',
		13071 => '1',
		13072 => '1',
		13073 => '1',
		13074 => '0',
		13075 => '0',
		13076 => '1',
		13077 => '1',
		13078 => '1',
		13079 => '0',
		13080 => '0',
		13081 => '1',
		13082 => '1',
		13083 => '1',
		13084 => '0',
		13085 => '0',
		13086 => '1',
		13087 => '1',
		13088 => '1',
		13089 => '0',
		13090 => '0',
		13091 => '1',
		13092 => '1',
		13093 => '1',
		13094 => '0',
		13095 => '0',
		13096 => '1',
		13097 => '1',
		13098 => '1',
		13099 => '1',
		13100 => '1',
		13101 => '1',
		13102 => '0',
		13103 => '1',
		13104 => '1',
		13105 => '1',
		13106 => '1',
		13107 => '1',
		13108 => '1',
		13109 => '0',
		13110 => '0',
		13111 => '1',
		13112 => '1',
		13113 => '1',
		13114 => '0',
		13115 => '0',
		13116 => '1',
		13117 => '1',
		13118 => '1',
		13119 => '0',
		13120 => '0',
		13121 => '1',
		13122 => '1',
		13123 => '1',
		13124 => '0',
		13125 => '0',
		13126 => '1',
		13127 => '1',
		13128 => '1',
		13129 => '0',
		13130 => '0',
		13131 => '1',
		13132 => '1',
		13133 => '1',
		13134 => '0',
		13135 => '0',
		13136 => '1',
		13137 => '1',
		13138 => '1',
		13139 => '0',
		13140 => '0',
		13141 => '1',
		13142 => '1',
		13143 => '1',
		13144 => '0',
		13145 => '0',
		13146 => '1',
		13147 => '1',
		13148 => '1',
		13149 => '0',
		13150 => '0',
		13151 => '1',
		13152 => '1',
		13153 => '1',
		13154 => '0',
		13155 => '0',
		13156 => '1',
		13157 => '1',
		13158 => '1',
		13159 => '1',
		13160 => '1',
		13161 => '1',
		13162 => '1',
		13163 => '1',
		13164 => '0',
		13165 => '0',
		13166 => '1',
		13167 => '1',
		13168 => '1',
		13169 => '0',
		13170 => '0',
		13171 => '1',
		13172 => '1',
		13173 => '1',
		13174 => '0',
		13175 => '0',
		13184 => '1',
		13185 => '1',
		13186 => '1',
		13187 => '0',
		13188 => '0',
		13189 => '1',
		13190 => '1',
		13191 => '1',
		13192 => '0',
		13193 => '0',
		13194 => '1',
		13195 => '1',
		13196 => '1',
		13197 => '0',
		13198 => '0',
		13199 => '1',
		13200 => '1',
		13201 => '1',
		13202 => '0',
		13203 => '0',
		13204 => '1',
		13205 => '1',
		13206 => '1',
		13207 => '0',
		13208 => '0',
		13209 => '1',
		13210 => '1',
		13211 => '1',
		13212 => '0',
		13213 => '0',
		13214 => '1',
		13215 => '1',
		13216 => '1',
		13217 => '0',
		13218 => '0',
		13219 => '1',
		13220 => '1',
		13221 => '1',
		13222 => '0',
		13223 => '0',
		13224 => '1',
		13225 => '1',
		13226 => '1',
		13227 => '1',
		13228 => '1',
		13229 => '1',
		13230 => '0',
		13231 => '1',
		13232 => '1',
		13233 => '1',
		13234 => '1',
		13235 => '1',
		13236 => '1',
		13237 => '0',
		13238 => '0',
		13239 => '1',
		13240 => '1',
		13241 => '1',
		13242 => '0',
		13243 => '0',
		13244 => '1',
		13245 => '1',
		13246 => '1',
		13247 => '0',
		13248 => '0',
		13249 => '1',
		13250 => '1',
		13251 => '1',
		13252 => '0',
		13253 => '0',
		13254 => '1',
		13255 => '1',
		13256 => '1',
		13257 => '0',
		13258 => '0',
		13259 => '1',
		13260 => '1',
		13261 => '1',
		13262 => '0',
		13263 => '0',
		13264 => '1',
		13265 => '1',
		13266 => '1',
		13267 => '0',
		13268 => '0',
		13269 => '1',
		13270 => '1',
		13271 => '1',
		13272 => '0',
		13273 => '0',
		13274 => '1',
		13275 => '1',
		13276 => '1',
		13277 => '0',
		13278 => '0',
		13279 => '1',
		13280 => '1',
		13281 => '1',
		13282 => '0',
		13283 => '0',
		13284 => '1',
		13285 => '1',
		13286 => '1',
		13287 => '1',
		13288 => '1',
		13289 => '1',
		13290 => '1',
		13291 => '1',
		13292 => '0',
		13293 => '0',
		13294 => '1',
		13295 => '1',
		13296 => '1',
		13297 => '0',
		13298 => '0',
		13299 => '1',
		13300 => '1',
		13301 => '1',
		13302 => '0',
		13303 => '0',
		13312 => '1',
		13313 => '1',
		13314 => '1',
		13315 => '0',
		13316 => '0',
		13317 => '1',
		13318 => '1',
		13319 => '1',
		13320 => '0',
		13321 => '0',
		13322 => '1',
		13323 => '1',
		13324 => '1',
		13325 => '0',
		13326 => '0',
		13327 => '1',
		13328 => '1',
		13329 => '1',
		13330 => '0',
		13331 => '0',
		13332 => '1',
		13333 => '1',
		13334 => '1',
		13335 => '0',
		13336 => '0',
		13337 => '1',
		13338 => '1',
		13339 => '1',
		13340 => '0',
		13341 => '0',
		13342 => '1',
		13343 => '1',
		13344 => '1',
		13345 => '1',
		13346 => '1',
		13347 => '1',
		13348 => '1',
		13349 => '1',
		13350 => '0',
		13351 => '0',
		13352 => '0',
		13353 => '0',
		13354 => '0',
		13355 => '1',
		13356 => '1',
		13357 => '1',
		13358 => '0',
		13359 => '1',
		13360 => '1',
		13361 => '1',
		13362 => '0',
		13363 => '0',
		13364 => '0',
		13365 => '0',
		13366 => '0',
		13367 => '1',
		13368 => '1',
		13369 => '1',
		13370 => '0',
		13371 => '0',
		13372 => '1',
		13373 => '1',
		13374 => '1',
		13375 => '0',
		13376 => '0',
		13377 => '1',
		13378 => '1',
		13379 => '1',
		13380 => '0',
		13381 => '0',
		13382 => '1',
		13383 => '1',
		13384 => '1',
		13385 => '0',
		13386 => '0',
		13387 => '1',
		13388 => '1',
		13389 => '1',
		13390 => '0',
		13391 => '0',
		13392 => '1',
		13393 => '1',
		13394 => '1',
		13395 => '0',
		13396 => '0',
		13397 => '0',
		13398 => '0',
		13399 => '0',
		13400 => '1',
		13401 => '1',
		13402 => '1',
		13403 => '1',
		13404 => '1',
		13405 => '0',
		13406 => '0',
		13407 => '1',
		13408 => '1',
		13409 => '1',
		13410 => '0',
		13411 => '0',
		13412 => '0',
		13413 => '0',
		13414 => '0',
		13415 => '0',
		13416 => '0',
		13417 => '1',
		13418 => '1',
		13419 => '1',
		13420 => '0',
		13421 => '0',
		13422 => '1',
		13423 => '1',
		13424 => '1',
		13425 => '0',
		13426 => '0',
		13427 => '1',
		13428 => '1',
		13429 => '1',
		13430 => '0',
		13431 => '0',
		13440 => '1',
		13441 => '1',
		13442 => '1',
		13443 => '0',
		13444 => '0',
		13445 => '1',
		13446 => '1',
		13447 => '1',
		13448 => '0',
		13449 => '0',
		13450 => '1',
		13451 => '1',
		13452 => '1',
		13453 => '0',
		13454 => '0',
		13455 => '1',
		13456 => '1',
		13457 => '1',
		13458 => '0',
		13459 => '0',
		13460 => '1',
		13461 => '1',
		13462 => '1',
		13463 => '0',
		13464 => '0',
		13465 => '1',
		13466 => '1',
		13467 => '1',
		13468 => '0',
		13469 => '0',
		13470 => '1',
		13471 => '1',
		13472 => '1',
		13473 => '1',
		13474 => '1',
		13475 => '1',
		13476 => '1',
		13477 => '1',
		13478 => '0',
		13479 => '0',
		13480 => '0',
		13481 => '0',
		13482 => '0',
		13483 => '1',
		13484 => '1',
		13485 => '1',
		13486 => '0',
		13487 => '1',
		13488 => '1',
		13489 => '1',
		13490 => '0',
		13491 => '0',
		13492 => '0',
		13493 => '0',
		13494 => '0',
		13495 => '1',
		13496 => '1',
		13497 => '1',
		13498 => '0',
		13499 => '0',
		13500 => '1',
		13501 => '1',
		13502 => '1',
		13503 => '0',
		13504 => '0',
		13505 => '1',
		13506 => '1',
		13507 => '1',
		13508 => '0',
		13509 => '0',
		13510 => '1',
		13511 => '1',
		13512 => '1',
		13513 => '0',
		13514 => '0',
		13515 => '1',
		13516 => '1',
		13517 => '1',
		13518 => '0',
		13519 => '0',
		13520 => '1',
		13521 => '1',
		13522 => '1',
		13523 => '0',
		13524 => '0',
		13525 => '0',
		13526 => '0',
		13527 => '0',
		13528 => '1',
		13529 => '1',
		13530 => '1',
		13531 => '1',
		13532 => '1',
		13533 => '0',
		13534 => '0',
		13535 => '1',
		13536 => '1',
		13537 => '1',
		13538 => '0',
		13539 => '0',
		13540 => '0',
		13541 => '0',
		13542 => '0',
		13543 => '0',
		13544 => '0',
		13545 => '1',
		13546 => '1',
		13547 => '1',
		13548 => '0',
		13549 => '0',
		13550 => '1',
		13551 => '1',
		13552 => '1',
		13553 => '0',
		13554 => '0',
		13555 => '1',
		13556 => '1',
		13557 => '1',
		13558 => '0',
		13559 => '0',
		13568 => '1',
		13569 => '1',
		13570 => '1',
		13571 => '0',
		13572 => '0',
		13573 => '1',
		13574 => '1',
		13575 => '1',
		13576 => '0',
		13577 => '0',
		13578 => '1',
		13579 => '1',
		13580 => '1',
		13581 => '0',
		13582 => '0',
		13583 => '1',
		13584 => '1',
		13585 => '1',
		13586 => '0',
		13587 => '0',
		13588 => '1',
		13589 => '1',
		13590 => '1',
		13591 => '0',
		13592 => '0',
		13593 => '1',
		13594 => '1',
		13595 => '1',
		13596 => '0',
		13597 => '0',
		13598 => '1',
		13599 => '1',
		13600 => '1',
		13601 => '1',
		13602 => '1',
		13603 => '1',
		13604 => '1',
		13605 => '1',
		13606 => '0',
		13607 => '0',
		13608 => '0',
		13609 => '0',
		13610 => '0',
		13611 => '1',
		13612 => '1',
		13613 => '1',
		13614 => '0',
		13615 => '1',
		13616 => '1',
		13617 => '1',
		13618 => '0',
		13619 => '0',
		13620 => '0',
		13621 => '0',
		13622 => '0',
		13623 => '1',
		13624 => '1',
		13625 => '1',
		13626 => '0',
		13627 => '0',
		13628 => '1',
		13629 => '1',
		13630 => '1',
		13631 => '0',
		13632 => '0',
		13633 => '1',
		13634 => '1',
		13635 => '1',
		13636 => '0',
		13637 => '0',
		13638 => '1',
		13639 => '1',
		13640 => '1',
		13641 => '0',
		13642 => '0',
		13643 => '1',
		13644 => '1',
		13645 => '1',
		13646 => '0',
		13647 => '0',
		13648 => '1',
		13649 => '1',
		13650 => '1',
		13651 => '0',
		13652 => '0',
		13653 => '1',
		13654 => '1',
		13655 => '1',
		13656 => '1',
		13657 => '1',
		13658 => '1',
		13659 => '1',
		13660 => '1',
		13661 => '0',
		13662 => '0',
		13663 => '1',
		13664 => '1',
		13665 => '1',
		13666 => '0',
		13667 => '0',
		13668 => '1',
		13669 => '1',
		13670 => '1',
		13671 => '1',
		13672 => '1',
		13673 => '1',
		13674 => '1',
		13675 => '1',
		13676 => '0',
		13677 => '0',
		13678 => '1',
		13679 => '1',
		13680 => '1',
		13681 => '1',
		13682 => '1',
		13683 => '1',
		13684 => '1',
		13685 => '1',
		13686 => '0',
		13687 => '0',
		13696 => '1',
		13697 => '1',
		13698 => '1',
		13699 => '0',
		13700 => '0',
		13701 => '1',
		13702 => '1',
		13703 => '1',
		13704 => '0',
		13705 => '0',
		13706 => '1',
		13707 => '1',
		13708 => '1',
		13709 => '0',
		13710 => '0',
		13711 => '1',
		13712 => '1',
		13713 => '1',
		13714 => '0',
		13715 => '0',
		13716 => '1',
		13717 => '1',
		13718 => '1',
		13719 => '0',
		13720 => '0',
		13721 => '1',
		13722 => '1',
		13723 => '1',
		13724 => '0',
		13725 => '0',
		13726 => '1',
		13727 => '1',
		13728 => '1',
		13729 => '0',
		13730 => '0',
		13731 => '1',
		13732 => '1',
		13733 => '1',
		13734 => '0',
		13735 => '0',
		13736 => '0',
		13737 => '0',
		13738 => '0',
		13739 => '1',
		13740 => '1',
		13741 => '1',
		13742 => '0',
		13743 => '1',
		13744 => '1',
		13745 => '1',
		13746 => '0',
		13747 => '0',
		13748 => '0',
		13749 => '0',
		13750 => '0',
		13751 => '1',
		13752 => '1',
		13753 => '1',
		13754 => '0',
		13755 => '0',
		13756 => '1',
		13757 => '1',
		13758 => '1',
		13759 => '0',
		13760 => '0',
		13761 => '1',
		13762 => '1',
		13763 => '1',
		13764 => '0',
		13765 => '0',
		13766 => '1',
		13767 => '1',
		13768 => '1',
		13769 => '0',
		13770 => '0',
		13771 => '1',
		13772 => '1',
		13773 => '1',
		13774 => '0',
		13775 => '0',
		13776 => '1',
		13777 => '1',
		13778 => '1',
		13779 => '0',
		13780 => '0',
		13781 => '1',
		13782 => '1',
		13783 => '1',
		13784 => '0',
		13785 => '0',
		13786 => '1',
		13787 => '1',
		13788 => '1',
		13789 => '0',
		13790 => '0',
		13791 => '1',
		13792 => '1',
		13793 => '1',
		13794 => '0',
		13795 => '0',
		13796 => '1',
		13797 => '1',
		13798 => '1',
		13799 => '1',
		13800 => '1',
		13801 => '1',
		13802 => '1',
		13803 => '1',
		13804 => '0',
		13805 => '0',
		13806 => '1',
		13807 => '1',
		13808 => '1',
		13809 => '1',
		13810 => '1',
		13811 => '1',
		13812 => '1',
		13813 => '1',
		13814 => '0',
		13815 => '0',
		13824 => '1',
		13825 => '1',
		13826 => '1',
		13827 => '0',
		13828 => '0',
		13829 => '1',
		13830 => '1',
		13831 => '1',
		13832 => '0',
		13833 => '0',
		13834 => '1',
		13835 => '1',
		13836 => '1',
		13837 => '0',
		13838 => '0',
		13839 => '1',
		13840 => '1',
		13841 => '1',
		13842 => '0',
		13843 => '0',
		13844 => '1',
		13845 => '1',
		13846 => '1',
		13847 => '0',
		13848 => '0',
		13849 => '1',
		13850 => '1',
		13851 => '1',
		13852 => '0',
		13853 => '0',
		13854 => '1',
		13855 => '1',
		13856 => '1',
		13857 => '0',
		13858 => '0',
		13859 => '1',
		13860 => '1',
		13861 => '1',
		13862 => '0',
		13863 => '0',
		13864 => '0',
		13865 => '0',
		13866 => '0',
		13867 => '1',
		13868 => '1',
		13869 => '1',
		13870 => '0',
		13871 => '1',
		13872 => '1',
		13873 => '1',
		13874 => '0',
		13875 => '0',
		13876 => '0',
		13877 => '0',
		13878 => '0',
		13879 => '1',
		13880 => '1',
		13881 => '1',
		13882 => '0',
		13883 => '0',
		13884 => '1',
		13885 => '1',
		13886 => '1',
		13887 => '0',
		13888 => '0',
		13889 => '1',
		13890 => '1',
		13891 => '1',
		13892 => '0',
		13893 => '0',
		13894 => '1',
		13895 => '1',
		13896 => '1',
		13897 => '0',
		13898 => '0',
		13899 => '1',
		13900 => '1',
		13901 => '1',
		13902 => '0',
		13903 => '0',
		13904 => '1',
		13905 => '1',
		13906 => '1',
		13907 => '0',
		13908 => '0',
		13909 => '1',
		13910 => '1',
		13911 => '1',
		13912 => '0',
		13913 => '0',
		13914 => '1',
		13915 => '1',
		13916 => '1',
		13917 => '0',
		13918 => '0',
		13919 => '1',
		13920 => '1',
		13921 => '1',
		13922 => '0',
		13923 => '0',
		13924 => '1',
		13925 => '1',
		13926 => '1',
		13927 => '1',
		13928 => '1',
		13929 => '1',
		13930 => '1',
		13931 => '1',
		13932 => '0',
		13933 => '0',
		13934 => '1',
		13935 => '1',
		13936 => '1',
		13937 => '1',
		13938 => '1',
		13939 => '1',
		13940 => '1',
		13941 => '1',
		13942 => '0',
		13943 => '0',
		13952 => '1',
		13953 => '1',
		13954 => '1',
		13955 => '1',
		13956 => '1',
		13957 => '0',
		13958 => '0',
		13959 => '0',
		13960 => '1',
		13961 => '1',
		13962 => '1',
		13963 => '1',
		13964 => '1',
		13965 => '0',
		13966 => '0',
		13967 => '1',
		13968 => '1',
		13969 => '1',
		13970 => '0',
		13971 => '0',
		13972 => '1',
		13973 => '1',
		13974 => '1',
		13975 => '0',
		13976 => '0',
		13977 => '1',
		13978 => '1',
		13979 => '1',
		13980 => '0',
		13981 => '0',
		13982 => '0',
		13983 => '0',
		13984 => '0',
		13985 => '0',
		13986 => '0',
		13987 => '1',
		13988 => '1',
		13989 => '1',
		13990 => '0',
		13991 => '0',
		13992 => '0',
		13993 => '0',
		13994 => '0',
		13995 => '1',
		13996 => '1',
		13997 => '1',
		13998 => '0',
		13999 => '1',
		14000 => '1',
		14001 => '1',
		14002 => '0',
		14003 => '0',
		14004 => '0',
		14005 => '0',
		14006 => '0',
		14007 => '1',
		14008 => '1',
		14009 => '1',
		14010 => '0',
		14011 => '0',
		14012 => '0',
		14013 => '0',
		14014 => '0',
		14015 => '0',
		14016 => '0',
		14017 => '1',
		14018 => '1',
		14019 => '1',
		14020 => '0',
		14021 => '0',
		14022 => '1',
		14023 => '1',
		14024 => '1',
		14025 => '0',
		14026 => '0',
		14027 => '1',
		14028 => '1',
		14029 => '1',
		14030 => '0',
		14031 => '0',
		14032 => '1',
		14033 => '1',
		14034 => '1',
		14035 => '0',
		14036 => '0',
		14037 => '1',
		14038 => '1',
		14039 => '1',
		14040 => '0',
		14041 => '0',
		14042 => '1',
		14043 => '1',
		14044 => '1',
		14045 => '0',
		14046 => '0',
		14047 => '1',
		14048 => '1',
		14049 => '1',
		14050 => '0',
		14051 => '0',
		14052 => '0',
		14053 => '0',
		14054 => '0',
		14055 => '0',
		14056 => '0',
		14057 => '1',
		14058 => '1',
		14059 => '1',
		14060 => '0',
		14061 => '0',
		14062 => '1',
		14063 => '1',
		14064 => '1',
		14065 => '0',
		14066 => '0',
		14067 => '1',
		14068 => '1',
		14069 => '1',
		14070 => '0',
		14071 => '0',
		14080 => '1',
		14081 => '1',
		14082 => '1',
		14083 => '1',
		14084 => '1',
		14085 => '0',
		14086 => '0',
		14087 => '0',
		14088 => '1',
		14089 => '1',
		14090 => '1',
		14091 => '1',
		14092 => '1',
		14093 => '0',
		14094 => '0',
		14095 => '1',
		14096 => '1',
		14097 => '1',
		14098 => '0',
		14099 => '0',
		14100 => '1',
		14101 => '1',
		14102 => '1',
		14103 => '0',
		14104 => '0',
		14105 => '1',
		14106 => '1',
		14107 => '1',
		14108 => '0',
		14109 => '0',
		14110 => '0',
		14111 => '0',
		14112 => '0',
		14113 => '0',
		14114 => '0',
		14115 => '1',
		14116 => '1',
		14117 => '1',
		14118 => '0',
		14119 => '0',
		14120 => '0',
		14121 => '0',
		14122 => '0',
		14123 => '1',
		14124 => '1',
		14125 => '1',
		14126 => '0',
		14127 => '1',
		14128 => '1',
		14129 => '1',
		14130 => '0',
		14131 => '0',
		14132 => '0',
		14133 => '0',
		14134 => '0',
		14135 => '1',
		14136 => '1',
		14137 => '1',
		14138 => '0',
		14139 => '0',
		14140 => '0',
		14141 => '0',
		14142 => '0',
		14143 => '0',
		14144 => '0',
		14145 => '1',
		14146 => '1',
		14147 => '1',
		14148 => '0',
		14149 => '0',
		14150 => '1',
		14151 => '1',
		14152 => '1',
		14153 => '0',
		14154 => '0',
		14155 => '1',
		14156 => '1',
		14157 => '1',
		14158 => '0',
		14159 => '0',
		14160 => '1',
		14161 => '1',
		14162 => '1',
		14163 => '0',
		14164 => '0',
		14165 => '1',
		14166 => '1',
		14167 => '1',
		14168 => '0',
		14169 => '0',
		14170 => '1',
		14171 => '1',
		14172 => '1',
		14173 => '0',
		14174 => '0',
		14175 => '1',
		14176 => '1',
		14177 => '1',
		14178 => '0',
		14179 => '0',
		14180 => '0',
		14181 => '0',
		14182 => '0',
		14183 => '0',
		14184 => '0',
		14185 => '1',
		14186 => '1',
		14187 => '1',
		14188 => '0',
		14189 => '0',
		14190 => '1',
		14191 => '1',
		14192 => '1',
		14193 => '0',
		14194 => '0',
		14195 => '1',
		14196 => '1',
		14197 => '1',
		14198 => '0',
		14199 => '0',
		14208 => '0',
		14209 => '0',
		14210 => '0',
		14211 => '1',
		14212 => '1',
		14213 => '1',
		14214 => '1',
		14215 => '1',
		14216 => '1',
		14217 => '1',
		14218 => '0',
		14219 => '0',
		14220 => '0',
		14221 => '0',
		14222 => '0',
		14223 => '1',
		14224 => '1',
		14225 => '1',
		14226 => '1',
		14227 => '1',
		14228 => '1',
		14229 => '1',
		14230 => '1',
		14231 => '0',
		14232 => '0',
		14233 => '1',
		14234 => '1',
		14235 => '1',
		14236 => '1',
		14237 => '1',
		14238 => '1',
		14239 => '1',
		14240 => '1',
		14241 => '1',
		14242 => '1',
		14243 => '1',
		14244 => '1',
		14245 => '1',
		14246 => '0',
		14247 => '0',
		14248 => '0',
		14249 => '0',
		14250 => '0',
		14251 => '1',
		14252 => '1',
		14253 => '1',
		14254 => '1',
		14255 => '1',
		14256 => '1',
		14257 => '1',
		14258 => '0',
		14259 => '0',
		14260 => '0',
		14261 => '0',
		14262 => '0',
		14263 => '1',
		14264 => '1',
		14265 => '1',
		14266 => '1',
		14267 => '1',
		14268 => '1',
		14269 => '1',
		14270 => '1',
		14271 => '1',
		14272 => '1',
		14273 => '1',
		14274 => '1',
		14275 => '1',
		14276 => '0',
		14277 => '0',
		14278 => '1',
		14279 => '1',
		14280 => '1',
		14281 => '1',
		14282 => '1',
		14283 => '1',
		14284 => '1',
		14285 => '1',
		14286 => '0',
		14287 => '0',
		14288 => '1',
		14289 => '1',
		14290 => '1',
		14291 => '1',
		14292 => '1',
		14293 => '1',
		14294 => '1',
		14295 => '1',
		14296 => '1',
		14297 => '1',
		14298 => '1',
		14299 => '1',
		14300 => '1',
		14301 => '0',
		14302 => '0',
		14303 => '1',
		14304 => '1',
		14305 => '1',
		14306 => '1',
		14307 => '1',
		14308 => '1',
		14309 => '1',
		14310 => '1',
		14311 => '1',
		14312 => '1',
		14313 => '1',
		14314 => '1',
		14315 => '1',
		14316 => '0',
		14317 => '0',
		14318 => '1',
		14319 => '1',
		14320 => '1',
		14321 => '1',
		14322 => '1',
		14323 => '1',
		14324 => '1',
		14325 => '1',
		14326 => '0',
		14327 => '0',
		14336 => '0',
		14337 => '0',
		14338 => '0',
		14339 => '1',
		14340 => '1',
		14341 => '1',
		14342 => '1',
		14343 => '1',
		14344 => '1',
		14345 => '1',
		14346 => '0',
		14347 => '0',
		14348 => '0',
		14349 => '0',
		14350 => '0',
		14351 => '1',
		14352 => '1',
		14353 => '1',
		14354 => '1',
		14355 => '1',
		14356 => '1',
		14357 => '1',
		14358 => '1',
		14359 => '0',
		14360 => '0',
		14361 => '1',
		14362 => '1',
		14363 => '1',
		14364 => '1',
		14365 => '1',
		14366 => '1',
		14367 => '1',
		14368 => '1',
		14369 => '1',
		14370 => '1',
		14371 => '1',
		14372 => '1',
		14373 => '1',
		14374 => '0',
		14375 => '0',
		14376 => '0',
		14377 => '0',
		14378 => '0',
		14379 => '1',
		14380 => '1',
		14381 => '1',
		14382 => '1',
		14383 => '1',
		14384 => '1',
		14385 => '1',
		14386 => '0',
		14387 => '0',
		14388 => '0',
		14389 => '0',
		14390 => '0',
		14391 => '1',
		14392 => '1',
		14393 => '1',
		14394 => '1',
		14395 => '1',
		14396 => '1',
		14397 => '1',
		14398 => '1',
		14399 => '1',
		14400 => '1',
		14401 => '1',
		14402 => '1',
		14403 => '1',
		14404 => '0',
		14405 => '0',
		14406 => '1',
		14407 => '1',
		14408 => '1',
		14409 => '1',
		14410 => '1',
		14411 => '1',
		14412 => '1',
		14413 => '1',
		14414 => '0',
		14415 => '0',
		14416 => '1',
		14417 => '1',
		14418 => '1',
		14419 => '1',
		14420 => '1',
		14421 => '1',
		14422 => '1',
		14423 => '1',
		14424 => '1',
		14425 => '1',
		14426 => '1',
		14427 => '1',
		14428 => '1',
		14429 => '0',
		14430 => '0',
		14431 => '1',
		14432 => '1',
		14433 => '1',
		14434 => '1',
		14435 => '1',
		14436 => '1',
		14437 => '1',
		14438 => '1',
		14439 => '1',
		14440 => '1',
		14441 => '1',
		14442 => '1',
		14443 => '1',
		14444 => '0',
		14445 => '0',
		14446 => '1',
		14447 => '1',
		14448 => '1',
		14449 => '1',
		14450 => '1',
		14451 => '1',
		14452 => '1',
		14453 => '1',
		14454 => '0',
		14455 => '0',
		14464 => '0',
		14465 => '0',
		14466 => '0',
		14467 => '1',
		14468 => '1',
		14469 => '1',
		14470 => '1',
		14471 => '1',
		14472 => '1',
		14473 => '1',
		14474 => '0',
		14475 => '0',
		14476 => '0',
		14477 => '0',
		14478 => '0',
		14479 => '1',
		14480 => '1',
		14481 => '1',
		14482 => '1',
		14483 => '1',
		14484 => '1',
		14485 => '1',
		14486 => '1',
		14487 => '0',
		14488 => '0',
		14489 => '1',
		14490 => '1',
		14491 => '1',
		14492 => '1',
		14493 => '1',
		14494 => '1',
		14495 => '1',
		14496 => '1',
		14497 => '1',
		14498 => '1',
		14499 => '1',
		14500 => '1',
		14501 => '1',
		14502 => '0',
		14503 => '0',
		14504 => '0',
		14505 => '0',
		14506 => '0',
		14507 => '1',
		14508 => '1',
		14509 => '1',
		14510 => '1',
		14511 => '1',
		14512 => '1',
		14513 => '1',
		14514 => '0',
		14515 => '0',
		14516 => '0',
		14517 => '0',
		14518 => '0',
		14519 => '1',
		14520 => '1',
		14521 => '1',
		14522 => '1',
		14523 => '1',
		14524 => '1',
		14525 => '1',
		14526 => '1',
		14527 => '1',
		14528 => '1',
		14529 => '1',
		14530 => '1',
		14531 => '1',
		14532 => '0',
		14533 => '0',
		14534 => '1',
		14535 => '1',
		14536 => '1',
		14537 => '1',
		14538 => '1',
		14539 => '1',
		14540 => '1',
		14541 => '1',
		14542 => '0',
		14543 => '0',
		14544 => '1',
		14545 => '1',
		14546 => '1',
		14547 => '1',
		14548 => '1',
		14549 => '1',
		14550 => '1',
		14551 => '1',
		14552 => '1',
		14553 => '1',
		14554 => '1',
		14555 => '1',
		14556 => '1',
		14557 => '0',
		14558 => '0',
		14559 => '1',
		14560 => '1',
		14561 => '1',
		14562 => '1',
		14563 => '1',
		14564 => '1',
		14565 => '1',
		14566 => '1',
		14567 => '1',
		14568 => '1',
		14569 => '1',
		14570 => '1',
		14571 => '1',
		14572 => '0',
		14573 => '0',
		14574 => '1',
		14575 => '1',
		14576 => '1',
		14577 => '1',
		14578 => '1',
		14579 => '1',
		14580 => '1',
		14581 => '1',
		14582 => '0',
		14583 => '0',
		14592 => '0',
		14593 => '0',
		14594 => '0',
		14595 => '0',
		14596 => '0',
		14597 => '0',
		14598 => '0',
		14599 => '0',
		14600 => '0',
		14601 => '0',
		14602 => '0',
		14603 => '0',
		14604 => '0',
		14605 => '0',
		14606 => '0',
		14607 => '0',
		14608 => '0',
		14609 => '0',
		14610 => '0',
		14611 => '0',
		14612 => '0',
		14613 => '0',
		14614 => '0',
		14615 => '0',
		14616 => '0',
		14617 => '0',
		14618 => '0',
		14619 => '0',
		14620 => '0',
		14621 => '0',
		14622 => '0',
		14623 => '0',
		14624 => '0',
		14625 => '0',
		14626 => '0',
		14627 => '0',
		14628 => '0',
		14629 => '0',
		14630 => '0',
		14631 => '0',
		14632 => '0',
		14633 => '0',
		14634 => '0',
		14635 => '0',
		14636 => '0',
		14637 => '0',
		14638 => '0',
		14639 => '0',
		14640 => '0',
		14641 => '0',
		14642 => '0',
		14643 => '0',
		14644 => '0',
		14645 => '0',
		14646 => '0',
		14647 => '0',
		14648 => '0',
		14649 => '0',
		14650 => '0',
		14651 => '0',
		14652 => '0',
		14653 => '0',
		14654 => '0',
		14655 => '0',
		14656 => '0',
		14657 => '0',
		14658 => '0',
		14659 => '0',
		14660 => '0',
		14661 => '0',
		14662 => '0',
		14663 => '0',
		14664 => '0',
		14665 => '0',
		14666 => '0',
		14667 => '0',
		14668 => '0',
		14669 => '0',
		14670 => '0',
		14671 => '0',
		14672 => '0',
		14673 => '0',
		14674 => '0',
		14675 => '0',
		14676 => '0',
		14677 => '0',
		14678 => '0',
		14679 => '0',
		14680 => '0',
		14681 => '0',
		14682 => '0',
		14683 => '0',
		14684 => '0',
		14685 => '0',
		14686 => '0',
		14687 => '0',
		14688 => '0',
		14689 => '0',
		14690 => '0',
		14691 => '0',
		14692 => '0',
		14693 => '0',
		14694 => '0',
		14695 => '0',
		14696 => '0',
		14697 => '0',
		14698 => '0',
		14699 => '0',
		14700 => '0',
		14701 => '0',
		14702 => '0',
		14703 => '0',
		14704 => '0',
		14705 => '0',
		14706 => '0',
		14707 => '0',
		14708 => '0',
		14709 => '0',
		14710 => '0',
		14711 => '0',
		14720 => '0',
		14721 => '0',
		14722 => '0',
		14723 => '0',
		14724 => '0',
		14725 => '0',
		14726 => '0',
		14727 => '0',
		14728 => '0',
		14729 => '0',
		14730 => '0',
		14731 => '0',
		14732 => '0',
		14733 => '0',
		14734 => '0',
		14735 => '0',
		14736 => '0',
		14737 => '0',
		14738 => '0',
		14739 => '0',
		14740 => '0',
		14741 => '0',
		14742 => '0',
		14743 => '0',
		14744 => '0',
		14745 => '0',
		14746 => '0',
		14747 => '0',
		14748 => '0',
		14749 => '0',
		14750 => '0',
		14751 => '0',
		14752 => '0',
		14753 => '0',
		14754 => '0',
		14755 => '0',
		14756 => '0',
		14757 => '0',
		14758 => '0',
		14759 => '0',
		14760 => '0',
		14761 => '0',
		14762 => '0',
		14763 => '0',
		14764 => '0',
		14765 => '0',
		14766 => '0',
		14767 => '0',
		14768 => '0',
		14769 => '0',
		14770 => '0',
		14771 => '0',
		14772 => '0',
		14773 => '0',
		14774 => '0',
		14775 => '0',
		14776 => '0',
		14777 => '0',
		14778 => '0',
		14779 => '0',
		14780 => '0',
		14781 => '0',
		14782 => '0',
		14783 => '0',
		14784 => '0',
		14785 => '0',
		14786 => '0',
		14787 => '0',
		14788 => '0',
		14789 => '0',
		14790 => '0',
		14791 => '0',
		14792 => '0',
		14793 => '0',
		14794 => '0',
		14795 => '0',
		14796 => '0',
		14797 => '0',
		14798 => '0',
		14799 => '0',
		14800 => '0',
		14801 => '0',
		14802 => '0',
		14803 => '0',
		14804 => '0',
		14805 => '0',
		14806 => '0',
		14807 => '0',
		14808 => '0',
		14809 => '0',
		14810 => '0',
		14811 => '0',
		14812 => '0',
		14813 => '0',
		14814 => '0',
		14815 => '0',
		14816 => '0',
		14817 => '0',
		14818 => '0',
		14819 => '0',
		14820 => '0',
		14821 => '0',
		14822 => '0',
		14823 => '0',
		14824 => '0',
		14825 => '0',
		14826 => '0',
		14827 => '0',
		14828 => '0',
		14829 => '0',
		14830 => '0',
		14831 => '0',
		14832 => '0',
		14833 => '0',
		14834 => '0',
		14835 => '0',
		14836 => '0',
		14837 => '0',
		14838 => '0',
		14839 => '0',
		14848 => '0',
		14849 => '0',
		14850 => '0',
		14851 => '0',
		14852 => '0',
		14853 => '0',
		14854 => '0',
		14855 => '0',
		14856 => '0',
		14857 => '0',
		14858 => '0',
		14859 => '0',
		14860 => '0',
		14861 => '0',
		14862 => '0',
		14863 => '0',
		14864 => '0',
		14865 => '0',
		14866 => '0',
		14867 => '0',
		14868 => '0',
		14869 => '0',
		14870 => '0',
		14871 => '0',
		14872 => '0',
		14873 => '0',
		14874 => '0',
		14875 => '0',
		14876 => '0',
		14877 => '0',
		14878 => '0',
		14879 => '0',
		14880 => '0',
		14881 => '0',
		14882 => '0',
		14883 => '0',
		14884 => '0',
		14885 => '0',
		14886 => '0',
		14887 => '0',
		14888 => '0',
		14889 => '0',
		14890 => '0',
		14891 => '0',
		14892 => '0',
		14893 => '0',
		14894 => '0',
		14895 => '0',
		14896 => '0',
		14897 => '0',
		14898 => '0',
		14899 => '0',
		14900 => '0',
		14901 => '0',
		14902 => '0',
		14903 => '0',
		14904 => '0',
		14905 => '0',
		14906 => '0',
		14907 => '0',
		14908 => '0',
		14909 => '0',
		14910 => '0',
		14911 => '0',
		14912 => '0',
		14913 => '0',
		14914 => '0',
		14915 => '0',
		14916 => '0',
		14917 => '0',
		14918 => '0',
		14919 => '0',
		14920 => '0',
		14921 => '0',
		14922 => '0',
		14923 => '0',
		14924 => '0',
		14925 => '0',
		14926 => '0',
		14927 => '0',
		14928 => '0',
		14929 => '0',
		14930 => '0',
		14931 => '0',
		14932 => '0',
		14933 => '0',
		14934 => '0',
		14935 => '0',
		14936 => '0',
		14937 => '0',
		14938 => '0',
		14939 => '0',
		14940 => '0',
		14941 => '0',
		14942 => '0',
		14943 => '0',
		14944 => '0',
		14945 => '0',
		14946 => '0',
		14947 => '0',
		14948 => '0',
		14949 => '0',
		14950 => '0',
		14951 => '0',
		14952 => '0',
		14953 => '0',
		14954 => '0',
		14955 => '0',
		14956 => '0',
		14957 => '0',
		14958 => '0',
		14959 => '0',
		14960 => '0',
		14961 => '0',
		14962 => '0',
		14963 => '0',
		14964 => '0',
		14965 => '0',
		14966 => '0',
		14967 => '0',
		14976 => '0',
		14977 => '0',
		14978 => '0',
		14979 => '0',
		14980 => '0',
		14981 => '0',
		14982 => '0',
		14983 => '0',
		14984 => '0',
		14985 => '0',
		14986 => '0',
		14987 => '0',
		14988 => '0',
		14989 => '0',
		14990 => '0',
		14991 => '0',
		14992 => '0',
		14993 => '0',
		14994 => '0',
		14995 => '0',
		14996 => '0',
		14997 => '0',
		14998 => '0',
		14999 => '0',
		15000 => '0',
		15001 => '0',
		15002 => '0',
		15003 => '0',
		15004 => '0',
		15005 => '0',
		15006 => '0',
		15007 => '0',
		15008 => '0',
		15009 => '0',
		15010 => '0',
		15011 => '0',
		15012 => '0',
		15013 => '0',
		15014 => '0',
		15015 => '0',
		15016 => '0',
		15017 => '0',
		15018 => '0',
		15019 => '0',
		15020 => '0',
		15021 => '0',
		15022 => '0',
		15023 => '0',
		15024 => '0',
		15025 => '0',
		15026 => '0',
		15027 => '0',
		15028 => '0',
		15029 => '0',
		15030 => '0',
		15031 => '0',
		15032 => '0',
		15033 => '0',
		15034 => '0',
		15035 => '0',
		15036 => '0',
		15037 => '0',
		15038 => '0',
		15039 => '0',
		15040 => '0',
		15041 => '0',
		15042 => '0',
		15043 => '0',
		15044 => '0',
		15045 => '0',
		15046 => '0',
		15047 => '0',
		15048 => '0',
		15049 => '0',
		15050 => '0',
		15051 => '0',
		15052 => '0',
		15053 => '0',
		15054 => '0',
		15055 => '0',
		15056 => '0',
		15057 => '0',
		15058 => '0',
		15059 => '0',
		15060 => '0',
		15061 => '0',
		15062 => '0',
		15063 => '0',
		15064 => '0',
		15065 => '0',
		15066 => '0',
		15067 => '0',
		15068 => '0',
		15069 => '0',
		15070 => '0',
		15071 => '0',
		15072 => '0',
		15073 => '0',
		15074 => '0',
		15075 => '0',
		15076 => '0',
		15077 => '0',
		15078 => '0',
		15079 => '0',
		15080 => '0',
		15081 => '0',
		15082 => '0',
		15083 => '0',
		15084 => '0',
		15085 => '0',
		15086 => '0',
		15087 => '0',
		15088 => '0',
		15089 => '0',
		15090 => '0',
		15091 => '0',
		15092 => '0',
		15093 => '0',
		15094 => '0',
		15095 => '0',
		15104 => '0',
		15105 => '0',
		15106 => '0',
		15107 => '0',
		15108 => '0',
		15109 => '0',
		15110 => '0',
		15111 => '0',
		15112 => '0',
		15113 => '0',
		15114 => '0',
		15115 => '0',
		15116 => '0',
		15117 => '0',
		15118 => '0',
		15119 => '0',
		15120 => '0',
		15121 => '0',
		15122 => '0',
		15123 => '0',
		15124 => '0',
		15125 => '0',
		15126 => '0',
		15127 => '0',
		15128 => '0',
		15129 => '0',
		15130 => '0',
		15131 => '0',
		15132 => '0',
		15133 => '0',
		15134 => '0',
		15135 => '0',
		15136 => '0',
		15137 => '0',
		15138 => '0',
		15139 => '0',
		15140 => '0',
		15141 => '0',
		15142 => '0',
		15143 => '0',
		15144 => '0',
		15145 => '0',
		15146 => '0',
		15147 => '0',
		15148 => '0',
		15149 => '0',
		15150 => '0',
		15151 => '0',
		15152 => '0',
		15153 => '0',
		15154 => '0',
		15155 => '0',
		15156 => '0',
		15157 => '0',
		15158 => '0',
		15159 => '0',
		15160 => '0',
		15161 => '0',
		15162 => '0',
		15163 => '0',
		15164 => '0',
		15165 => '0',
		15166 => '0',
		15167 => '0',
		15168 => '0',
		15169 => '0',
		15170 => '0',
		15171 => '0',
		15172 => '0',
		15173 => '0',
		15174 => '0',
		15175 => '0',
		15176 => '0',
		15177 => '0',
		15178 => '0',
		15179 => '0',
		15180 => '0',
		15181 => '0',
		15182 => '0',
		15183 => '0',
		15184 => '0',
		15185 => '0',
		15186 => '0',
		15187 => '0',
		15188 => '0',
		15189 => '0',
		15190 => '0',
		15191 => '0',
		15192 => '0',
		15193 => '0',
		15194 => '0',
		15195 => '0',
		15196 => '0',
		15197 => '0',
		15198 => '0',
		15199 => '0',
		15200 => '0',
		15201 => '0',
		15202 => '0',
		15203 => '0',
		15204 => '0',
		15205 => '0',
		15206 => '0',
		15207 => '0',
		15208 => '0',
		15209 => '0',
		15210 => '0',
		15211 => '0',
		15212 => '0',
		15213 => '0',
		15214 => '0',
		15215 => '0',
		15216 => '0',
		15217 => '0',
		15218 => '0',
		15219 => '0',
		15220 => '0',
		15221 => '0',
		15222 => '0',
		15223 => '0',
		15232 => '0',
		15233 => '0',
		15234 => '0',
		15235 => '0',
		15236 => '0',
		15237 => '0',
		15238 => '0',
		15239 => '0',
		15240 => '0',
		15241 => '0',
		15242 => '0',
		15243 => '0',
		15244 => '0',
		15245 => '0',
		15246 => '0',
		15247 => '0',
		15248 => '0',
		15249 => '0',
		15250 => '0',
		15251 => '0',
		15252 => '0',
		15253 => '0',
		15254 => '0',
		15255 => '0',
		15256 => '0',
		15257 => '0',
		15258 => '0',
		15259 => '0',
		15260 => '0',
		15261 => '0',
		15262 => '0',
		15263 => '0',
		15264 => '0',
		15265 => '0',
		15266 => '0',
		15267 => '0',
		15268 => '0',
		15269 => '0',
		15270 => '0',
		15271 => '0',
		15272 => '0',
		15273 => '0',
		15274 => '0',
		15275 => '0',
		15276 => '0',
		15277 => '0',
		15278 => '0',
		15279 => '0',
		15280 => '0',
		15281 => '0',
		15282 => '0',
		15283 => '0',
		15284 => '0',
		15285 => '0',
		15286 => '0',
		15287 => '0',
		15288 => '0',
		15289 => '0',
		15290 => '0',
		15291 => '0',
		15292 => '0',
		15293 => '0',
		15294 => '0',
		15295 => '0',
		15296 => '0',
		15297 => '0',
		15298 => '0',
		15299 => '0',
		15300 => '0',
		15301 => '0',
		15302 => '0',
		15303 => '0',
		15304 => '0',
		15305 => '0',
		15306 => '0',
		15307 => '0',
		15308 => '0',
		15309 => '0',
		15310 => '0',
		15311 => '0',
		15312 => '0',
		15313 => '0',
		15314 => '0',
		15315 => '0',
		15316 => '0',
		15317 => '0',
		15318 => '0',
		15319 => '0',
		15320 => '0',
		15321 => '0',
		15322 => '0',
		15323 => '0',
		15324 => '0',
		15325 => '0',
		15326 => '0',
		15327 => '0',
		15328 => '0',
		15329 => '0',
		15330 => '0',
		15331 => '0',
		15332 => '0',
		15333 => '0',
		15334 => '0',
		15335 => '0',
		15336 => '0',
		15337 => '0',
		15338 => '0',
		15339 => '0',
		15340 => '0',
		15341 => '0',
		15342 => '0',
		15343 => '0',
		15344 => '0',
		15345 => '0',
		15346 => '0',
		15347 => '0',
		15348 => '0',
		15349 => '0',
		15350 => '0',
		15351 => '0',

	others => '0'
);

begin
	
	-- process ROM
	process (CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (EN = '1') then
				DATA <= ROM(to_integer(unsigned(ADDR)));
			end if;
		end if;
	end process;
	
end Behavioral;

