----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:16:29 04/19/2013 
-- Design Name: 
-- Module Name:    VRAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity VRAM is
	port (Clk		: in 	std_logic;
			CE			: in 	std_logic;
			Enable_w	: in 	std_logic;
			Addr_w	: in 	std_logic_vector	(18 downto 0);
			Addr_r	: in 	std_logic_vector	(18 downto 0);
			Data_in	: in 	std_logic_vector	(7 downto 0);
			Data_out	: out std_logic_vector	(7 downto 0));
end VRAM;

architecture Behavioral of VRAM is
	type ram_type is array ((2**16)-1 downto 0) of std_logic_vector (7 downto 0);
	signal VRAM: ram_type := (
		19555 to 19994 => "11111111",
		20579 to 21018 => "11111111",
		21603 to 22042 => "11111111",
		22627 to 23066 => "11111111",
		23651 to 24090 => "11111111",
		24675 to 24679 => "11111111",
		24820 to 24824 => "11111111",
		24965 to 24969 => "11111111",
		25110 to 25114 => "11111111",
		25699 to 25703 => "11111111",
		25844 to 25848 => "11111111",
		25989 to 25993 => "11111111",
		26134 to 26138 => "11111111",
		26723 to 26727 => "11111111",
		26868 to 26872 => "11111111",
		27013 to 27017 => "11111111",
		27158 to 27162 => "11111111",
		27747 to 27751 => "11111111",
		27892 to 27896 => "11111111",
		28037 to 28041 => "11111111",
		28182 to 28186 => "11111111",
		28771 to 28775 => "11111111",
		28916 to 28920 => "11111111",
		29061 to 29065 => "11111111",
		29206 to 29210 => "11111111",
		29795 to 29799 => "11111111",
		29940 to 29944 => "11111111",
		30085 to 30089 => "11111111",
		30230 to 30234 => "11111111",
		30819 to 30823 => "11111111",
		30964 to 30968 => "11111111",
		31109 to 31113 => "11111111",
		31254 to 31258 => "11111111",
		31843 to 31847 => "11111111",
		31988 to 31992 => "11111111",
		32133 to 32137 => "11111111",
		32278 to 32282 => "11111111",
		32867 to 32871 => "11111111",
		33012 to 33016 => "11111111",
		33157 to 33161 => "11111111",
		33302 to 33306 => "11111111",
		33891 to 33895 => "11111111",
		34036 to 34040 => "11111111",
		34181 to 34185 => "11111111",
		34326 to 34330 => "11111111",
		34915 to 34919 => "11111111",
		35060 to 35064 => "11111111",
		35205 to 35209 => "11111111",
		35350 to 35354 => "11111111",
		35939 to 35943 => "11111111",
		36084 to 36088 => "11111111",
		36229 to 36233 => "11111111",
		36374 to 36378 => "11111111",
		36963 to 36967 => "11111111",
		37108 to 37112 => "11111111",
		37253 to 37257 => "11111111",
		37398 to 37402 => "11111111",
		37987 to 37991 => "11111111",
		38132 to 38136 => "11111111",
		38277 to 38281 => "11111111",
		38422 to 38426 => "11111111",
		39011 to 39015 => "11111111",
		39156 to 39160 => "11111111",
		39301 to 39305 => "11111111",
		39446 to 39450 => "11111111",
		40035 to 40039 => "11111111",
		40180 to 40184 => "11111111",
		40325 to 40329 => "11111111",
		40470 to 40474 => "11111111",
		41059 to 41063 => "11111111",
		41204 to 41208 => "11111111",
		41349 to 41353 => "11111111",
		41494 to 41498 => "11111111",
		42083 to 42087 => "11111111",
		42228 to 42232 => "11111111",
		42373 to 42377 => "11111111",
		42518 to 42522 => "11111111",
		43107 to 43111 => "11111111",
		43252 to 43256 => "11111111",
		43397 to 43401 => "11111111",
		43542 to 43546 => "11111111",
		44131 to 44135 => "11111111",
		44276 to 44280 => "11111111",
		44421 to 44425 => "11111111",
		44566 to 44570 => "11111111",
		45155 to 45159 => "11111111",
		45300 to 45304 => "11111111",
		45445 to 45449 => "11111111",
		45590 to 45594 => "11111111",
		46179 to 46183 => "11111111",
		46324 to 46328 => "11111111",
		46469 to 46473 => "11111111",
		46614 to 46618 => "11111111",
		47203 to 47207 => "11111111",
		47348 to 47352 => "11111111",
		47493 to 47497 => "11111111",
		47638 to 47642 => "11111111",
		48227 to 48231 => "11111111",
		48372 to 48376 => "11111111",
		48517 to 48521 => "11111111",
		48662 to 48666 => "11111111",
		49251 to 49255 => "11111111",
		49396 to 49400 => "11111111",
		49541 to 49545 => "11111111",
		49686 to 49690 => "11111111",
		50275 to 50279 => "11111111",
		50420 to 50424 => "11111111",
		50565 to 50569 => "11111111",
		50710 to 50714 => "11111111",
		51299 to 51303 => "11111111",
		51444 to 51448 => "11111111",
		51589 to 51593 => "11111111",
		51734 to 51738 => "11111111",
		52323 to 52327 => "11111111",
		52468 to 52472 => "11111111",
		52613 to 52617 => "11111111",
		52758 to 52762 => "11111111",
		53347 to 53351 => "11111111",
		53492 to 53496 => "11111111",
		53637 to 53641 => "11111111",
		53782 to 53786 => "11111111",
		54371 to 54375 => "11111111",
		54516 to 54520 => "11111111",
		54661 to 54665 => "11111111",
		54806 to 54810 => "11111111",
		55395 to 55399 => "11111111",
		55540 to 55544 => "11111111",
		55685 to 55689 => "11111111",
		55830 to 55834 => "11111111",
		56419 to 56423 => "11111111",
		56564 to 56568 => "11111111",
		56709 to 56713 => "11111111",
		56854 to 56858 => "11111111",
		57443 to 57447 => "11111111",
		57588 to 57592 => "11111111",
		57733 to 57737 => "11111111",
		57878 to 57882 => "11111111",
		58467 to 58471 => "11111111",
		58612 to 58616 => "11111111",
		58757 to 58761 => "11111111",
		58902 to 58906 => "11111111",
		59491 to 59495 => "11111111",
		59636 to 59640 => "11111111",
		59781 to 59785 => "11111111",
		59926 to 59930 => "11111111",
		60515 to 60519 => "11111111",
		60660 to 60664 => "11111111",
		60805 to 60809 => "11111111",
		60950 to 60954 => "11111111",
		61539 to 61543 => "11111111",
		61684 to 61688 => "11111111",
		61829 to 61833 => "11111111",
		61974 to 61978 => "11111111",
		62563 to 62567 => "11111111",
		62708 to 62712 => "11111111",
		62853 to 62857 => "11111111",
		62998 to 63002 => "11111111",
		63587 to 63591 => "11111111",
		63732 to 63736 => "11111111",
		63877 to 63881 => "11111111",
		64022 to 64026 => "11111111",
		64611 to 64615 => "11111111",
		64756 to 64760 => "11111111",
		64901 to 64905 => "11111111",
		65046 to 65050 => "11111111",
--		65635 to 65639 => "11111111",
--		65780 to 65784 => "11111111",
--		65925 to 65929 => "11111111",
--		66070 to 66074 => "11111111",
--		66659 to 66663 => "11111111",
--		66804 to 66808 => "11111111",
--		66949 to 66953 => "11111111",
--		67094 to 67098 => "11111111",
--		67683 to 67687 => "11111111",
--		67828 to 67832 => "11111111",
--		67973 to 67977 => "11111111",
--		68118 to 68122 => "11111111",
--		68707 to 68711 => "11111111",
--		68852 to 68856 => "11111111",
--		68997 to 69001 => "11111111",
--		69142 to 69146 => "11111111",
--		69731 to 69735 => "11111111",
--		69876 to 69880 => "11111111",
--		70021 to 70025 => "11111111",
--		70166 to 70170 => "11111111",
--		70755 to 70759 => "11111111",
--		70900 to 70904 => "11111111",
--		71045 to 71049 => "11111111",
--		71190 to 71194 => "11111111",
--		71779 to 71783 => "11111111",
--		71924 to 71928 => "11111111",
--		72069 to 72073 => "11111111",
--		72214 to 72218 => "11111111",
--		72803 to 72807 => "11111111",
--		72948 to 72952 => "11111111",
--		73093 to 73097 => "11111111",
--		73238 to 73242 => "11111111",
--		73827 to 73831 => "11111111",
--		73972 to 73976 => "11111111",
--		74117 to 74121 => "11111111",
--		74262 to 74266 => "11111111",
--		74851 to 74855 => "11111111",
--		74996 to 75000 => "11111111",
--		75141 to 75145 => "11111111",
--		75286 to 75290 => "11111111",
--		75875 to 75879 => "11111111",
--		76020 to 76024 => "11111111",
--		76165 to 76169 => "11111111",
--		76310 to 76314 => "11111111",
--		76899 to 76903 => "11111111",
--		77044 to 77048 => "11111111",
--		77189 to 77193 => "11111111",
--		77334 to 77338 => "11111111",
--		77923 to 77927 => "11111111",
--		78068 to 78072 => "11111111",
--		78213 to 78217 => "11111111",
--		78358 to 78362 => "11111111",
--		78947 to 78951 => "11111111",
--		79092 to 79096 => "11111111",
--		79237 to 79241 => "11111111",
--		79382 to 79386 => "11111111",
--		79971 to 79975 => "11111111",
--		80116 to 80120 => "11111111",
--		80261 to 80265 => "11111111",
--		80406 to 80410 => "11111111",
--		80995 to 80999 => "11111111",
--		81140 to 81144 => "11111111",
--		81285 to 81289 => "11111111",
--		81430 to 81434 => "11111111",
--		82019 to 82023 => "11111111",
--		82164 to 82168 => "11111111",
--		82309 to 82313 => "11111111",
--		82454 to 82458 => "11111111",
--		83043 to 83047 => "11111111",
--		83188 to 83192 => "11111111",
--		83333 to 83337 => "11111111",
--		83478 to 83482 => "11111111",
--		84067 to 84071 => "11111111",
--		84212 to 84216 => "11111111",
--		84357 to 84361 => "11111111",
--		84502 to 84506 => "11111111",
--		85091 to 85095 => "11111111",
--		85236 to 85240 => "11111111",
--		85381 to 85385 => "11111111",
--		85526 to 85530 => "11111111",
--		86115 to 86119 => "11111111",
--		86260 to 86264 => "11111111",
--		86405 to 86409 => "11111111",
--		86550 to 86554 => "11111111",
--		87139 to 87143 => "11111111",
--		87284 to 87288 => "11111111",
--		87429 to 87433 => "11111111",
--		87574 to 87578 => "11111111",
--		88163 to 88167 => "11111111",
--		88308 to 88312 => "11111111",
--		88453 to 88457 => "11111111",
--		88598 to 88602 => "11111111",
--		89187 to 89191 => "11111111",
--		89332 to 89336 => "11111111",
--		89477 to 89481 => "11111111",
--		89622 to 89626 => "11111111",
--		90211 to 90215 => "11111111",
--		90356 to 90360 => "11111111",
--		90501 to 90505 => "11111111",
--		90646 to 90650 => "11111111",
--		91235 to 91239 => "11111111",
--		91380 to 91384 => "11111111",
--		91525 to 91529 => "11111111",
--		91670 to 91674 => "11111111",
--		92259 to 92263 => "11111111",
--		92404 to 92408 => "11111111",
--		92549 to 92553 => "11111111",
--		92694 to 92698 => "11111111",
--		93283 to 93287 => "11111111",
--		93428 to 93432 => "11111111",
--		93573 to 93577 => "11111111",
--		93718 to 93722 => "11111111",
--		94307 to 94311 => "11111111",
--		94452 to 94456 => "11111111",
--		94597 to 94601 => "11111111",
--		94742 to 94746 => "11111111",
--		95331 to 95335 => "11111111",
--		95476 to 95480 => "11111111",
--		95621 to 95625 => "11111111",
--		95766 to 95770 => "11111111",
--		96355 to 96359 => "11111111",
--		96500 to 96504 => "11111111",
--		96645 to 96649 => "11111111",
--		96790 to 96794 => "11111111",
--		97379 to 97383 => "11111111",
--		97524 to 97528 => "11111111",
--		97669 to 97673 => "11111111",
--		97814 to 97818 => "11111111",
--		98403 to 98407 => "11111111",
--		98548 to 98552 => "11111111",
--		98693 to 98697 => "11111111",
--		98838 to 98842 => "11111111",
--		99427 to 99431 => "11111111",
--		99572 to 99576 => "11111111",
--		99717 to 99721 => "11111111",
--		99862 to 99866 => "11111111",
--		100451 to 100455 => "11111111",
--		100596 to 100600 => "11111111",
--		100741 to 100745 => "11111111",
--		100886 to 100890 => "11111111",
--		101475 to 101479 => "11111111",
--		101620 to 101624 => "11111111",
--		101765 to 101769 => "11111111",
--		101910 to 101914 => "11111111",
--		102499 to 102503 => "11111111",
--		102644 to 102648 => "11111111",
--		102789 to 102793 => "11111111",
--		102934 to 102938 => "11111111",
--		103523 to 103527 => "11111111",
--		103668 to 103672 => "11111111",
--		103813 to 103817 => "11111111",
--		103958 to 103962 => "11111111",
--		104547 to 104551 => "11111111",
--		104692 to 104696 => "11111111",
--		104837 to 104841 => "11111111",
--		104982 to 104986 => "11111111",
--		105571 to 105575 => "11111111",
--		105716 to 105720 => "11111111",
--		105861 to 105865 => "11111111",
--		106006 to 106010 => "11111111",
--		106595 to 106599 => "11111111",
--		106740 to 106744 => "11111111",
--		106885 to 106889 => "11111111",
--		107030 to 107034 => "11111111",
--		107619 to 107623 => "11111111",
--		107764 to 107768 => "11111111",
--		107909 to 107913 => "11111111",
--		108054 to 108058 => "11111111",
--		108643 to 108647 => "11111111",
--		108788 to 108792 => "11111111",
--		108933 to 108937 => "11111111",
--		109078 to 109082 => "11111111",
--		109667 to 109671 => "11111111",
--		109812 to 109816 => "11111111",
--		109957 to 109961 => "11111111",
--		110102 to 110106 => "11111111",
--		110691 to 110695 => "11111111",
--		110836 to 110840 => "11111111",
--		110981 to 110985 => "11111111",
--		111126 to 111130 => "11111111",
--		111715 to 111719 => "11111111",
--		111860 to 111864 => "11111111",
--		112005 to 112009 => "11111111",
--		112150 to 112154 => "11111111",
--		112739 to 112743 => "11111111",
--		112884 to 112888 => "11111111",
--		113029 to 113033 => "11111111",
--		113174 to 113178 => "11111111",
--		113763 to 113767 => "11111111",
--		113908 to 113912 => "11111111",
--		114053 to 114057 => "11111111",
--		114198 to 114202 => "11111111",
--		114787 to 114791 => "11111111",
--		114932 to 114936 => "11111111",
--		115077 to 115081 => "11111111",
--		115222 to 115226 => "11111111",
--		115811 to 115815 => "11111111",
--		115956 to 115960 => "11111111",
--		116101 to 116105 => "11111111",
--		116246 to 116250 => "11111111",
--		116835 to 116839 => "11111111",
--		116980 to 116984 => "11111111",
--		117125 to 117129 => "11111111",
--		117270 to 117274 => "11111111",
--		117859 to 117863 => "11111111",
--		118004 to 118008 => "11111111",
--		118149 to 118153 => "11111111",
--		118294 to 118298 => "11111111",
--		118883 to 118887 => "11111111",
--		119028 to 119032 => "11111111",
--		119173 to 119177 => "11111111",
--		119318 to 119322 => "11111111",
--		119907 to 119911 => "11111111",
--		120052 to 120056 => "11111111",
--		120197 to 120201 => "11111111",
--		120342 to 120346 => "11111111",
--		120931 to 120935 => "11111111",
--		121076 to 121080 => "11111111",
--		121221 to 121225 => "11111111",
--		121366 to 121370 => "11111111",
--		121955 to 121959 => "11111111",
--		122100 to 122104 => "11111111",
--		122245 to 122249 => "11111111",
--		122390 to 122394 => "11111111",
--		122979 to 122983 => "11111111",
--		123124 to 123128 => "11111111",
--		123269 to 123273 => "11111111",
--		123414 to 123418 => "11111111",
--		124003 to 124007 => "11111111",
--		124148 to 124152 => "11111111",
--		124293 to 124297 => "11111111",
--		124438 to 124442 => "11111111",
--		125027 to 125031 => "11111111",
--		125172 to 125176 => "11111111",
--		125317 to 125321 => "11111111",
--		125462 to 125466 => "11111111",
--		126051 to 126055 => "11111111",
--		126196 to 126200 => "11111111",
--		126341 to 126345 => "11111111",
--		126486 to 126490 => "11111111",
--		127075 to 127079 => "11111111",
--		127220 to 127224 => "11111111",
--		127365 to 127369 => "11111111",
--		127510 to 127514 => "11111111",
--		128099 to 128103 => "11111111",
--		128244 to 128248 => "11111111",
--		128389 to 128393 => "11111111",
--		128534 to 128538 => "11111111",
--		129123 to 129127 => "11111111",
--		129268 to 129272 => "11111111",
--		129413 to 129417 => "11111111",
--		129558 to 129562 => "11111111",
--		130147 to 130151 => "11111111",
--		130292 to 130296 => "11111111",
--		130437 to 130441 => "11111111",
--		130582 to 130586 => "11111111",
--		131171 to 131175 => "11111111",
--		131316 to 131320 => "11111111",
--		131461 to 131465 => "11111111",
--		131606 to 131610 => "11111111",
--		132195 to 132199 => "11111111",
--		132340 to 132344 => "11111111",
--		132485 to 132489 => "11111111",
--		132630 to 132634 => "11111111",
--		133219 to 133223 => "11111111",
--		133364 to 133368 => "11111111",
--		133509 to 133513 => "11111111",
--		133654 to 133658 => "11111111",
--		134243 to 134247 => "11111111",
--		134388 to 134392 => "11111111",
--		134533 to 134537 => "11111111",
--		134678 to 134682 => "11111111",
--		135267 to 135271 => "11111111",
--		135412 to 135416 => "11111111",
--		135557 to 135561 => "11111111",
--		135702 to 135706 => "11111111",
--		136291 to 136295 => "11111111",
--		136436 to 136440 => "11111111",
--		136581 to 136585 => "11111111",
--		136726 to 136730 => "11111111",
--		137315 to 137319 => "11111111",
--		137460 to 137464 => "11111111",
--		137605 to 137609 => "11111111",
--		137750 to 137754 => "11111111",
--		138339 to 138343 => "11111111",
--		138484 to 138488 => "11111111",
--		138629 to 138633 => "11111111",
--		138774 to 138778 => "11111111",
--		139363 to 139367 => "11111111",
--		139508 to 139512 => "11111111",
--		139653 to 139657 => "11111111",
--		139798 to 139802 => "11111111",
--		140387 to 140391 => "11111111",
--		140532 to 140536 => "11111111",
--		140677 to 140681 => "11111111",
--		140822 to 140826 => "11111111",
--		141411 to 141415 => "11111111",
--		141556 to 141560 => "11111111",
--		141701 to 141705 => "11111111",
--		141846 to 141850 => "11111111",
--		142435 to 142439 => "11111111",
--		142580 to 142584 => "11111111",
--		142725 to 142729 => "11111111",
--		142870 to 142874 => "11111111",
--		143459 to 143463 => "11111111",
--		143604 to 143608 => "11111111",
--		143749 to 143753 => "11111111",
--		143894 to 143898 => "11111111",
--		144483 to 144487 => "11111111",
--		144628 to 144632 => "11111111",
--		144773 to 144777 => "11111111",
--		144918 to 144922 => "11111111",
--		145507 to 145511 => "11111111",
--		145652 to 145656 => "11111111",
--		145797 to 145801 => "11111111",
--		145942 to 145946 => "11111111",
--		146531 to 146535 => "11111111",
--		146676 to 146680 => "11111111",
--		146821 to 146825 => "11111111",
--		146966 to 146970 => "11111111",
--		147555 to 147559 => "11111111",
--		147700 to 147704 => "11111111",
--		147845 to 147849 => "11111111",
--		147990 to 147994 => "11111111",
--		148579 to 148583 => "11111111",
--		148724 to 148728 => "11111111",
--		148869 to 148873 => "11111111",
--		149014 to 149018 => "11111111",
--		149603 to 149607 => "11111111",
--		149748 to 149752 => "11111111",
--		149893 to 149897 => "11111111",
--		150038 to 150042 => "11111111",
--		150627 to 150631 => "11111111",
--		150772 to 150776 => "11111111",
--		150917 to 150921 => "11111111",
--		151062 to 151066 => "11111111",
--		151651 to 151655 => "11111111",
--		151796 to 151800 => "11111111",
--		151941 to 151945 => "11111111",
--		152086 to 152090 => "11111111",
--		152675 to 152679 => "11111111",
--		152820 to 152824 => "11111111",
--		152965 to 152969 => "11111111",
--		153110 to 153114 => "11111111",
--		153699 to 153703 => "11111111",
--		153844 to 153848 => "11111111",
--		153989 to 153993 => "11111111",
--		154134 to 154138 => "11111111",
--		154723 to 154727 => "11111111",
--		154868 to 154872 => "11111111",
--		155013 to 155017 => "11111111",
--		155158 to 155162 => "11111111",
--		155747 to 155751 => "11111111",
--		155892 to 155896 => "11111111",
--		156037 to 156041 => "11111111",
--		156182 to 156186 => "11111111",
--		156771 to 156775 => "11111111",
--		156916 to 156920 => "11111111",
--		157061 to 157065 => "11111111",
--		157206 to 157210 => "11111111",
--		157795 to 157799 => "11111111",
--		157940 to 157944 => "11111111",
--		158085 to 158089 => "11111111",
--		158230 to 158234 => "11111111",
--		158819 to 158823 => "11111111",
--		158964 to 158968 => "11111111",
--		159109 to 159113 => "11111111",
--		159254 to 159258 => "11111111",
--		159843 to 159847 => "11111111",
--		159988 to 159992 => "11111111",
--		160133 to 160137 => "11111111",
--		160278 to 160282 => "11111111",
--		160867 to 160871 => "11111111",
--		161012 to 161016 => "11111111",
--		161157 to 161161 => "11111111",
--		161302 to 161306 => "11111111",
--		161891 to 161895 => "11111111",
--		162036 to 162040 => "11111111",
--		162181 to 162185 => "11111111",
--		162326 to 162330 => "11111111",
--		162915 to 162919 => "11111111",
--		163060 to 163064 => "11111111",
--		163205 to 163209 => "11111111",
--		163350 to 163354 => "11111111",
--		163939 to 163943 => "11111111",
--		164084 to 164088 => "11111111",
--		164229 to 164233 => "11111111",
--		164374 to 164378 => "11111111",
--		164963 to 164967 => "11111111",
--		165108 to 165112 => "11111111",
--		165253 to 165257 => "11111111",
--		165398 to 165402 => "11111111",
--		165987 to 165991 => "11111111",
--		166132 to 166136 => "11111111",
--		166277 to 166281 => "11111111",
--		166422 to 166426 => "11111111",
--		167011 to 167015 => "11111111",
--		167156 to 167160 => "11111111",
--		167301 to 167305 => "11111111",
--		167446 to 167450 => "11111111",
--		168035 to 168474 => "11111111",
--		169059 to 169498 => "11111111",
--		170083 to 170522 => "11111111",
--		171107 to 171546 => "11111111",
--		172131 to 172570 => "11111111",
--		173155 to 173159 => "11111111",
--		173300 to 173304 => "11111111",
--		173445 to 173449 => "11111111",
--		173590 to 173594 => "11111111",
--		174179 to 174183 => "11111111",
--		174324 to 174328 => "11111111",
--		174469 to 174473 => "11111111",
--		174614 to 174618 => "11111111",
--		175203 to 175207 => "11111111",
--		175348 to 175352 => "11111111",
--		175493 to 175497 => "11111111",
--		175638 to 175642 => "11111111",
--		176227 to 176231 => "11111111",
--		176372 to 176376 => "11111111",
--		176517 to 176521 => "11111111",
--		176662 to 176666 => "11111111",
--		177251 to 177255 => "11111111",
--		177396 to 177400 => "11111111",
--		177541 to 177545 => "11111111",
--		177686 to 177690 => "11111111",
--		178275 to 178279 => "11111111",
--		178420 to 178424 => "11111111",
--		178565 to 178569 => "11111111",
--		178710 to 178714 => "11111111",
--		179299 to 179303 => "11111111",
--		179444 to 179448 => "11111111",
--		179589 to 179593 => "11111111",
--		179734 to 179738 => "11111111",
--		180323 to 180327 => "11111111",
--		180468 to 180472 => "11111111",
--		180613 to 180617 => "11111111",
--		180758 to 180762 => "11111111",
--		181347 to 181351 => "11111111",
--		181492 to 181496 => "11111111",
--		181637 to 181641 => "11111111",
--		181782 to 181786 => "11111111",
--		182371 to 182375 => "11111111",
--		182516 to 182520 => "11111111",
--		182661 to 182665 => "11111111",
--		182806 to 182810 => "11111111",
--		183395 to 183399 => "11111111",
--		183540 to 183544 => "11111111",
--		183685 to 183689 => "11111111",
--		183830 to 183834 => "11111111",
--		184419 to 184423 => "11111111",
--		184564 to 184568 => "11111111",
--		184709 to 184713 => "11111111",
--		184854 to 184858 => "11111111",
--		185443 to 185447 => "11111111",
--		185588 to 185592 => "11111111",
--		185733 to 185737 => "11111111",
--		185878 to 185882 => "11111111",
--		186467 to 186471 => "11111111",
--		186612 to 186616 => "11111111",
--		186757 to 186761 => "11111111",
--		186902 to 186906 => "11111111",
--		187491 to 187495 => "11111111",
--		187636 to 187640 => "11111111",
--		187781 to 187785 => "11111111",
--		187926 to 187930 => "11111111",
--		188515 to 188519 => "11111111",
--		188660 to 188664 => "11111111",
--		188805 to 188809 => "11111111",
--		188950 to 188954 => "11111111",
--		189539 to 189543 => "11111111",
--		189684 to 189688 => "11111111",
--		189829 to 189833 => "11111111",
--		189974 to 189978 => "11111111",
--		190563 to 190567 => "11111111",
--		190708 to 190712 => "11111111",
--		190853 to 190857 => "11111111",
--		190998 to 191002 => "11111111",
--		191587 to 191591 => "11111111",
--		191732 to 191736 => "11111111",
--		191877 to 191881 => "11111111",
--		192022 to 192026 => "11111111",
--		192611 to 192615 => "11111111",
--		192756 to 192760 => "11111111",
--		192901 to 192905 => "11111111",
--		193046 to 193050 => "11111111",
--		193635 to 193639 => "11111111",
--		193780 to 193784 => "11111111",
--		193925 to 193929 => "11111111",
--		194070 to 194074 => "11111111",
--		194659 to 194663 => "11111111",
--		194804 to 194808 => "11111111",
--		194949 to 194953 => "11111111",
--		195094 to 195098 => "11111111",
--		195683 to 195687 => "11111111",
--		195828 to 195832 => "11111111",
--		195973 to 195977 => "11111111",
--		196118 to 196122 => "11111111",
--		196707 to 196711 => "11111111",
--		196852 to 196856 => "11111111",
--		196997 to 197001 => "11111111",
--		197142 to 197146 => "11111111",
--		197731 to 197735 => "11111111",
--		197876 to 197880 => "11111111",
--		198021 to 198025 => "11111111",
--		198166 to 198170 => "11111111",
--		198755 to 198759 => "11111111",
--		198900 to 198904 => "11111111",
--		199045 to 199049 => "11111111",
--		199190 to 199194 => "11111111",
--		199779 to 199783 => "11111111",
--		199924 to 199928 => "11111111",
--		200069 to 200073 => "11111111",
--		200214 to 200218 => "11111111",
--		200803 to 200807 => "11111111",
--		200948 to 200952 => "11111111",
--		201093 to 201097 => "11111111",
--		201238 to 201242 => "11111111",
--		201827 to 201831 => "11111111",
--		201972 to 201976 => "11111111",
--		202117 to 202121 => "11111111",
--		202262 to 202266 => "11111111",
--		202851 to 202855 => "11111111",
--		202996 to 203000 => "11111111",
--		203141 to 203145 => "11111111",
--		203286 to 203290 => "11111111",
--		203875 to 203879 => "11111111",
--		204020 to 204024 => "11111111",
--		204165 to 204169 => "11111111",
--		204310 to 204314 => "11111111",
--		204899 to 204903 => "11111111",
--		205044 to 205048 => "11111111",
--		205189 to 205193 => "11111111",
--		205334 to 205338 => "11111111",
--		205923 to 205927 => "11111111",
--		206068 to 206072 => "11111111",
--		206213 to 206217 => "11111111",
--		206358 to 206362 => "11111111",
--		206947 to 206951 => "11111111",
--		207092 to 207096 => "11111111",
--		207237 to 207241 => "11111111",
--		207382 to 207386 => "11111111",
--		207971 to 207975 => "11111111",
--		208116 to 208120 => "11111111",
--		208261 to 208265 => "11111111",
--		208406 to 208410 => "11111111",
--		208995 to 208999 => "11111111",
--		209140 to 209144 => "11111111",
--		209285 to 209289 => "11111111",
--		209430 to 209434 => "11111111",
--		210019 to 210023 => "11111111",
--		210164 to 210168 => "11111111",
--		210309 to 210313 => "11111111",
--		210454 to 210458 => "11111111",
--		211043 to 211047 => "11111111",
--		211188 to 211192 => "11111111",
--		211333 to 211337 => "11111111",
--		211478 to 211482 => "11111111",
--		212067 to 212071 => "11111111",
--		212212 to 212216 => "11111111",
--		212357 to 212361 => "11111111",
--		212502 to 212506 => "11111111",
--		213091 to 213095 => "11111111",
--		213236 to 213240 => "11111111",
--		213381 to 213385 => "11111111",
--		213526 to 213530 => "11111111",
--		214115 to 214119 => "11111111",
--		214260 to 214264 => "11111111",
--		214405 to 214409 => "11111111",
--		214550 to 214554 => "11111111",
--		215139 to 215143 => "11111111",
--		215284 to 215288 => "11111111",
--		215429 to 215433 => "11111111",
--		215574 to 215578 => "11111111",
--		216163 to 216167 => "11111111",
--		216308 to 216312 => "11111111",
--		216453 to 216457 => "11111111",
--		216598 to 216602 => "11111111",
--		217187 to 217191 => "11111111",
--		217332 to 217336 => "11111111",
--		217477 to 217481 => "11111111",
--		217622 to 217626 => "11111111",
--		218211 to 218215 => "11111111",
--		218356 to 218360 => "11111111",
--		218501 to 218505 => "11111111",
--		218646 to 218650 => "11111111",
--		219235 to 219239 => "11111111",
--		219380 to 219384 => "11111111",
--		219525 to 219529 => "11111111",
--		219670 to 219674 => "11111111",
--		220259 to 220263 => "11111111",
--		220404 to 220408 => "11111111",
--		220549 to 220553 => "11111111",
--		220694 to 220698 => "11111111",
--		221283 to 221287 => "11111111",
--		221428 to 221432 => "11111111",
--		221573 to 221577 => "11111111",
--		221718 to 221722 => "11111111",
--		222307 to 222311 => "11111111",
--		222452 to 222456 => "11111111",
--		222597 to 222601 => "11111111",
--		222742 to 222746 => "11111111",
--		223331 to 223335 => "11111111",
--		223476 to 223480 => "11111111",
--		223621 to 223625 => "11111111",
--		223766 to 223770 => "11111111",
--		224355 to 224359 => "11111111",
--		224500 to 224504 => "11111111",
--		224645 to 224649 => "11111111",
--		224790 to 224794 => "11111111",
--		225379 to 225383 => "11111111",
--		225524 to 225528 => "11111111",
--		225669 to 225673 => "11111111",
--		225814 to 225818 => "11111111",
--		226403 to 226407 => "11111111",
--		226548 to 226552 => "11111111",
--		226693 to 226697 => "11111111",
--		226838 to 226842 => "11111111",
--		227427 to 227431 => "11111111",
--		227572 to 227576 => "11111111",
--		227717 to 227721 => "11111111",
--		227862 to 227866 => "11111111",
--		228451 to 228455 => "11111111",
--		228596 to 228600 => "11111111",
--		228741 to 228745 => "11111111",
--		228886 to 228890 => "11111111",
--		229475 to 229479 => "11111111",
--		229620 to 229624 => "11111111",
--		229765 to 229769 => "11111111",
--		229910 to 229914 => "11111111",
--		230499 to 230503 => "11111111",
--		230644 to 230648 => "11111111",
--		230789 to 230793 => "11111111",
--		230934 to 230938 => "11111111",
--		231523 to 231527 => "11111111",
--		231668 to 231672 => "11111111",
--		231813 to 231817 => "11111111",
--		231958 to 231962 => "11111111",
--		232547 to 232551 => "11111111",
--		232692 to 232696 => "11111111",
--		232837 to 232841 => "11111111",
--		232982 to 232986 => "11111111",
--		233571 to 233575 => "11111111",
--		233716 to 233720 => "11111111",
--		233861 to 233865 => "11111111",
--		234006 to 234010 => "11111111",
--		234595 to 234599 => "11111111",
--		234740 to 234744 => "11111111",
--		234885 to 234889 => "11111111",
--		235030 to 235034 => "11111111",
--		235619 to 235623 => "11111111",
--		235764 to 235768 => "11111111",
--		235909 to 235913 => "11111111",
--		236054 to 236058 => "11111111",
--		236643 to 236647 => "11111111",
--		236788 to 236792 => "11111111",
--		236933 to 236937 => "11111111",
--		237078 to 237082 => "11111111",
--		237667 to 237671 => "11111111",
--		237812 to 237816 => "11111111",
--		237957 to 237961 => "11111111",
--		238102 to 238106 => "11111111",
--		238691 to 238695 => "11111111",
--		238836 to 238840 => "11111111",
--		238981 to 238985 => "11111111",
--		239126 to 239130 => "11111111",
--		239715 to 239719 => "11111111",
--		239860 to 239864 => "11111111",
--		240005 to 240009 => "11111111",
--		240150 to 240154 => "11111111",
--		240739 to 240743 => "11111111",
--		240884 to 240888 => "11111111",
--		241029 to 241033 => "11111111",
--		241174 to 241178 => "11111111",
--		241763 to 241767 => "11111111",
--		241908 to 241912 => "11111111",
--		242053 to 242057 => "11111111",
--		242198 to 242202 => "11111111",
--		242787 to 242791 => "11111111",
--		242932 to 242936 => "11111111",
--		243077 to 243081 => "11111111",
--		243222 to 243226 => "11111111",
--		243811 to 243815 => "11111111",
--		243956 to 243960 => "11111111",
--		244101 to 244105 => "11111111",
--		244246 to 244250 => "11111111",
--		244835 to 244839 => "11111111",
--		244980 to 244984 => "11111111",
--		245125 to 245129 => "11111111",
--		245270 to 245274 => "11111111",
--		245859 to 245863 => "11111111",
--		246004 to 246008 => "11111111",
--		246149 to 246153 => "11111111",
--		246294 to 246298 => "11111111",
--		246883 to 246887 => "11111111",
--		247028 to 247032 => "11111111",
--		247173 to 247177 => "11111111",
--		247318 to 247322 => "11111111",
--		247907 to 247911 => "11111111",
--		248052 to 248056 => "11111111",
--		248197 to 248201 => "11111111",
--		248342 to 248346 => "11111111",
--		248931 to 248935 => "11111111",
--		249076 to 249080 => "11111111",
--		249221 to 249225 => "11111111",
--		249366 to 249370 => "11111111",
--		249955 to 249959 => "11111111",
--		250100 to 250104 => "11111111",
--		250245 to 250249 => "11111111",
--		250390 to 250394 => "11111111",
--		250979 to 250983 => "11111111",
--		251124 to 251128 => "11111111",
--		251269 to 251273 => "11111111",
--		251414 to 251418 => "11111111",
--		252003 to 252007 => "11111111",
--		252148 to 252152 => "11111111",
--		252293 to 252297 => "11111111",
--		252438 to 252442 => "11111111",
--		253027 to 253031 => "11111111",
--		253172 to 253176 => "11111111",
--		253317 to 253321 => "11111111",
--		253462 to 253466 => "11111111",
--		254051 to 254055 => "11111111",
--		254196 to 254200 => "11111111",
--		254341 to 254345 => "11111111",
--		254486 to 254490 => "11111111",
--		255075 to 255079 => "11111111",
--		255220 to 255224 => "11111111",
--		255365 to 255369 => "11111111",
--		255510 to 255514 => "11111111",
--		256099 to 256103 => "11111111",
--		256244 to 256248 => "11111111",
--		256389 to 256393 => "11111111",
--		256534 to 256538 => "11111111",
--		257123 to 257127 => "11111111",
--		257268 to 257272 => "11111111",
--		257413 to 257417 => "11111111",
--		257558 to 257562 => "11111111",
--		258147 to 258151 => "11111111",
--		258292 to 258296 => "11111111",
--		258437 to 258441 => "11111111",
--		258582 to 258586 => "11111111",
--		259171 to 259175 => "11111111",
--		259316 to 259320 => "11111111",
--		259461 to 259465 => "11111111",
--		259606 to 259610 => "11111111",
--		260195 to 260199 => "11111111",
--		260340 to 260344 => "11111111",
--		260485 to 260489 => "11111111",
--		260630 to 260634 => "11111111",
--		261219 to 261223 => "11111111",
--		261364 to 261368 => "11111111",
--		261509 to 261513 => "11111111",
--		261654 to 261658 => "11111111",
--		262243 to 262247 => "11111111",
--		262388 to 262392 => "11111111",
--		262533 to 262537 => "11111111",
--		262678 to 262682 => "11111111",
--		263267 to 263271 => "11111111",
--		263412 to 263416 => "11111111",
--		263557 to 263561 => "11111111",
--		263702 to 263706 => "11111111",
--		264291 to 264295 => "11111111",
--		264436 to 264440 => "11111111",
--		264581 to 264585 => "11111111",
--		264726 to 264730 => "11111111",
--		265315 to 265319 => "11111111",
--		265460 to 265464 => "11111111",
--		265605 to 265609 => "11111111",
--		265750 to 265754 => "11111111",
--		266339 to 266343 => "11111111",
--		266484 to 266488 => "11111111",
--		266629 to 266633 => "11111111",
--		266774 to 266778 => "11111111",
--		267363 to 267367 => "11111111",
--		267508 to 267512 => "11111111",
--		267653 to 267657 => "11111111",
--		267798 to 267802 => "11111111",
--		268387 to 268391 => "11111111",
--		268532 to 268536 => "11111111",
--		268677 to 268681 => "11111111",
--		268822 to 268826 => "11111111",
--		269411 to 269415 => "11111111",
--		269556 to 269560 => "11111111",
--		269701 to 269705 => "11111111",
--		269846 to 269850 => "11111111",
--		270435 to 270439 => "11111111",
--		270580 to 270584 => "11111111",
--		270725 to 270729 => "11111111",
--		270870 to 270874 => "11111111",
--		271459 to 271463 => "11111111",
--		271604 to 271608 => "11111111",
--		271749 to 271753 => "11111111",
--		271894 to 271898 => "11111111",
--		272483 to 272487 => "11111111",
--		272628 to 272632 => "11111111",
--		272773 to 272777 => "11111111",
--		272918 to 272922 => "11111111",
--		273507 to 273511 => "11111111",
--		273652 to 273656 => "11111111",
--		273797 to 273801 => "11111111",
--		273942 to 273946 => "11111111",
--		274531 to 274535 => "11111111",
--		274676 to 274680 => "11111111",
--		274821 to 274825 => "11111111",
--		274966 to 274970 => "11111111",
--		275555 to 275559 => "11111111",
--		275700 to 275704 => "11111111",
--		275845 to 275849 => "11111111",
--		275990 to 275994 => "11111111",
--		276579 to 276583 => "11111111",
--		276724 to 276728 => "11111111",
--		276869 to 276873 => "11111111",
--		277014 to 277018 => "11111111",
--		277603 to 277607 => "11111111",
--		277748 to 277752 => "11111111",
--		277893 to 277897 => "11111111",
--		278038 to 278042 => "11111111",
--		278627 to 278631 => "11111111",
--		278772 to 278776 => "11111111",
--		278917 to 278921 => "11111111",
--		279062 to 279066 => "11111111",
--		279651 to 279655 => "11111111",
--		279796 to 279800 => "11111111",
--		279941 to 279945 => "11111111",
--		280086 to 280090 => "11111111",
--		280675 to 280679 => "11111111",
--		280820 to 280824 => "11111111",
--		280965 to 280969 => "11111111",
--		281110 to 281114 => "11111111",
--		281699 to 281703 => "11111111",
--		281844 to 281848 => "11111111",
--		281989 to 281993 => "11111111",
--		282134 to 282138 => "11111111",
--		282723 to 282727 => "11111111",
--		282868 to 282872 => "11111111",
--		283013 to 283017 => "11111111",
--		283158 to 283162 => "11111111",
--		283747 to 283751 => "11111111",
--		283892 to 283896 => "11111111",
--		284037 to 284041 => "11111111",
--		284182 to 284186 => "11111111",
--		284771 to 284775 => "11111111",
--		284916 to 284920 => "11111111",
--		285061 to 285065 => "11111111",
--		285206 to 285210 => "11111111",
--		285795 to 285799 => "11111111",
--		285940 to 285944 => "11111111",
--		286085 to 286089 => "11111111",
--		286230 to 286234 => "11111111",
--		286819 to 286823 => "11111111",
--		286964 to 286968 => "11111111",
--		287109 to 287113 => "11111111",
--		287254 to 287258 => "11111111",
--		287843 to 287847 => "11111111",
--		287988 to 287992 => "11111111",
--		288133 to 288137 => "11111111",
--		288278 to 288282 => "11111111",
--		288867 to 288871 => "11111111",
--		289012 to 289016 => "11111111",
--		289157 to 289161 => "11111111",
--		289302 to 289306 => "11111111",
--		289891 to 289895 => "11111111",
--		290036 to 290040 => "11111111",
--		290181 to 290185 => "11111111",
--		290326 to 290330 => "11111111",
--		290915 to 290919 => "11111111",
--		291060 to 291064 => "11111111",
--		291205 to 291209 => "11111111",
--		291350 to 291354 => "11111111",
--		291939 to 291943 => "11111111",
--		292084 to 292088 => "11111111",
--		292229 to 292233 => "11111111",
--		292374 to 292378 => "11111111",
--		292963 to 292967 => "11111111",
--		293108 to 293112 => "11111111",
--		293253 to 293257 => "11111111",
--		293398 to 293402 => "11111111",
--		293987 to 293991 => "11111111",
--		294132 to 294136 => "11111111",
--		294277 to 294281 => "11111111",
--		294422 to 294426 => "11111111",
--		295011 to 295015 => "11111111",
--		295156 to 295160 => "11111111",
--		295301 to 295305 => "11111111",
--		295446 to 295450 => "11111111",
--		296035 to 296039 => "11111111",
--		296180 to 296184 => "11111111",
--		296325 to 296329 => "11111111",
--		296470 to 296474 => "11111111",
--		297059 to 297063 => "11111111",
--		297204 to 297208 => "11111111",
--		297349 to 297353 => "11111111",
--		297494 to 297498 => "11111111",
--		298083 to 298087 => "11111111",
--		298228 to 298232 => "11111111",
--		298373 to 298377 => "11111111",
--		298518 to 298522 => "11111111",
--		299107 to 299111 => "11111111",
--		299252 to 299256 => "11111111",
--		299397 to 299401 => "11111111",
--		299542 to 299546 => "11111111",
--		300131 to 300135 => "11111111",
--		300276 to 300280 => "11111111",
--		300421 to 300425 => "11111111",
--		300566 to 300570 => "11111111",
--		301155 to 301159 => "11111111",
--		301300 to 301304 => "11111111",
--		301445 to 301449 => "11111111",
--		301590 to 301594 => "11111111",
--		302179 to 302183 => "11111111",
--		302324 to 302328 => "11111111",
--		302469 to 302473 => "11111111",
--		302614 to 302618 => "11111111",
--		303203 to 303207 => "11111111",
--		303348 to 303352 => "11111111",
--		303493 to 303497 => "11111111",
--		303638 to 303642 => "11111111",
--		304227 to 304231 => "11111111",
--		304372 to 304376 => "11111111",
--		304517 to 304521 => "11111111",
--		304662 to 304666 => "11111111",
--		305251 to 305255 => "11111111",
--		305396 to 305400 => "11111111",
--		305541 to 305545 => "11111111",
--		305686 to 305690 => "11111111",
--		306275 to 306279 => "11111111",
--		306420 to 306424 => "11111111",
--		306565 to 306569 => "11111111",
--		306710 to 306714 => "11111111",
--		307299 to 307303 => "11111111",
--		307444 to 307448 => "11111111",
--		307589 to 307593 => "11111111",
--		307734 to 307738 => "11111111",
--		308323 to 308327 => "11111111",
--		308468 to 308472 => "11111111",
--		308613 to 308617 => "11111111",
--		308758 to 308762 => "11111111",
--		309347 to 309351 => "11111111",
--		309492 to 309496 => "11111111",
--		309637 to 309641 => "11111111",
--		309782 to 309786 => "11111111",
--		310371 to 310375 => "11111111",
--		310516 to 310520 => "11111111",
--		310661 to 310665 => "11111111",
--		310806 to 310810 => "11111111",
--		311395 to 311399 => "11111111",
--		311540 to 311544 => "11111111",
--		311685 to 311689 => "11111111",
--		311830 to 311834 => "11111111",
--		312419 to 312423 => "11111111",
--		312564 to 312568 => "11111111",
--		312709 to 312713 => "11111111",
--		312854 to 312858 => "11111111",
--		313443 to 313447 => "11111111",
--		313588 to 313592 => "11111111",
--		313733 to 313737 => "11111111",
--		313878 to 313882 => "11111111",
--		314467 to 314471 => "11111111",
--		314612 to 314616 => "11111111",
--		314757 to 314761 => "11111111",
--		314902 to 314906 => "11111111",
--		315491 to 315495 => "11111111",
--		315636 to 315640 => "11111111",
--		315781 to 315785 => "11111111",
--		315926 to 315930 => "11111111",
--		316515 to 316954 => "11111111",
--		317539 to 317978 => "11111111",
--		318563 to 319002 => "11111111",
--		319587 to 320026 => "11111111",
--		320611 to 321050 => "11111111",
--		321635 to 321639 => "11111111",
--		321780 to 321784 => "11111111",
--		321925 to 321929 => "11111111",
--		322070 to 322074 => "11111111",
--		322659 to 322663 => "11111111",
--		322804 to 322808 => "11111111",
--		322949 to 322953 => "11111111",
--		323094 to 323098 => "11111111",
--		323683 to 323687 => "11111111",
--		323828 to 323832 => "11111111",
--		323973 to 323977 => "11111111",
--		324118 to 324122 => "11111111",
--		324707 to 324711 => "11111111",
--		324852 to 324856 => "11111111",
--		324997 to 325001 => "11111111",
--		325142 to 325146 => "11111111",
--		325731 to 325735 => "11111111",
--		325876 to 325880 => "11111111",
--		326021 to 326025 => "11111111",
--		326166 to 326170 => "11111111",
--		326755 to 326759 => "11111111",
--		326900 to 326904 => "11111111",
--		327045 to 327049 => "11111111",
--		327190 to 327194 => "11111111",
--		327779 to 327783 => "11111111",
--		327924 to 327928 => "11111111",
--		328069 to 328073 => "11111111",
--		328214 to 328218 => "11111111",
--		328803 to 328807 => "11111111",
--		328948 to 328952 => "11111111",
--		329093 to 329097 => "11111111",
--		329238 to 329242 => "11111111",
--		329827 to 329831 => "11111111",
--		329972 to 329976 => "11111111",
--		330117 to 330121 => "11111111",
--		330262 to 330266 => "11111111",
--		330851 to 330855 => "11111111",
--		330996 to 331000 => "11111111",
--		331141 to 331145 => "11111111",
--		331286 to 331290 => "11111111",
--		331875 to 331879 => "11111111",
--		332020 to 332024 => "11111111",
--		332165 to 332169 => "11111111",
--		332310 to 332314 => "11111111",
--		332899 to 332903 => "11111111",
--		333044 to 333048 => "11111111",
--		333189 to 333193 => "11111111",
--		333334 to 333338 => "11111111",
--		333923 to 333927 => "11111111",
--		334068 to 334072 => "11111111",
--		334213 to 334217 => "11111111",
--		334358 to 334362 => "11111111",
--		334947 to 334951 => "11111111",
--		335092 to 335096 => "11111111",
--		335237 to 335241 => "11111111",
--		335382 to 335386 => "11111111",
--		335971 to 335975 => "11111111",
--		336116 to 336120 => "11111111",
--		336261 to 336265 => "11111111",
--		336406 to 336410 => "11111111",
--		336995 to 336999 => "11111111",
--		337140 to 337144 => "11111111",
--		337285 to 337289 => "11111111",
--		337430 to 337434 => "11111111",
--		338019 to 338023 => "11111111",
--		338164 to 338168 => "11111111",
--		338309 to 338313 => "11111111",
--		338454 to 338458 => "11111111",
--		339043 to 339047 => "11111111",
--		339188 to 339192 => "11111111",
--		339333 to 339337 => "11111111",
--		339478 to 339482 => "11111111",
--		340067 to 340071 => "11111111",
--		340212 to 340216 => "11111111",
--		340357 to 340361 => "11111111",
--		340502 to 340506 => "11111111",
--		341091 to 341095 => "11111111",
--		341236 to 341240 => "11111111",
--		341381 to 341385 => "11111111",
--		341526 to 341530 => "11111111",
--		342115 to 342119 => "11111111",
--		342260 to 342264 => "11111111",
--		342405 to 342409 => "11111111",
--		342550 to 342554 => "11111111",
--		343139 to 343143 => "11111111",
--		343284 to 343288 => "11111111",
--		343429 to 343433 => "11111111",
--		343574 to 343578 => "11111111",
--		344163 to 344167 => "11111111",
--		344308 to 344312 => "11111111",
--		344453 to 344457 => "11111111",
--		344598 to 344602 => "11111111",
--		345187 to 345191 => "11111111",
--		345332 to 345336 => "11111111",
--		345477 to 345481 => "11111111",
--		345622 to 345626 => "11111111",
--		346211 to 346215 => "11111111",
--		346356 to 346360 => "11111111",
--		346501 to 346505 => "11111111",
--		346646 to 346650 => "11111111",
--		347235 to 347239 => "11111111",
--		347380 to 347384 => "11111111",
--		347525 to 347529 => "11111111",
--		347670 to 347674 => "11111111",
--		348259 to 348263 => "11111111",
--		348404 to 348408 => "11111111",
--		348549 to 348553 => "11111111",
--		348694 to 348698 => "11111111",
--		349283 to 349287 => "11111111",
--		349428 to 349432 => "11111111",
--		349573 to 349577 => "11111111",
--		349718 to 349722 => "11111111",
--		350307 to 350311 => "11111111",
--		350452 to 350456 => "11111111",
--		350597 to 350601 => "11111111",
--		350742 to 350746 => "11111111",
--		351331 to 351335 => "11111111",
--		351476 to 351480 => "11111111",
--		351621 to 351625 => "11111111",
--		351766 to 351770 => "11111111",
--		352355 to 352359 => "11111111",
--		352500 to 352504 => "11111111",
--		352645 to 352649 => "11111111",
--		352790 to 352794 => "11111111",
--		353379 to 353383 => "11111111",
--		353524 to 353528 => "11111111",
--		353669 to 353673 => "11111111",
--		353814 to 353818 => "11111111",
--		354403 to 354407 => "11111111",
--		354548 to 354552 => "11111111",
--		354693 to 354697 => "11111111",
--		354838 to 354842 => "11111111",
--		355427 to 355431 => "11111111",
--		355572 to 355576 => "11111111",
--		355717 to 355721 => "11111111",
--		355862 to 355866 => "11111111",
--		356451 to 356455 => "11111111",
--		356596 to 356600 => "11111111",
--		356741 to 356745 => "11111111",
--		356886 to 356890 => "11111111",
--		357475 to 357479 => "11111111",
--		357620 to 357624 => "11111111",
--		357765 to 357769 => "11111111",
--		357910 to 357914 => "11111111",
--		358499 to 358503 => "11111111",
--		358644 to 358648 => "11111111",
--		358789 to 358793 => "11111111",
--		358934 to 358938 => "11111111",
--		359523 to 359527 => "11111111",
--		359668 to 359672 => "11111111",
--		359813 to 359817 => "11111111",
--		359958 to 359962 => "11111111",
--		360547 to 360551 => "11111111",
--		360692 to 360696 => "11111111",
--		360837 to 360841 => "11111111",
--		360982 to 360986 => "11111111",
--		361571 to 361575 => "11111111",
--		361716 to 361720 => "11111111",
--		361861 to 361865 => "11111111",
--		362006 to 362010 => "11111111",
--		362595 to 362599 => "11111111",
--		362740 to 362744 => "11111111",
--		362885 to 362889 => "11111111",
--		363030 to 363034 => "11111111",
--		363619 to 363623 => "11111111",
--		363764 to 363768 => "11111111",
--		363909 to 363913 => "11111111",
--		364054 to 364058 => "11111111",
--		364643 to 364647 => "11111111",
--		364788 to 364792 => "11111111",
--		364933 to 364937 => "11111111",
--		365078 to 365082 => "11111111",
--		365667 to 365671 => "11111111",
--		365812 to 365816 => "11111111",
--		365957 to 365961 => "11111111",
--		366102 to 366106 => "11111111",
--		366691 to 366695 => "11111111",
--		366836 to 366840 => "11111111",
--		366981 to 366985 => "11111111",
--		367126 to 367130 => "11111111",
--		367715 to 367719 => "11111111",
--		367860 to 367864 => "11111111",
--		368005 to 368009 => "11111111",
--		368150 to 368154 => "11111111",
--		368739 to 368743 => "11111111",
--		368884 to 368888 => "11111111",
--		369029 to 369033 => "11111111",
--		369174 to 369178 => "11111111",
--		369763 to 369767 => "11111111",
--		369908 to 369912 => "11111111",
--		370053 to 370057 => "11111111",
--		370198 to 370202 => "11111111",
--		370787 to 370791 => "11111111",
--		370932 to 370936 => "11111111",
--		371077 to 371081 => "11111111",
--		371222 to 371226 => "11111111",
--		371811 to 371815 => "11111111",
--		371956 to 371960 => "11111111",
--		372101 to 372105 => "11111111",
--		372246 to 372250 => "11111111",
--		372835 to 372839 => "11111111",
--		372980 to 372984 => "11111111",
--		373125 to 373129 => "11111111",
--		373270 to 373274 => "11111111",
--		373859 to 373863 => "11111111",
--		374004 to 374008 => "11111111",
--		374149 to 374153 => "11111111",
--		374294 to 374298 => "11111111",
--		374883 to 374887 => "11111111",
--		375028 to 375032 => "11111111",
--		375173 to 375177 => "11111111",
--		375318 to 375322 => "11111111",
--		375907 to 375911 => "11111111",
--		376052 to 376056 => "11111111",
--		376197 to 376201 => "11111111",
--		376342 to 376346 => "11111111",
--		376931 to 376935 => "11111111",
--		377076 to 377080 => "11111111",
--		377221 to 377225 => "11111111",
--		377366 to 377370 => "11111111",
--		377955 to 377959 => "11111111",
--		378100 to 378104 => "11111111",
--		378245 to 378249 => "11111111",
--		378390 to 378394 => "11111111",
--		378979 to 378983 => "11111111",
--		379124 to 379128 => "11111111",
--		379269 to 379273 => "11111111",
--		379414 to 379418 => "11111111",
--		380003 to 380007 => "11111111",
--		380148 to 380152 => "11111111",
--		380293 to 380297 => "11111111",
--		380438 to 380442 => "11111111",
--		381027 to 381031 => "11111111",
--		381172 to 381176 => "11111111",
--		381317 to 381321 => "11111111",
--		381462 to 381466 => "11111111",
--		382051 to 382055 => "11111111",
--		382196 to 382200 => "11111111",
--		382341 to 382345 => "11111111",
--		382486 to 382490 => "11111111",
--		383075 to 383079 => "11111111",
--		383220 to 383224 => "11111111",
--		383365 to 383369 => "11111111",
--		383510 to 383514 => "11111111",
--		384099 to 384103 => "11111111",
--		384244 to 384248 => "11111111",
--		384389 to 384393 => "11111111",
--		384534 to 384538 => "11111111",
--		385123 to 385127 => "11111111",
--		385268 to 385272 => "11111111",
--		385413 to 385417 => "11111111",
--		385558 to 385562 => "11111111",
--		386147 to 386151 => "11111111",
--		386292 to 386296 => "11111111",
--		386437 to 386441 => "11111111",
--		386582 to 386586 => "11111111",
--		387171 to 387175 => "11111111",
--		387316 to 387320 => "11111111",
--		387461 to 387465 => "11111111",
--		387606 to 387610 => "11111111",
--		388195 to 388199 => "11111111",
--		388340 to 388344 => "11111111",
--		388485 to 388489 => "11111111",
--		388630 to 388634 => "11111111",
--		389219 to 389223 => "11111111",
--		389364 to 389368 => "11111111",
--		389509 to 389513 => "11111111",
--		389654 to 389658 => "11111111",
--		390243 to 390247 => "11111111",
--		390388 to 390392 => "11111111",
--		390533 to 390537 => "11111111",
--		390678 to 390682 => "11111111",
--		391267 to 391271 => "11111111",
--		391412 to 391416 => "11111111",
--		391557 to 391561 => "11111111",
--		391702 to 391706 => "11111111",
--		392291 to 392295 => "11111111",
--		392436 to 392440 => "11111111",
--		392581 to 392585 => "11111111",
--		392726 to 392730 => "11111111",
--		393315 to 393319 => "11111111",
--		393460 to 393464 => "11111111",
--		393605 to 393609 => "11111111",
--		393750 to 393754 => "11111111",
--		394339 to 394343 => "11111111",
--		394484 to 394488 => "11111111",
--		394629 to 394633 => "11111111",
--		394774 to 394778 => "11111111",
--		395363 to 395367 => "11111111",
--		395508 to 395512 => "11111111",
--		395653 to 395657 => "11111111",
--		395798 to 395802 => "11111111",
--		396387 to 396391 => "11111111",
--		396532 to 396536 => "11111111",
--		396677 to 396681 => "11111111",
--		396822 to 396826 => "11111111",
--		397411 to 397415 => "11111111",
--		397556 to 397560 => "11111111",
--		397701 to 397705 => "11111111",
--		397846 to 397850 => "11111111",
--		398435 to 398439 => "11111111",
--		398580 to 398584 => "11111111",
--		398725 to 398729 => "11111111",
--		398870 to 398874 => "11111111",
--		399459 to 399463 => "11111111",
--		399604 to 399608 => "11111111",
--		399749 to 399753 => "11111111",
--		399894 to 399898 => "11111111",
--		400483 to 400487 => "11111111",
--		400628 to 400632 => "11111111",
--		400773 to 400777 => "11111111",
--		400918 to 400922 => "11111111",
--		401507 to 401511 => "11111111",
--		401652 to 401656 => "11111111",
--		401797 to 401801 => "11111111",
--		401942 to 401946 => "11111111",
--		402531 to 402535 => "11111111",
--		402676 to 402680 => "11111111",
--		402821 to 402825 => "11111111",
--		402966 to 402970 => "11111111",
--		403555 to 403559 => "11111111",
--		403700 to 403704 => "11111111",
--		403845 to 403849 => "11111111",
--		403990 to 403994 => "11111111",
--		404579 to 404583 => "11111111",
--		404724 to 404728 => "11111111",
--		404869 to 404873 => "11111111",
--		405014 to 405018 => "11111111",
--		405603 to 405607 => "11111111",
--		405748 to 405752 => "11111111",
--		405893 to 405897 => "11111111",
--		406038 to 406042 => "11111111",
--		406627 to 406631 => "11111111",
--		406772 to 406776 => "11111111",
--		406917 to 406921 => "11111111",
--		407062 to 407066 => "11111111",
--		407651 to 407655 => "11111111",
--		407796 to 407800 => "11111111",
--		407941 to 407945 => "11111111",
--		408086 to 408090 => "11111111",
--		408675 to 408679 => "11111111",
--		408820 to 408824 => "11111111",
--		408965 to 408969 => "11111111",
--		409110 to 409114 => "11111111",
--		409699 to 409703 => "11111111",
--		409844 to 409848 => "11111111",
--		409989 to 409993 => "11111111",
--		410134 to 410138 => "11111111",
--		410723 to 410727 => "11111111",
--		410868 to 410872 => "11111111",
--		411013 to 411017 => "11111111",
--		411158 to 411162 => "11111111",
--		411747 to 411751 => "11111111",
--		411892 to 411896 => "11111111",
--		412037 to 412041 => "11111111",
--		412182 to 412186 => "11111111",
--		412771 to 412775 => "11111111",
--		412916 to 412920 => "11111111",
--		413061 to 413065 => "11111111",
--		413206 to 413210 => "11111111",
--		413795 to 413799 => "11111111",
--		413940 to 413944 => "11111111",
--		414085 to 414089 => "11111111",
--		414230 to 414234 => "11111111",
--		414819 to 414823 => "11111111",
--		414964 to 414968 => "11111111",
--		415109 to 415113 => "11111111",
--		415254 to 415258 => "11111111",
--		415843 to 415847 => "11111111",
--		415988 to 415992 => "11111111",
--		416133 to 416137 => "11111111",
--		416278 to 416282 => "11111111",
--		416867 to 416871 => "11111111",
--		417012 to 417016 => "11111111",
--		417157 to 417161 => "11111111",
--		417302 to 417306 => "11111111",
--		417891 to 417895 => "11111111",
--		418036 to 418040 => "11111111",
--		418181 to 418185 => "11111111",
--		418326 to 418330 => "11111111",
--		418915 to 418919 => "11111111",
--		419060 to 419064 => "11111111",
--		419205 to 419209 => "11111111",
--		419350 to 419354 => "11111111",
--		419939 to 419943 => "11111111",
--		420084 to 420088 => "11111111",
--		420229 to 420233 => "11111111",
--		420374 to 420378 => "11111111",
--		420963 to 420967 => "11111111",
--		421108 to 421112 => "11111111",
--		421253 to 421257 => "11111111",
--		421398 to 421402 => "11111111",
--		421987 to 421991 => "11111111",
--		422132 to 422136 => "11111111",
--		422277 to 422281 => "11111111",
--		422422 to 422426 => "11111111",
--		423011 to 423015 => "11111111",
--		423156 to 423160 => "11111111",
--		423301 to 423305 => "11111111",
--		423446 to 423450 => "11111111",
--		424035 to 424039 => "11111111",
--		424180 to 424184 => "11111111",
--		424325 to 424329 => "11111111",
--		424470 to 424474 => "11111111",
--		425059 to 425063 => "11111111",
--		425204 to 425208 => "11111111",
--		425349 to 425353 => "11111111",
--		425494 to 425498 => "11111111",
--		426083 to 426087 => "11111111",
--		426228 to 426232 => "11111111",
--		426373 to 426377 => "11111111",
--		426518 to 426522 => "11111111",
--		427107 to 427111 => "11111111",
--		427252 to 427256 => "11111111",
--		427397 to 427401 => "11111111",
--		427542 to 427546 => "11111111",
--		428131 to 428135 => "11111111",
--		428276 to 428280 => "11111111",
--		428421 to 428425 => "11111111",
--		428566 to 428570 => "11111111",
--		429155 to 429159 => "11111111",
--		429300 to 429304 => "11111111",
--		429445 to 429449 => "11111111",
--		429590 to 429594 => "11111111",
--		430179 to 430183 => "11111111",
--		430324 to 430328 => "11111111",
--		430469 to 430473 => "11111111",
--		430614 to 430618 => "11111111",
--		431203 to 431207 => "11111111",
--		431348 to 431352 => "11111111",
--		431493 to 431497 => "11111111",
--		431638 to 431642 => "11111111",
--		432227 to 432231 => "11111111",
--		432372 to 432376 => "11111111",
--		432517 to 432521 => "11111111",
--		432662 to 432666 => "11111111",
--		433251 to 433255 => "11111111",
--		433396 to 433400 => "11111111",
--		433541 to 433545 => "11111111",
--		433686 to 433690 => "11111111",
--		434275 to 434279 => "11111111",
--		434420 to 434424 => "11111111",
--		434565 to 434569 => "11111111",
--		434710 to 434714 => "11111111",
--		435299 to 435303 => "11111111",
--		435444 to 435448 => "11111111",
--		435589 to 435593 => "11111111",
--		435734 to 435738 => "11111111",
--		436323 to 436327 => "11111111",
--		436468 to 436472 => "11111111",
--		436613 to 436617 => "11111111",
--		436758 to 436762 => "11111111",
--		437347 to 437351 => "11111111",
--		437492 to 437496 => "11111111",
--		437637 to 437641 => "11111111",
--		437782 to 437786 => "11111111",
--		438371 to 438375 => "11111111",
--		438516 to 438520 => "11111111",
--		438661 to 438665 => "11111111",
--		438806 to 438810 => "11111111",
--		439395 to 439399 => "11111111",
--		439540 to 439544 => "11111111",
--		439685 to 439689 => "11111111",
--		439830 to 439834 => "11111111",
--		440419 to 440423 => "11111111",
--		440564 to 440568 => "11111111",
--		440709 to 440713 => "11111111",
--		440854 to 440858 => "11111111",
--		441443 to 441447 => "11111111",
--		441588 to 441592 => "11111111",
--		441733 to 441737 => "11111111",
--		441878 to 441882 => "11111111",
--		442467 to 442471 => "11111111",
--		442612 to 442616 => "11111111",
--		442757 to 442761 => "11111111",
--		442902 to 442906 => "11111111",
--		443491 to 443495 => "11111111",
--		443636 to 443640 => "11111111",
--		443781 to 443785 => "11111111",
--		443926 to 443930 => "11111111",
--		444515 to 444519 => "11111111",
--		444660 to 444664 => "11111111",
--		444805 to 444809 => "11111111",
--		444950 to 444954 => "11111111",
--		445539 to 445543 => "11111111",
--		445684 to 445688 => "11111111",
--		445829 to 445833 => "11111111",
--		445974 to 445978 => "11111111",
--		446563 to 446567 => "11111111",
--		446708 to 446712 => "11111111",
--		446853 to 446857 => "11111111",
--		446998 to 447002 => "11111111",
--		447587 to 447591 => "11111111",
--		447732 to 447736 => "11111111",
--		447877 to 447881 => "11111111",
--		448022 to 448026 => "11111111",
--		448611 to 448615 => "11111111",
--		448756 to 448760 => "11111111",
--		448901 to 448905 => "11111111",
--		449046 to 449050 => "11111111",
--		449635 to 449639 => "11111111",
--		449780 to 449784 => "11111111",
--		449925 to 449929 => "11111111",
--		450070 to 450074 => "11111111",
--		450659 to 450663 => "11111111",
--		450804 to 450808 => "11111111",
--		450949 to 450953 => "11111111",
--		451094 to 451098 => "11111111",
--		451683 to 451687 => "11111111",
--		451828 to 451832 => "11111111",
--		451973 to 451977 => "11111111",
--		452118 to 452122 => "11111111",
--		452707 to 452711 => "11111111",
--		452852 to 452856 => "11111111",
--		452997 to 453001 => "11111111",
--		453142 to 453146 => "11111111",
--		453731 to 453735 => "11111111",
--		453876 to 453880 => "11111111",
--		454021 to 454025 => "11111111",
--		454166 to 454170 => "11111111",
--		454755 to 454759 => "11111111",
--		454900 to 454904 => "11111111",
--		455045 to 455049 => "11111111",
--		455190 to 455194 => "11111111",
--		455779 to 455783 => "11111111",
--		455924 to 455928 => "11111111",
--		456069 to 456073 => "11111111",
--		456214 to 456218 => "11111111",
--		456803 to 456807 => "11111111",
--		456948 to 456952 => "11111111",
--		457093 to 457097 => "11111111",
--		457238 to 457242 => "11111111",
--		457827 to 457831 => "11111111",
--		457972 to 457976 => "11111111",
--		458117 to 458121 => "11111111",
--		458262 to 458266 => "11111111",
--		458851 to 458855 => "11111111",
--		458996 to 459000 => "11111111",
--		459141 to 459145 => "11111111",
--		459286 to 459290 => "11111111",
--		459875 to 459879 => "11111111",
--		460020 to 460024 => "11111111",
--		460165 to 460169 => "11111111",
--		460310 to 460314 => "11111111",
--		460899 to 460903 => "11111111",
--		461044 to 461048 => "11111111",
--		461189 to 461193 => "11111111",
--		461334 to 461338 => "11111111",
--		461923 to 461927 => "11111111",
--		462068 to 462072 => "11111111",
--		462213 to 462217 => "11111111",
--		462358 to 462362 => "11111111",
--		462947 to 462951 => "11111111",
--		463092 to 463096 => "11111111",
--		463237 to 463241 => "11111111",
--		463382 to 463386 => "11111111",
--		463971 to 463975 => "11111111",
--		464116 to 464120 => "11111111",
--		464261 to 464265 => "11111111",
--		464406 to 464410 => "11111111",
--		464995 to 465434 => "11111111",
--		466019 to 466458 => "11111111",
--		467043 to 467482 => "11111111",
--		468067 to 468506 => "11111111",
--		469091 to 469530 => "11111111",
		others=> "00000000");
begin

	process (Clk)
	begin
		if (Clk'event and Clk = '1') then
			if (CE = '1') then
				if (Enable_w = '1') then
					VRAM (to_integer(unsigned(Addr_w))) <= Data_in;
				end if;
				Data_out <= VRAM(to_integer(unsigned(Addr_r)));
			else
				NULL;
			end if;
		end if;
	end process;

end Behavioral;

					
