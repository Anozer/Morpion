		4140 to 4369 => "11111111",
		5164 to 5393 => "11111111",
		6188 to 6417 => "11111111",
		7212 to 7441 => "11111111",
		8236 to 8465 => "11111111",
		9260 to 9264 => "11111111",
		9335 to 9339 => "11111111",
		9410 to 9414 => "11111111",
		9485 to 9489 => "11111111",
		10284 to 10288 => "11111111",
		10359 to 10363 => "11111111",
		10434 to 10438 => "11111111",
		10509 to 10513 => "11111111",
		11308 to 11312 => "11111111",
		11383 to 11387 => "11111111",
		11458 to 11462 => "11111111",
		11533 to 11537 => "11111111",
		12332 to 12336 => "11111111",
		12407 to 12411 => "11111111",
		12482 to 12486 => "11111111",
		12557 to 12561 => "11111111",
		13356 to 13360 => "11111111",
		13431 to 13435 => "11111111",
		13506 to 13510 => "11111111",
		13581 to 13585 => "11111111",
		14380 to 14384 => "11111111",
		14455 to 14459 => "11111111",
		14530 to 14534 => "11111111",
		14605 to 14609 => "11111111",
		15404 to 15408 => "11111111",
		15479 to 15483 => "11111111",
		15554 to 15558 => "11111111",
		15629 to 15633 => "11111111",
		16428 to 16432 => "11111111",
		16503 to 16507 => "11111111",
		16578 to 16582 => "11111111",
		16653 to 16657 => "11111111",
		17452 to 17456 => "11111111",
		17527 to 17531 => "11111111",
		17602 to 17606 => "11111111",
		17677 to 17681 => "11111111",
		18476 to 18480 => "11111111",
		18551 to 18555 => "11111111",
		18626 to 18630 => "11111111",
		18701 to 18705 => "11111111",
		19500 to 19504 => "11111111",
		19575 to 19579 => "11111111",
		19650 to 19654 => "11111111",
		19725 to 19729 => "11111111",
		20524 to 20528 => "11111111",
		20599 to 20603 => "11111111",
		20674 to 20678 => "11111111",
		20749 to 20753 => "11111111",
		21548 to 21552 => "11111111",
		21623 to 21627 => "11111111",
		21698 to 21702 => "11111111",
		21773 to 21777 => "11111111",
		22572 to 22576 => "11111111",
		22647 to 22651 => "11111111",
		22722 to 22726 => "11111111",
		22797 to 22801 => "11111111",
		23596 to 23600 => "11111111",
		23671 to 23675 => "11111111",
		23746 to 23750 => "11111111",
		23821 to 23825 => "11111111",
		24620 to 24624 => "11111111",
		24695 to 24699 => "11111111",
		24770 to 24774 => "11111111",
		24845 to 24849 => "11111111",
		25644 to 25648 => "11111111",
		25719 to 25723 => "11111111",
		25794 to 25798 => "11111111",
		25869 to 25873 => "11111111",
		26668 to 26672 => "11111111",
		26743 to 26747 => "11111111",
		26818 to 26822 => "11111111",
		26893 to 26897 => "11111111",
		27692 to 27696 => "11111111",
		27767 to 27771 => "11111111",
		27842 to 27846 => "11111111",
		27917 to 27921 => "11111111",
		28716 to 28720 => "11111111",
		28791 to 28795 => "11111111",
		28866 to 28870 => "11111111",
		28941 to 28945 => "11111111",
		29740 to 29744 => "11111111",
		29815 to 29819 => "11111111",
		29890 to 29894 => "11111111",
		29965 to 29969 => "11111111",
		30764 to 30768 => "11111111",
		30839 to 30843 => "11111111",
		30914 to 30918 => "11111111",
		30989 to 30993 => "11111111",
		31788 to 31792 => "11111111",
		31863 to 31867 => "11111111",
		31938 to 31942 => "11111111",
		32013 to 32017 => "11111111",
		32812 to 32816 => "11111111",
		32887 to 32891 => "11111111",
		32962 to 32966 => "11111111",
		33037 to 33041 => "11111111",
		33836 to 33840 => "11111111",
		33911 to 33915 => "11111111",
		33986 to 33990 => "11111111",
		34061 to 34065 => "11111111",
		34860 to 34864 => "11111111",
		34935 to 34939 => "11111111",
		35010 to 35014 => "11111111",
		35085 to 35089 => "11111111",
		35884 to 35888 => "11111111",
		35959 to 35963 => "11111111",
		36034 to 36038 => "11111111",
		36109 to 36113 => "11111111",
		36908 to 36912 => "11111111",
		36983 to 36987 => "11111111",
		37058 to 37062 => "11111111",
		37133 to 37137 => "11111111",
		37932 to 37936 => "11111111",
		38007 to 38011 => "11111111",
		38082 to 38086 => "11111111",
		38157 to 38161 => "11111111",
		38956 to 38960 => "11111111",
		39031 to 39035 => "11111111",
		39106 to 39110 => "11111111",
		39181 to 39185 => "11111111",
		39980 to 39984 => "11111111",
		40055 to 40059 => "11111111",
		40130 to 40134 => "11111111",
		40205 to 40209 => "11111111",
		41004 to 41008 => "11111111",
		41079 to 41083 => "11111111",
		41154 to 41158 => "11111111",
		41229 to 41233 => "11111111",
		42028 to 42032 => "11111111",
		42103 to 42107 => "11111111",
		42178 to 42182 => "11111111",
		42253 to 42257 => "11111111",
		43052 to 43056 => "11111111",
		43127 to 43131 => "11111111",
		43202 to 43206 => "11111111",
		43277 to 43281 => "11111111",
		44076 to 44080 => "11111111",
		44151 to 44155 => "11111111",
		44226 to 44230 => "11111111",
		44301 to 44305 => "11111111",
		45100 to 45104 => "11111111",
		45175 to 45179 => "11111111",
		45250 to 45254 => "11111111",
		45325 to 45329 => "11111111",
		46124 to 46128 => "11111111",
		46199 to 46203 => "11111111",
		46274 to 46278 => "11111111",
		46349 to 46353 => "11111111",
		47148 to 47152 => "11111111",
		47223 to 47227 => "11111111",
		47298 to 47302 => "11111111",
		47373 to 47377 => "11111111",
		48172 to 48176 => "11111111",
		48247 to 48251 => "11111111",
		48322 to 48326 => "11111111",
		48397 to 48401 => "11111111",
		49196 to 49200 => "11111111",
		49271 to 49275 => "11111111",
		49346 to 49350 => "11111111",
		49421 to 49425 => "11111111",
		50220 to 50224 => "11111111",
		50295 to 50299 => "11111111",
		50370 to 50374 => "11111111",
		50445 to 50449 => "11111111",
		51244 to 51248 => "11111111",
		51319 to 51323 => "11111111",
		51394 to 51398 => "11111111",
		51469 to 51473 => "11111111",
		52268 to 52272 => "11111111",
		52343 to 52347 => "11111111",
		52418 to 52422 => "11111111",
		52493 to 52497 => "11111111",
		53292 to 53296 => "11111111",
		53367 to 53371 => "11111111",
		53442 to 53446 => "11111111",
		53517 to 53521 => "11111111",
		54316 to 54320 => "11111111",
		54391 to 54395 => "11111111",
		54466 to 54470 => "11111111",
		54541 to 54545 => "11111111",
		55340 to 55344 => "11111111",
		55415 to 55419 => "11111111",
		55490 to 55494 => "11111111",
		55565 to 55569 => "11111111",
		56364 to 56368 => "11111111",
		56439 to 56443 => "11111111",
		56514 to 56518 => "11111111",
		56589 to 56593 => "11111111",
		57388 to 57392 => "11111111",
		57463 to 57467 => "11111111",
		57538 to 57542 => "11111111",
		57613 to 57617 => "11111111",
		58412 to 58416 => "11111111",
		58487 to 58491 => "11111111",
		58562 to 58566 => "11111111",
		58637 to 58641 => "11111111",
		59436 to 59440 => "11111111",
		59511 to 59515 => "11111111",
		59586 to 59590 => "11111111",
		59661 to 59665 => "11111111",
		60460 to 60464 => "11111111",
		60535 to 60539 => "11111111",
		60610 to 60614 => "11111111",
		60685 to 60689 => "11111111",
		61484 to 61488 => "11111111",
		61559 to 61563 => "11111111",
		61634 to 61638 => "11111111",
		61709 to 61713 => "11111111",
		62508 to 62512 => "11111111",
		62583 to 62587 => "11111111",
		62658 to 62662 => "11111111",
		62733 to 62737 => "11111111",
		63532 to 63536 => "11111111",
		63607 to 63611 => "11111111",
		63682 to 63686 => "11111111",
		63757 to 63761 => "11111111",
		64556 to 64560 => "11111111",
		64631 to 64635 => "11111111",
		64706 to 64710 => "11111111",
		64781 to 64785 => "11111111",
		65580 to 65584 => "11111111",
		65655 to 65659 => "11111111",
		65730 to 65734 => "11111111",
		65805 to 65809 => "11111111",
		66604 to 66608 => "11111111",
		66679 to 66683 => "11111111",
		66754 to 66758 => "11111111",
		66829 to 66833 => "11111111",
		67628 to 67632 => "11111111",
		67703 to 67707 => "11111111",
		67778 to 67782 => "11111111",
		67853 to 67857 => "11111111",
		68652 to 68656 => "11111111",
		68727 to 68731 => "11111111",
		68802 to 68806 => "11111111",
		68877 to 68881 => "11111111",
		69676 to 69680 => "11111111",
		69751 to 69755 => "11111111",
		69826 to 69830 => "11111111",
		69901 to 69905 => "11111111",
		70700 to 70704 => "11111111",
		70775 to 70779 => "11111111",
		70850 to 70854 => "11111111",
		70925 to 70929 => "11111111",
		71724 to 71728 => "11111111",
		71799 to 71803 => "11111111",
		71874 to 71878 => "11111111",
		71949 to 71953 => "11111111",
		72748 to 72752 => "11111111",
		72823 to 72827 => "11111111",
		72898 to 72902 => "11111111",
		72973 to 72977 => "11111111",
		73772 to 73776 => "11111111",
		73847 to 73851 => "11111111",
		73922 to 73926 => "11111111",
		73997 to 74001 => "11111111",
		74796 to 74800 => "11111111",
		74871 to 74875 => "11111111",
		74946 to 74950 => "11111111",
		75021 to 75025 => "11111111",
		75820 to 75824 => "11111111",
		75895 to 75899 => "11111111",
		75970 to 75974 => "11111111",
		76045 to 76049 => "11111111",
		76844 to 76848 => "11111111",
		76919 to 76923 => "11111111",
		76994 to 76998 => "11111111",
		77069 to 77073 => "11111111",
		77868 to 77872 => "11111111",
		77943 to 77947 => "11111111",
		78018 to 78022 => "11111111",
		78093 to 78097 => "11111111",
		78892 to 78896 => "11111111",
		78967 to 78971 => "11111111",
		79042 to 79046 => "11111111",
		79117 to 79121 => "11111111",
		79916 to 79920 => "11111111",
		79991 to 79995 => "11111111",
		80066 to 80070 => "11111111",
		80141 to 80145 => "11111111",
		80940 to 81169 => "11111111",
		81964 to 82193 => "11111111",
		82988 to 83217 => "11111111",
		84012 to 84241 => "11111111",
		85036 to 85265 => "11111111",
		86060 to 86064 => "11111111",
		86135 to 86139 => "11111111",
		86210 to 86214 => "11111111",
		86285 to 86289 => "11111111",
		87084 to 87088 => "11111111",
		87159 to 87163 => "11111111",
		87234 to 87238 => "11111111",
		87309 to 87313 => "11111111",
		88108 to 88112 => "11111111",
		88183 to 88187 => "11111111",
		88258 to 88262 => "11111111",
		88333 to 88337 => "11111111",
		89132 to 89136 => "11111111",
		89207 to 89211 => "11111111",
		89282 to 89286 => "11111111",
		89357 to 89361 => "11111111",
		90156 to 90160 => "11111111",
		90231 to 90235 => "11111111",
		90306 to 90310 => "11111111",
		90381 to 90385 => "11111111",
		91180 to 91184 => "11111111",
		91255 to 91259 => "11111111",
		91330 to 91334 => "11111111",
		91405 to 91409 => "11111111",
		92204 to 92208 => "11111111",
		92279 to 92283 => "11111111",
		92354 to 92358 => "11111111",
		92429 to 92433 => "11111111",
		93228 to 93232 => "11111111",
		93303 to 93307 => "11111111",
		93378 to 93382 => "11111111",
		93453 to 93457 => "11111111",
		94252 to 94256 => "11111111",
		94327 to 94331 => "11111111",
		94402 to 94406 => "11111111",
		94477 to 94481 => "11111111",
		95276 to 95280 => "11111111",
		95351 to 95355 => "11111111",
		95426 to 95430 => "11111111",
		95501 to 95505 => "11111111",
		96300 to 96304 => "11111111",
		96375 to 96379 => "11111111",
		96450 to 96454 => "11111111",
		96525 to 96529 => "11111111",
		97324 to 97328 => "11111111",
		97399 to 97403 => "11111111",
		97474 to 97478 => "11111111",
		97549 to 97553 => "11111111",
		98348 to 98352 => "11111111",
		98423 to 98427 => "11111111",
		98498 to 98502 => "11111111",
		98573 to 98577 => "11111111",
		99372 to 99376 => "11111111",
		99447 to 99451 => "11111111",
		99522 to 99526 => "11111111",
		99597 to 99601 => "11111111",
		100396 to 100400 => "11111111",
		100471 to 100475 => "11111111",
		100546 to 100550 => "11111111",
		100621 to 100625 => "11111111",
		101420 to 101424 => "11111111",
		101495 to 101499 => "11111111",
		101570 to 101574 => "11111111",
		101645 to 101649 => "11111111",
		102444 to 102448 => "11111111",
		102519 to 102523 => "11111111",
		102594 to 102598 => "11111111",
		102669 to 102673 => "11111111",
		103468 to 103472 => "11111111",
		103543 to 103547 => "11111111",
		103618 to 103622 => "11111111",
		103693 to 103697 => "11111111",
		104492 to 104496 => "11111111",
		104567 to 104571 => "11111111",
		104642 to 104646 => "11111111",
		104717 to 104721 => "11111111",
		105516 to 105520 => "11111111",
		105591 to 105595 => "11111111",
		105666 to 105670 => "11111111",
		105741 to 105745 => "11111111",
		106540 to 106544 => "11111111",
		106615 to 106619 => "11111111",
		106690 to 106694 => "11111111",
		106765 to 106769 => "11111111",
		107564 to 107568 => "11111111",
		107639 to 107643 => "11111111",
		107714 to 107718 => "11111111",
		107789 to 107793 => "11111111",
		108588 to 108592 => "11111111",
		108663 to 108667 => "11111111",
		108738 to 108742 => "11111111",
		108813 to 108817 => "11111111",
		109612 to 109616 => "11111111",
		109687 to 109691 => "11111111",
		109762 to 109766 => "11111111",
		109837 to 109841 => "11111111",
		110636 to 110640 => "11111111",
		110711 to 110715 => "11111111",
		110786 to 110790 => "11111111",
		110861 to 110865 => "11111111",
		111660 to 111664 => "11111111",
		111735 to 111739 => "11111111",
		111810 to 111814 => "11111111",
		111885 to 111889 => "11111111",
		112684 to 112688 => "11111111",
		112759 to 112763 => "11111111",
		112834 to 112838 => "11111111",
		112909 to 112913 => "11111111",
		113708 to 113712 => "11111111",
		113783 to 113787 => "11111111",
		113858 to 113862 => "11111111",
		113933 to 113937 => "11111111",
		114732 to 114736 => "11111111",
		114807 to 114811 => "11111111",
		114882 to 114886 => "11111111",
		114957 to 114961 => "11111111",
		115756 to 115760 => "11111111",
		115831 to 115835 => "11111111",
		115906 to 115910 => "11111111",
		115981 to 115985 => "11111111",
		116780 to 116784 => "11111111",
		116855 to 116859 => "11111111",
		116930 to 116934 => "11111111",
		117005 to 117009 => "11111111",
		117804 to 117808 => "11111111",
		117879 to 117883 => "11111111",
		117954 to 117958 => "11111111",
		118029 to 118033 => "11111111",
		118828 to 118832 => "11111111",
		118903 to 118907 => "11111111",
		118978 to 118982 => "11111111",
		119053 to 119057 => "11111111",
		119852 to 119856 => "11111111",
		119927 to 119931 => "11111111",
		120002 to 120006 => "11111111",
		120077 to 120081 => "11111111",
		120876 to 120880 => "11111111",
		120951 to 120955 => "11111111",
		121026 to 121030 => "11111111",
		121101 to 121105 => "11111111",
		121900 to 121904 => "11111111",
		121975 to 121979 => "11111111",
		122050 to 122054 => "11111111",
		122125 to 122129 => "11111111",
		122924 to 122928 => "11111111",
		122999 to 123003 => "11111111",
		123074 to 123078 => "11111111",
		123149 to 123153 => "11111111",
		123948 to 123952 => "11111111",
		124023 to 124027 => "11111111",
		124098 to 124102 => "11111111",
		124173 to 124177 => "11111111",
		124972 to 124976 => "11111111",
		125047 to 125051 => "11111111",
		125122 to 125126 => "11111111",
		125197 to 125201 => "11111111",
		125996 to 126000 => "11111111",
		126071 to 126075 => "11111111",
		126146 to 126150 => "11111111",
		126221 to 126225 => "11111111",
		127020 to 127024 => "11111111",
		127095 to 127099 => "11111111",
		127170 to 127174 => "11111111",
		127245 to 127249 => "11111111",
		128044 to 128048 => "11111111",
		128119 to 128123 => "11111111",
		128194 to 128198 => "11111111",
		128269 to 128273 => "11111111",
		129068 to 129072 => "11111111",
		129143 to 129147 => "11111111",
		129218 to 129222 => "11111111",
		129293 to 129297 => "11111111",
		130092 to 130096 => "11111111",
		130167 to 130171 => "11111111",
		130242 to 130246 => "11111111",
		130317 to 130321 => "11111111",
		131116 to 131120 => "11111111",
		131191 to 131195 => "11111111",
		131266 to 131270 => "11111111",
		131341 to 131345 => "11111111",
		132140 to 132144 => "11111111",
		132215 to 132219 => "11111111",
		132290 to 132294 => "11111111",
		132365 to 132369 => "11111111",
		133164 to 133168 => "11111111",
		133239 to 133243 => "11111111",
		133314 to 133318 => "11111111",
		133389 to 133393 => "11111111",
		134188 to 134192 => "11111111",
		134263 to 134267 => "11111111",
		134338 to 134342 => "11111111",
		134413 to 134417 => "11111111",
		135212 to 135216 => "11111111",
		135287 to 135291 => "11111111",
		135362 to 135366 => "11111111",
		135437 to 135441 => "11111111",
		136236 to 136240 => "11111111",
		136311 to 136315 => "11111111",
		136386 to 136390 => "11111111",
		136461 to 136465 => "11111111",
		137260 to 137264 => "11111111",
		137335 to 137339 => "11111111",
		137410 to 137414 => "11111111",
		137485 to 137489 => "11111111",
		138284 to 138288 => "11111111",
		138359 to 138363 => "11111111",
		138434 to 138438 => "11111111",
		138509 to 138513 => "11111111",
		139308 to 139312 => "11111111",
		139383 to 139387 => "11111111",
		139458 to 139462 => "11111111",
		139533 to 139537 => "11111111",
		140332 to 140336 => "11111111",
		140407 to 140411 => "11111111",
		140482 to 140486 => "11111111",
		140557 to 140561 => "11111111",
		141356 to 141360 => "11111111",
		141431 to 141435 => "11111111",
		141506 to 141510 => "11111111",
		141581 to 141585 => "11111111",
		142380 to 142384 => "11111111",
		142455 to 142459 => "11111111",
		142530 to 142534 => "11111111",
		142605 to 142609 => "11111111",
		143404 to 143408 => "11111111",
		143479 to 143483 => "11111111",
		143554 to 143558 => "11111111",
		143629 to 143633 => "11111111",
		144428 to 144432 => "11111111",
		144503 to 144507 => "11111111",
		144578 to 144582 => "11111111",
		144653 to 144657 => "11111111",
		145452 to 145456 => "11111111",
		145527 to 145531 => "11111111",
		145602 to 145606 => "11111111",
		145677 to 145681 => "11111111",
		146476 to 146480 => "11111111",
		146551 to 146555 => "11111111",
		146626 to 146630 => "11111111",
		146701 to 146705 => "11111111",
		147500 to 147504 => "11111111",
		147575 to 147579 => "11111111",
		147650 to 147654 => "11111111",
		147725 to 147729 => "11111111",
		148524 to 148528 => "11111111",
		148599 to 148603 => "11111111",
		148674 to 148678 => "11111111",
		148749 to 148753 => "11111111",
		149548 to 149552 => "11111111",
		149623 to 149627 => "11111111",
		149698 to 149702 => "11111111",
		149773 to 149777 => "11111111",
		150572 to 150576 => "11111111",
		150647 to 150651 => "11111111",
		150722 to 150726 => "11111111",
		150797 to 150801 => "11111111",
		151596 to 151600 => "11111111",
		151671 to 151675 => "11111111",
		151746 to 151750 => "11111111",
		151821 to 151825 => "11111111",
		152620 to 152624 => "11111111",
		152695 to 152699 => "11111111",
		152770 to 152774 => "11111111",
		152845 to 152849 => "11111111",
		153644 to 153648 => "11111111",
		153719 to 153723 => "11111111",
		153794 to 153798 => "11111111",
		153869 to 153873 => "11111111",
		154668 to 154672 => "11111111",
		154743 to 154747 => "11111111",
		154818 to 154822 => "11111111",
		154893 to 154897 => "11111111",
		155692 to 155696 => "11111111",
		155767 to 155771 => "11111111",
		155842 to 155846 => "11111111",
		155917 to 155921 => "11111111",
		156716 to 156720 => "11111111",
		156791 to 156795 => "11111111",
		156866 to 156870 => "11111111",
		156941 to 156945 => "11111111",
		157740 to 157969 => "11111111",
		158764 to 158993 => "11111111",
		159788 to 160017 => "11111111",
		160812 to 161041 => "11111111",
		161836 to 162065 => "11111111",
		162860 to 162864 => "11111111",
		162935 to 162939 => "11111111",
		163010 to 163014 => "11111111",
		163085 to 163089 => "11111111",
		163884 to 163888 => "11111111",
		163959 to 163963 => "11111111",
		164034 to 164038 => "11111111",
		164109 to 164113 => "11111111",
		164908 to 164912 => "11111111",
		164983 to 164987 => "11111111",
		165058 to 165062 => "11111111",
		165133 to 165137 => "11111111",
		165932 to 165936 => "11111111",
		166007 to 166011 => "11111111",
		166082 to 166086 => "11111111",
		166157 to 166161 => "11111111",
		166956 to 166960 => "11111111",
		167031 to 167035 => "11111111",
		167106 to 167110 => "11111111",
		167181 to 167185 => "11111111",
		167980 to 167984 => "11111111",
		168055 to 168059 => "11111111",
		168130 to 168134 => "11111111",
		168205 to 168209 => "11111111",
		169004 to 169008 => "11111111",
		169079 to 169083 => "11111111",
		169154 to 169158 => "11111111",
		169229 to 169233 => "11111111",
		170028 to 170032 => "11111111",
		170103 to 170107 => "11111111",
		170178 to 170182 => "11111111",
		170253 to 170257 => "11111111",
		171052 to 171056 => "11111111",
		171127 to 171131 => "11111111",
		171202 to 171206 => "11111111",
		171277 to 171281 => "11111111",
		172076 to 172080 => "11111111",
		172151 to 172155 => "11111111",
		172226 to 172230 => "11111111",
		172301 to 172305 => "11111111",
		173100 to 173104 => "11111111",
		173175 to 173179 => "11111111",
		173250 to 173254 => "11111111",
		173325 to 173329 => "11111111",
		174124 to 174128 => "11111111",
		174199 to 174203 => "11111111",
		174274 to 174278 => "11111111",
		174349 to 174353 => "11111111",
		175148 to 175152 => "11111111",
		175223 to 175227 => "11111111",
		175298 to 175302 => "11111111",
		175373 to 175377 => "11111111",
		176172 to 176176 => "11111111",
		176247 to 176251 => "11111111",
		176322 to 176326 => "11111111",
		176397 to 176401 => "11111111",
		177196 to 177200 => "11111111",
		177271 to 177275 => "11111111",
		177346 to 177350 => "11111111",
		177421 to 177425 => "11111111",
		178220 to 178224 => "11111111",
		178295 to 178299 => "11111111",
		178370 to 178374 => "11111111",
		178445 to 178449 => "11111111",
		179244 to 179248 => "11111111",
		179319 to 179323 => "11111111",
		179394 to 179398 => "11111111",
		179469 to 179473 => "11111111",
		180268 to 180272 => "11111111",
		180343 to 180347 => "11111111",
		180418 to 180422 => "11111111",
		180493 to 180497 => "11111111",
		181292 to 181296 => "11111111",
		181367 to 181371 => "11111111",
		181442 to 181446 => "11111111",
		181517 to 181521 => "11111111",
		182316 to 182320 => "11111111",
		182391 to 182395 => "11111111",
		182466 to 182470 => "11111111",
		182541 to 182545 => "11111111",
		183340 to 183344 => "11111111",
		183415 to 183419 => "11111111",
		183490 to 183494 => "11111111",
		183565 to 183569 => "11111111",
		184364 to 184368 => "11111111",
		184439 to 184443 => "11111111",
		184514 to 184518 => "11111111",
		184589 to 184593 => "11111111",
		185388 to 185392 => "11111111",
		185463 to 185467 => "11111111",
		185538 to 185542 => "11111111",
		185613 to 185617 => "11111111",
		186412 to 186416 => "11111111",
		186487 to 186491 => "11111111",
		186562 to 186566 => "11111111",
		186637 to 186641 => "11111111",
		187436 to 187440 => "11111111",
		187511 to 187515 => "11111111",
		187586 to 187590 => "11111111",
		187661 to 187665 => "11111111",
		188460 to 188464 => "11111111",
		188535 to 188539 => "11111111",
		188610 to 188614 => "11111111",
		188685 to 188689 => "11111111",
		189484 to 189488 => "11111111",
		189559 to 189563 => "11111111",
		189634 to 189638 => "11111111",
		189709 to 189713 => "11111111",
		190508 to 190512 => "11111111",
		190583 to 190587 => "11111111",
		190658 to 190662 => "11111111",
		190733 to 190737 => "11111111",
		191532 to 191536 => "11111111",
		191607 to 191611 => "11111111",
		191682 to 191686 => "11111111",
		191757 to 191761 => "11111111",
		192556 to 192560 => "11111111",
		192631 to 192635 => "11111111",
		192706 to 192710 => "11111111",
		192781 to 192785 => "11111111",
		193580 to 193584 => "11111111",
		193655 to 193659 => "11111111",
		193730 to 193734 => "11111111",
		193805 to 193809 => "11111111",
		194604 to 194608 => "11111111",
		194679 to 194683 => "11111111",
		194754 to 194758 => "11111111",
		194829 to 194833 => "11111111",
		195628 to 195632 => "11111111",
		195703 to 195707 => "11111111",
		195778 to 195782 => "11111111",
		195853 to 195857 => "11111111",
		196652 to 196656 => "11111111",
		196727 to 196731 => "11111111",
		196802 to 196806 => "11111111",
		196877 to 196881 => "11111111",
		197676 to 197680 => "11111111",
		197751 to 197755 => "11111111",
		197826 to 197830 => "11111111",
		197901 to 197905 => "11111111",
		198700 to 198704 => "11111111",
		198775 to 198779 => "11111111",
		198850 to 198854 => "11111111",
		198925 to 198929 => "11111111",
		199724 to 199728 => "11111111",
		199799 to 199803 => "11111111",
		199874 to 199878 => "11111111",
		199949 to 199953 => "11111111",
		200748 to 200752 => "11111111",
		200823 to 200827 => "11111111",
		200898 to 200902 => "11111111",
		200973 to 200977 => "11111111",
		201772 to 201776 => "11111111",
		201847 to 201851 => "11111111",
		201922 to 201926 => "11111111",
		201997 to 202001 => "11111111",
		202796 to 202800 => "11111111",
		202871 to 202875 => "11111111",
		202946 to 202950 => "11111111",
		203021 to 203025 => "11111111",
		203820 to 203824 => "11111111",
		203895 to 203899 => "11111111",
		203970 to 203974 => "11111111",
		204045 to 204049 => "11111111",
		204844 to 204848 => "11111111",
		204919 to 204923 => "11111111",
		204994 to 204998 => "11111111",
		205069 to 205073 => "11111111",
		205868 to 205872 => "11111111",
		205943 to 205947 => "11111111",
		206018 to 206022 => "11111111",
		206093 to 206097 => "11111111",
		206892 to 206896 => "11111111",
		206967 to 206971 => "11111111",
		207042 to 207046 => "11111111",
		207117 to 207121 => "11111111",
		207916 to 207920 => "11111111",
		207991 to 207995 => "11111111",
		208066 to 208070 => "11111111",
		208141 to 208145 => "11111111",
		208940 to 208944 => "11111111",
		209015 to 209019 => "11111111",
		209090 to 209094 => "11111111",
		209165 to 209169 => "11111111",
		209964 to 209968 => "11111111",
		210039 to 210043 => "11111111",
		210114 to 210118 => "11111111",
		210189 to 210193 => "11111111",
		210988 to 210992 => "11111111",
		211063 to 211067 => "11111111",
		211138 to 211142 => "11111111",
		211213 to 211217 => "11111111",
		212012 to 212016 => "11111111",
		212087 to 212091 => "11111111",
		212162 to 212166 => "11111111",
		212237 to 212241 => "11111111",
		213036 to 213040 => "11111111",
		213111 to 213115 => "11111111",
		213186 to 213190 => "11111111",
		213261 to 213265 => "11111111",
		214060 to 214064 => "11111111",
		214135 to 214139 => "11111111",
		214210 to 214214 => "11111111",
		214285 to 214289 => "11111111",
		215084 to 215088 => "11111111",
		215159 to 215163 => "11111111",
		215234 to 215238 => "11111111",
		215309 to 215313 => "11111111",
		216108 to 216112 => "11111111",
		216183 to 216187 => "11111111",
		216258 to 216262 => "11111111",
		216333 to 216337 => "11111111",
		217132 to 217136 => "11111111",
		217207 to 217211 => "11111111",
		217282 to 217286 => "11111111",
		217357 to 217361 => "11111111",
		218156 to 218160 => "11111111",
		218231 to 218235 => "11111111",
		218306 to 218310 => "11111111",
		218381 to 218385 => "11111111",
		219180 to 219184 => "11111111",
		219255 to 219259 => "11111111",
		219330 to 219334 => "11111111",
		219405 to 219409 => "11111111",
		220204 to 220208 => "11111111",
		220279 to 220283 => "11111111",
		220354 to 220358 => "11111111",
		220429 to 220433 => "11111111",
		221228 to 221232 => "11111111",
		221303 to 221307 => "11111111",
		221378 to 221382 => "11111111",
		221453 to 221457 => "11111111",
		222252 to 222256 => "11111111",
		222327 to 222331 => "11111111",
		222402 to 222406 => "11111111",
		222477 to 222481 => "11111111",
		223276 to 223280 => "11111111",
		223351 to 223355 => "11111111",
		223426 to 223430 => "11111111",
		223501 to 223505 => "11111111",
		224300 to 224304 => "11111111",
		224375 to 224379 => "11111111",
		224450 to 224454 => "11111111",
		224525 to 224529 => "11111111",
		225324 to 225328 => "11111111",
		225399 to 225403 => "11111111",
		225474 to 225478 => "11111111",
		225549 to 225553 => "11111111",
		226348 to 226352 => "11111111",
		226423 to 226427 => "11111111",
		226498 to 226502 => "11111111",
		226573 to 226577 => "11111111",
		227372 to 227376 => "11111111",
		227447 to 227451 => "11111111",
		227522 to 227526 => "11111111",
		227597 to 227601 => "11111111",
		228396 to 228400 => "11111111",
		228471 to 228475 => "11111111",
		228546 to 228550 => "11111111",
		228621 to 228625 => "11111111",
		229420 to 229424 => "11111111",
		229495 to 229499 => "11111111",
		229570 to 229574 => "11111111",
		229645 to 229649 => "11111111",
		230444 to 230448 => "11111111",
		230519 to 230523 => "11111111",
		230594 to 230598 => "11111111",
		230669 to 230673 => "11111111",
		231468 to 231472 => "11111111",
		231543 to 231547 => "11111111",
		231618 to 231622 => "11111111",
		231693 to 231697 => "11111111",
		232492 to 232496 => "11111111",
		232567 to 232571 => "11111111",
		232642 to 232646 => "11111111",
		232717 to 232721 => "11111111",
		233516 to 233520 => "11111111",
		233591 to 233595 => "11111111",
		233666 to 233670 => "11111111",
		233741 to 233745 => "11111111",
		234540 to 234769 => "11111111",
		235564 to 235793 => "11111111",
		236588 to 236817 => "11111111",
		237612 to 237841 => "11111111",
		238636 to 238865 => "11111111",
