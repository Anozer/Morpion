		49270 => x"FF",
		49271 => x"FF",
		49272 => x"FF",
		49273 => x"FF",
		49274 => x"FF",
		49275 => x"FF",
		49276 => x"FF",
		49277 => x"FF",
		49278 => x"FF",
		49279 => x"FF",
		49280 => x"FF",
		49281 => x"FF",
		49282 => x"FF",
		49283 => x"FF",
		49284 => x"FF",
		49285 => x"FF",
		49286 => x"FF",
		49287 => x"FF",
		49288 => x"FF",
		49289 => x"FF",
		49290 => x"FF",
		49291 => x"FF",
		49292 => x"FF",
		49293 => x"FF",
		49294 => x"FF",
		49295 => x"FF",
		49296 => x"FF",
		49297 => x"FF",
		49298 => x"FF",
		49299 => x"FF",
		49300 => x"FF",
		49301 => x"FF",
		49302 => x"FF",
		49303 => x"FF",
		49304 => x"FF",
		49305 => x"FF",
		49306 => x"FF",
		49307 => x"FF",
		49308 => x"FF",
		49309 => x"FF",
		49310 => x"FF",
		49311 => x"FF",
		49312 => x"FF",
		49313 => x"FF",
		49314 => x"FF",
		49315 => x"FF",
		49316 => x"FF",
		49317 => x"FF",
		49318 => x"FF",
		49319 => x"FF",
		49320 => x"FF",
		49321 => x"FF",
		49322 => x"FF",
		49323 => x"FF",
		49324 => x"FF",
		49325 => x"FF",
		49326 => x"FF",
		49327 => x"FF",
		49328 => x"FF",
		49329 => x"FF",
		49330 => x"FF",
		49331 => x"FF",
		49332 => x"FF",
		49333 => x"FF",
		49334 => x"FF",
		49335 => x"FF",
		49336 => x"FF",
		49337 => x"FF",
		49338 => x"FF",
		49339 => x"FF",
		49340 => x"FF",
		49341 => x"FF",
		49342 => x"FF",
		49343 => x"FF",
		49344 => x"FF",
		49345 => x"FF",
		49346 => x"FF",
		49347 => x"FF",
		49348 => x"FF",
		49349 => x"FF",
		49350 => x"FF",
		49351 => x"FF",
		49352 => x"FF",
		49353 => x"FF",
		49354 => x"FF",
		49355 => x"FF",
		49356 => x"FF",
		49357 => x"FF",
		49358 => x"FF",
		49359 => x"FF",
		49360 => x"FF",
		49361 => x"FF",
		49362 => x"FF",
		49363 => x"FF",
		49364 => x"FF",
		49365 => x"FF",
		49366 => x"FF",
		49367 => x"FF",
		49368 => x"FF",
		49369 => x"FF",
		49370 => x"FF",
		49371 => x"FF",
		49372 => x"FF",
		49373 => x"FF",
		49374 => x"FF",
		49375 => x"FF",
		49376 => x"FF",
		49377 => x"FF",
		49378 => x"FF",
		49379 => x"FF",
		49380 => x"FF",
		49381 => x"FF",
		49382 => x"FF",
		49383 => x"FF",
		49384 => x"FF",
		49385 => x"FF",
		49386 => x"FF",
		49387 => x"FF",
		49388 => x"FF",
		49389 => x"FF",
		49390 => x"FF",
		49391 => x"FF",
		49392 => x"FF",
		49393 => x"FF",
		49394 => x"FF",
		49395 => x"FF",
		49396 => x"FF",
		49397 => x"FF",
		49398 => x"FF",
		49399 => x"FF",
		49400 => x"FF",
		49401 => x"FF",
		49402 => x"FF",
		49403 => x"FF",
		49404 => x"FF",
		49405 => x"FF",
		49406 => x"FF",
		49407 => x"FF",
		49408 => x"FF",
		49409 => x"FF",
		49410 => x"FF",
		49411 => x"FF",
		49412 => x"FF",
		49413 => x"FF",
		49414 => x"FF",
		49415 => x"FF",
		49416 => x"FF",
		49417 => x"FF",
		49418 => x"FF",
		49419 => x"FF",
		49420 => x"FF",
		49421 => x"FF",
		49422 => x"FF",
		49423 => x"FF",
		49424 => x"FF",
		49425 => x"FF",
		49426 => x"FF",
		49427 => x"FF",
		49428 => x"FF",
		49429 => x"FF",
		49430 => x"FF",
		49431 => x"FF",
		49432 => x"FF",
		49433 => x"FF",
		49434 => x"FF",
		49435 => x"FF",
		49436 => x"FF",
		49437 => x"FF",
		49438 => x"FF",
		49439 => x"FF",
		49440 => x"FF",
		49441 => x"FF",
		49442 => x"FF",
		49443 => x"FF",
		49444 => x"FF",
		49445 => x"FF",
		49446 => x"FF",
		49447 => x"FF",
		49448 => x"FF",
		49449 => x"FF",
		49450 => x"FF",
		49451 => x"FF",
		49452 => x"FF",
		49453 => x"FF",
		49454 => x"FF",
		49455 => x"FF",
		49456 => x"FF",
		49457 => x"FF",
		49458 => x"FF",
		49459 => x"FF",
		49460 => x"FF",
		49461 => x"FF",
		49462 => x"FF",
		49463 => x"FF",
		49464 => x"FF",
		49465 => x"FF",
		49466 => x"FF",
		49467 => x"FF",
		49468 => x"FF",
		49469 => x"FF",
		49470 => x"FF",
		49471 => x"FF",
		49472 => x"FF",
		49473 => x"FF",
		49474 => x"FF",
		49475 => x"FF",
		49476 => x"FF",
		49477 => x"FF",
		49478 => x"FF",
		49479 => x"FF",
		49480 => x"FF",
		49481 => x"FF",
		49482 => x"FF",
		49483 => x"FF",
		49484 => x"FF",
		49485 => x"FF",
		49486 => x"FF",
		49487 => x"FF",
		49488 => x"FF",
		49489 => x"FF",
		49490 => x"FF",
		49491 => x"FF",
		49492 => x"FF",
		49493 => x"FF",
		49494 => x"FF",
		49495 => x"FF",
		49496 => x"FF",
		49497 => x"FF",
		49498 => x"FF",
		49499 => x"FF",
		49500 => x"FF",
		49501 => x"FF",
		49502 => x"FF",
		49503 => x"FF",
		49504 => x"FF",
		49505 => x"FF",
		49506 => x"FF",
		49507 => x"FF",
		49508 => x"FF",
		49509 => x"FF",
		49510 => x"FF",
		49511 => x"FF",
		49512 => x"FF",
		49513 => x"FF",
		49514 => x"FF",
		49515 => x"FF",
		49516 => x"FF",
		49517 => x"FF",
		49518 => x"FF",
		49519 => x"FF",
		49520 => x"FF",
		49521 => x"FF",
		49522 => x"FF",
		49523 => x"FF",
		49524 => x"FF",
		49525 => x"FF",
		49526 => x"FF",
		49527 => x"FF",
		49528 => x"FF",
		49529 => x"FF",
		49530 => x"FF",
		49531 => x"FF",
		49532 => x"FF",
		49533 => x"FF",
		49534 => x"FF",
		49535 => x"FF",
		49536 => x"FF",
		49537 => x"FF",
		49538 => x"FF",
		49539 => x"FF",
		49540 => x"FF",
		49541 => x"FF",
		49542 => x"FF",
		49543 => x"FF",
		49544 => x"FF",
		49545 => x"FF",
		49546 => x"FF",
		49547 => x"FF",
		49548 => x"FF",
		49549 => x"FF",
		49550 => x"FF",
		49551 => x"FF",
		49552 => x"FF",
		49553 => x"FF",
		49554 => x"FF",
		49555 => x"FF",
		49556 => x"FF",
		49557 => x"FF",
		49558 => x"FF",
		49559 => x"FF",
		49560 => x"FF",
		49561 => x"FF",
		49562 => x"FF",
		49563 => x"FF",
		49564 => x"FF",
		49565 => x"FF",
		49566 => x"FF",
		49567 => x"FF",
		49568 => x"FF",
		49569 => x"FF",
		49570 => x"FF",
		49571 => x"FF",
		49572 => x"FF",
		49573 => x"FF",
		49574 => x"FF",
		49575 => x"FF",
		49576 => x"FF",
		49577 => x"FF",
		49578 => x"FF",
		49579 => x"FF",
		49580 => x"FF",
		49581 => x"FF",
		49582 => x"FF",
		49583 => x"FF",
		49584 => x"FF",
		49585 => x"FF",
		49586 => x"FF",
		49587 => x"FF",
		49588 => x"FF",
		49589 => x"FF",
		49590 => x"FF",
		49591 => x"FF",
		49592 => x"FF",
		49593 => x"FF",
		49594 => x"FF",
		49595 => x"FF",
		49596 => x"FF",
		49597 => x"FF",
		49598 => x"FF",
		49599 => x"FF",
		49600 => x"FF",
		49601 => x"FF",
		49602 => x"FF",
		49603 => x"FF",
		49604 => x"FF",
		49605 => x"FF",
		49606 => x"FF",
		49607 => x"FF",
		49608 => x"FF",
		49609 => x"FF",
		49610 => x"FF",
		49611 => x"FF",
		49612 => x"FF",
		49613 => x"FF",
		49614 => x"FF",
		49615 => x"FF",
		49616 => x"FF",
		49617 => x"FF",
		49618 => x"FF",
		49619 => x"FF",
		49620 => x"FF",
		49621 => x"FF",
		49622 => x"FF",
		49623 => x"FF",
		49624 => x"FF",
		49625 => x"FF",
		49626 => x"FF",
		49627 => x"FF",
		49628 => x"FF",
		49629 => x"FF",
		49630 => x"FF",
		49631 => x"FF",
		49632 => x"FF",
		49633 => x"FF",
		49634 => x"FF",
		49635 => x"FF",
		49636 => x"FF",
		49637 => x"FF",
		49638 => x"FF",
		49639 => x"FF",
		49640 => x"FF",
		49641 => x"FF",
		49642 => x"FF",
		49643 => x"FF",
		49644 => x"FF",
		49645 => x"FF",
		49646 => x"FF",
		49647 => x"FF",
		49648 => x"FF",
		49649 => x"FF",
		50294 => x"FF",
		50295 => x"FF",
		50296 => x"FF",
		50297 => x"FF",
		50298 => x"FF",
		50299 => x"FF",
		50300 => x"FF",
		50301 => x"FF",
		50302 => x"FF",
		50303 => x"FF",
		50304 => x"FF",
		50305 => x"FF",
		50306 => x"FF",
		50307 => x"FF",
		50308 => x"FF",
		50309 => x"FF",
		50310 => x"FF",
		50311 => x"FF",
		50312 => x"FF",
		50313 => x"FF",
		50314 => x"FF",
		50315 => x"FF",
		50316 => x"FF",
		50317 => x"FF",
		50318 => x"FF",
		50319 => x"FF",
		50320 => x"FF",
		50321 => x"FF",
		50322 => x"FF",
		50323 => x"FF",
		50324 => x"FF",
		50325 => x"FF",
		50326 => x"FF",
		50327 => x"FF",
		50328 => x"FF",
		50329 => x"FF",
		50330 => x"FF",
		50331 => x"FF",
		50332 => x"FF",
		50333 => x"FF",
		50334 => x"FF",
		50335 => x"FF",
		50336 => x"FF",
		50337 => x"FF",
		50338 => x"FF",
		50339 => x"FF",
		50340 => x"FF",
		50341 => x"FF",
		50342 => x"FF",
		50343 => x"FF",
		50344 => x"FF",
		50345 => x"FF",
		50346 => x"FF",
		50347 => x"FF",
		50348 => x"FF",
		50349 => x"FF",
		50350 => x"FF",
		50351 => x"FF",
		50352 => x"FF",
		50353 => x"FF",
		50354 => x"FF",
		50355 => x"FF",
		50356 => x"FF",
		50357 => x"FF",
		50358 => x"FF",
		50359 => x"FF",
		50360 => x"FF",
		50361 => x"FF",
		50362 => x"FF",
		50363 => x"FF",
		50364 => x"FF",
		50365 => x"FF",
		50366 => x"FF",
		50367 => x"FF",
		50368 => x"FF",
		50369 => x"FF",
		50370 => x"FF",
		50371 => x"FF",
		50372 => x"FF",
		50373 => x"FF",
		50374 => x"FF",
		50375 => x"FF",
		50376 => x"FF",
		50377 => x"FF",
		50378 => x"FF",
		50379 => x"FF",
		50380 => x"FF",
		50381 => x"FF",
		50382 => x"FF",
		50383 => x"FF",
		50384 => x"FF",
		50385 => x"FF",
		50386 => x"FF",
		50387 => x"FF",
		50388 => x"FF",
		50389 => x"FF",
		50390 => x"FF",
		50391 => x"FF",
		50392 => x"FF",
		50393 => x"FF",
		50394 => x"FF",
		50395 => x"FF",
		50396 => x"FF",
		50397 => x"FF",
		50398 => x"FF",
		50399 => x"FF",
		50400 => x"FF",
		50401 => x"FF",
		50402 => x"FF",
		50403 => x"FF",
		50404 => x"FF",
		50405 => x"FF",
		50406 => x"FF",
		50407 => x"FF",
		50408 => x"FF",
		50409 => x"FF",
		50410 => x"FF",
		50411 => x"FF",
		50412 => x"FF",
		50413 => x"FF",
		50414 => x"FF",
		50415 => x"FF",
		50416 => x"FF",
		50417 => x"FF",
		50418 => x"FF",
		50419 => x"FF",
		50420 => x"FF",
		50421 => x"FF",
		50422 => x"FF",
		50423 => x"FF",
		50424 => x"FF",
		50425 => x"FF",
		50426 => x"FF",
		50427 => x"FF",
		50428 => x"FF",
		50429 => x"FF",
		50430 => x"FF",
		50431 => x"FF",
		50432 => x"FF",
		50433 => x"FF",
		50434 => x"FF",
		50435 => x"FF",
		50436 => x"FF",
		50437 => x"FF",
		50438 => x"FF",
		50439 => x"FF",
		50440 => x"FF",
		50441 => x"FF",
		50442 => x"FF",
		50443 => x"FF",
		50444 => x"FF",
		50445 => x"FF",
		50446 => x"FF",
		50447 => x"FF",
		50448 => x"FF",
		50449 => x"FF",
		50450 => x"FF",
		50451 => x"FF",
		50452 => x"FF",
		50453 => x"FF",
		50454 => x"FF",
		50455 => x"FF",
		50456 => x"FF",
		50457 => x"FF",
		50458 => x"FF",
		50459 => x"FF",
		50460 => x"FF",
		50461 => x"FF",
		50462 => x"FF",
		50463 => x"FF",
		50464 => x"FF",
		50465 => x"FF",
		50466 => x"FF",
		50467 => x"FF",
		50468 => x"FF",
		50469 => x"FF",
		50470 => x"FF",
		50471 => x"FF",
		50472 => x"FF",
		50473 => x"FF",
		50474 => x"FF",
		50475 => x"FF",
		50476 => x"FF",
		50477 => x"FF",
		50478 => x"FF",
		50479 => x"FF",
		50480 => x"FF",
		50481 => x"FF",
		50482 => x"FF",
		50483 => x"FF",
		50484 => x"FF",
		50485 => x"FF",
		50486 => x"FF",
		50487 => x"FF",
		50488 => x"FF",
		50489 => x"FF",
		50490 => x"FF",
		50491 => x"FF",
		50492 => x"FF",
		50493 => x"FF",
		50494 => x"FF",
		50495 => x"FF",
		50496 => x"FF",
		50497 => x"FF",
		50498 => x"FF",
		50499 => x"FF",
		50500 => x"FF",
		50501 => x"FF",
		50502 => x"FF",
		50503 => x"FF",
		50504 => x"FF",
		50505 => x"FF",
		50506 => x"FF",
		50507 => x"FF",
		50508 => x"FF",
		50509 => x"FF",
		50510 => x"FF",
		50511 => x"FF",
		50512 => x"FF",
		50513 => x"FF",
		50514 => x"FF",
		50515 => x"FF",
		50516 => x"FF",
		50517 => x"FF",
		50518 => x"FF",
		50519 => x"FF",
		50520 => x"FF",
		50521 => x"FF",
		50522 => x"FF",
		50523 => x"FF",
		50524 => x"FF",
		50525 => x"FF",
		50526 => x"FF",
		50527 => x"FF",
		50528 => x"FF",
		50529 => x"FF",
		50530 => x"FF",
		50531 => x"FF",
		50532 => x"FF",
		50533 => x"FF",
		50534 => x"FF",
		50535 => x"FF",
		50536 => x"FF",
		50537 => x"FF",
		50538 => x"FF",
		50539 => x"FF",
		50540 => x"FF",
		50541 => x"FF",
		50542 => x"FF",
		50543 => x"FF",
		50544 => x"FF",
		50545 => x"FF",
		50546 => x"FF",
		50547 => x"FF",
		50548 => x"FF",
		50549 => x"FF",
		50550 => x"FF",
		50551 => x"FF",
		50552 => x"FF",
		50553 => x"FF",
		50554 => x"FF",
		50555 => x"FF",
		50556 => x"FF",
		50557 => x"FF",
		50558 => x"FF",
		50559 => x"FF",
		50560 => x"FF",
		50561 => x"FF",
		50562 => x"FF",
		50563 => x"FF",
		50564 => x"FF",
		50565 => x"FF",
		50566 => x"FF",
		50567 => x"FF",
		50568 => x"FF",
		50569 => x"FF",
		50570 => x"FF",
		50571 => x"FF",
		50572 => x"FF",
		50573 => x"FF",
		50574 => x"FF",
		50575 => x"FF",
		50576 => x"FF",
		50577 => x"FF",
		50578 => x"FF",
		50579 => x"FF",
		50580 => x"FF",
		50581 => x"FF",
		50582 => x"FF",
		50583 => x"FF",
		50584 => x"FF",
		50585 => x"FF",
		50586 => x"FF",
		50587 => x"FF",
		50588 => x"FF",
		50589 => x"FF",
		50590 => x"FF",
		50591 => x"FF",
		50592 => x"FF",
		50593 => x"FF",
		50594 => x"FF",
		50595 => x"FF",
		50596 => x"FF",
		50597 => x"FF",
		50598 => x"FF",
		50599 => x"FF",
		50600 => x"FF",
		50601 => x"FF",
		50602 => x"FF",
		50603 => x"FF",
		50604 => x"FF",
		50605 => x"FF",
		50606 => x"FF",
		50607 => x"FF",
		50608 => x"FF",
		50609 => x"FF",
		50610 => x"FF",
		50611 => x"FF",
		50612 => x"FF",
		50613 => x"FF",
		50614 => x"FF",
		50615 => x"FF",
		50616 => x"FF",
		50617 => x"FF",
		50618 => x"FF",
		50619 => x"FF",
		50620 => x"FF",
		50621 => x"FF",
		50622 => x"FF",
		50623 => x"FF",
		50624 => x"FF",
		50625 => x"FF",
		50626 => x"FF",
		50627 => x"FF",
		50628 => x"FF",
		50629 => x"FF",
		50630 => x"FF",
		50631 => x"FF",
		50632 => x"FF",
		50633 => x"FF",
		50634 => x"FF",
		50635 => x"FF",
		50636 => x"FF",
		50637 => x"FF",
		50638 => x"FF",
		50639 => x"FF",
		50640 => x"FF",
		50641 => x"FF",
		50642 => x"FF",
		50643 => x"FF",
		50644 => x"FF",
		50645 => x"FF",
		50646 => x"FF",
		50647 => x"FF",
		50648 => x"FF",
		50649 => x"FF",
		50650 => x"FF",
		50651 => x"FF",
		50652 => x"FF",
		50653 => x"FF",
		50654 => x"FF",
		50655 => x"FF",
		50656 => x"FF",
		50657 => x"FF",
		50658 => x"FF",
		50659 => x"FF",
		50660 => x"FF",
		50661 => x"FF",
		50662 => x"FF",
		50663 => x"FF",
		50664 => x"FF",
		50665 => x"FF",
		50666 => x"FF",
		50667 => x"FF",
		50668 => x"FF",
		50669 => x"FF",
		50670 => x"FF",
		50671 => x"FF",
		50672 => x"FF",
		50673 => x"FF",
		51318 => x"FF",
		51319 => x"FF",
		51320 => x"FF",
		51321 => x"FF",
		51322 => x"FF",
		51323 => x"FF",
		51324 => x"FF",
		51325 => x"FF",
		51326 => x"FF",
		51327 => x"FF",
		51328 => x"FF",
		51329 => x"FF",
		51330 => x"FF",
		51331 => x"FF",
		51332 => x"FF",
		51333 => x"FF",
		51334 => x"FF",
		51335 => x"FF",
		51336 => x"FF",
		51337 => x"FF",
		51338 => x"FF",
		51339 => x"FF",
		51340 => x"FF",
		51341 => x"FF",
		51342 => x"FF",
		51343 => x"FF",
		51344 => x"FF",
		51345 => x"FF",
		51346 => x"FF",
		51347 => x"FF",
		51348 => x"FF",
		51349 => x"FF",
		51350 => x"FF",
		51351 => x"FF",
		51352 => x"FF",
		51353 => x"FF",
		51354 => x"FF",
		51355 => x"FF",
		51356 => x"FF",
		51357 => x"FF",
		51358 => x"FF",
		51359 => x"FF",
		51360 => x"FF",
		51361 => x"FF",
		51362 => x"FF",
		51363 => x"FF",
		51364 => x"FF",
		51365 => x"FF",
		51366 => x"FF",
		51367 => x"FF",
		51368 => x"FF",
		51369 => x"FF",
		51370 => x"FF",
		51371 => x"FF",
		51372 => x"FF",
		51373 => x"FF",
		51374 => x"FF",
		51375 => x"FF",
		51376 => x"FF",
		51377 => x"FF",
		51378 => x"FF",
		51379 => x"FF",
		51380 => x"FF",
		51381 => x"FF",
		51382 => x"FF",
		51383 => x"FF",
		51384 => x"FF",
		51385 => x"FF",
		51386 => x"FF",
		51387 => x"FF",
		51388 => x"FF",
		51389 => x"FF",
		51390 => x"FF",
		51391 => x"FF",
		51392 => x"FF",
		51393 => x"FF",
		51394 => x"FF",
		51395 => x"FF",
		51396 => x"FF",
		51397 => x"FF",
		51398 => x"FF",
		51399 => x"FF",
		51400 => x"FF",
		51401 => x"FF",
		51402 => x"FF",
		51403 => x"FF",
		51404 => x"FF",
		51405 => x"FF",
		51406 => x"FF",
		51407 => x"FF",
		51408 => x"FF",
		51409 => x"FF",
		51410 => x"FF",
		51411 => x"FF",
		51412 => x"FF",
		51413 => x"FF",
		51414 => x"FF",
		51415 => x"FF",
		51416 => x"FF",
		51417 => x"FF",
		51418 => x"FF",
		51419 => x"FF",
		51420 => x"FF",
		51421 => x"FF",
		51422 => x"FF",
		51423 => x"FF",
		51424 => x"FF",
		51425 => x"FF",
		51426 => x"FF",
		51427 => x"FF",
		51428 => x"FF",
		51429 => x"FF",
		51430 => x"FF",
		51431 => x"FF",
		51432 => x"FF",
		51433 => x"FF",
		51434 => x"FF",
		51435 => x"FF",
		51436 => x"FF",
		51437 => x"FF",
		51438 => x"FF",
		51439 => x"FF",
		51440 => x"FF",
		51441 => x"FF",
		51442 => x"FF",
		51443 => x"FF",
		51444 => x"FF",
		51445 => x"FF",
		51446 => x"FF",
		51447 => x"FF",
		51448 => x"FF",
		51449 => x"FF",
		51450 => x"FF",
		51451 => x"FF",
		51452 => x"FF",
		51453 => x"FF",
		51454 => x"FF",
		51455 => x"FF",
		51456 => x"FF",
		51457 => x"FF",
		51458 => x"FF",
		51459 => x"FF",
		51460 => x"FF",
		51461 => x"FF",
		51462 => x"FF",
		51463 => x"FF",
		51464 => x"FF",
		51465 => x"FF",
		51466 => x"FF",
		51467 => x"FF",
		51468 => x"FF",
		51469 => x"FF",
		51470 => x"FF",
		51471 => x"FF",
		51472 => x"FF",
		51473 => x"FF",
		51474 => x"FF",
		51475 => x"FF",
		51476 => x"FF",
		51477 => x"FF",
		51478 => x"FF",
		51479 => x"FF",
		51480 => x"FF",
		51481 => x"FF",
		51482 => x"FF",
		51483 => x"FF",
		51484 => x"FF",
		51485 => x"FF",
		51486 => x"FF",
		51487 => x"FF",
		51488 => x"FF",
		51489 => x"FF",
		51490 => x"FF",
		51491 => x"FF",
		51492 => x"FF",
		51493 => x"FF",
		51494 => x"FF",
		51495 => x"FF",
		51496 => x"FF",
		51497 => x"FF",
		51498 => x"FF",
		51499 => x"FF",
		51500 => x"FF",
		51501 => x"FF",
		51502 => x"FF",
		51503 => x"FF",
		51504 => x"FF",
		51505 => x"FF",
		51506 => x"FF",
		51507 => x"FF",
		51508 => x"FF",
		51509 => x"FF",
		51510 => x"FF",
		51511 => x"FF",
		51512 => x"FF",
		51513 => x"FF",
		51514 => x"FF",
		51515 => x"FF",
		51516 => x"FF",
		51517 => x"FF",
		51518 => x"FF",
		51519 => x"FF",
		51520 => x"FF",
		51521 => x"FF",
		51522 => x"FF",
		51523 => x"FF",
		51524 => x"FF",
		51525 => x"FF",
		51526 => x"FF",
		51527 => x"FF",
		51528 => x"FF",
		51529 => x"FF",
		51530 => x"FF",
		51531 => x"FF",
		51532 => x"FF",
		51533 => x"FF",
		51534 => x"FF",
		51535 => x"FF",
		51536 => x"FF",
		51537 => x"FF",
		51538 => x"FF",
		51539 => x"FF",
		51540 => x"FF",
		51541 => x"FF",
		51542 => x"FF",
		51543 => x"FF",
		51544 => x"FF",
		51545 => x"FF",
		51546 => x"FF",
		51547 => x"FF",
		51548 => x"FF",
		51549 => x"FF",
		51550 => x"FF",
		51551 => x"FF",
		51552 => x"FF",
		51553 => x"FF",
		51554 => x"FF",
		51555 => x"FF",
		51556 => x"FF",
		51557 => x"FF",
		51558 => x"FF",
		51559 => x"FF",
		51560 => x"FF",
		51561 => x"FF",
		51562 => x"FF",
		51563 => x"FF",
		51564 => x"FF",
		51565 => x"FF",
		51566 => x"FF",
		51567 => x"FF",
		51568 => x"FF",
		51569 => x"FF",
		51570 => x"FF",
		51571 => x"FF",
		51572 => x"FF",
		51573 => x"FF",
		51574 => x"FF",
		51575 => x"FF",
		51576 => x"FF",
		51577 => x"FF",
		51578 => x"FF",
		51579 => x"FF",
		51580 => x"FF",
		51581 => x"FF",
		51582 => x"FF",
		51583 => x"FF",
		51584 => x"FF",
		51585 => x"FF",
		51586 => x"FF",
		51587 => x"FF",
		51588 => x"FF",
		51589 => x"FF",
		51590 => x"FF",
		51591 => x"FF",
		51592 => x"FF",
		51593 => x"FF",
		51594 => x"FF",
		51595 => x"FF",
		51596 => x"FF",
		51597 => x"FF",
		51598 => x"FF",
		51599 => x"FF",
		51600 => x"FF",
		51601 => x"FF",
		51602 => x"FF",
		51603 => x"FF",
		51604 => x"FF",
		51605 => x"FF",
		51606 => x"FF",
		51607 => x"FF",
		51608 => x"FF",
		51609 => x"FF",
		51610 => x"FF",
		51611 => x"FF",
		51612 => x"FF",
		51613 => x"FF",
		51614 => x"FF",
		51615 => x"FF",
		51616 => x"FF",
		51617 => x"FF",
		51618 => x"FF",
		51619 => x"FF",
		51620 => x"FF",
		51621 => x"FF",
		51622 => x"FF",
		51623 => x"FF",
		51624 => x"FF",
		51625 => x"FF",
		51626 => x"FF",
		51627 => x"FF",
		51628 => x"FF",
		51629 => x"FF",
		51630 => x"FF",
		51631 => x"FF",
		51632 => x"FF",
		51633 => x"FF",
		51634 => x"FF",
		51635 => x"FF",
		51636 => x"FF",
		51637 => x"FF",
		51638 => x"FF",
		51639 => x"FF",
		51640 => x"FF",
		51641 => x"FF",
		51642 => x"FF",
		51643 => x"FF",
		51644 => x"FF",
		51645 => x"FF",
		51646 => x"FF",
		51647 => x"FF",
		51648 => x"FF",
		51649 => x"FF",
		51650 => x"FF",
		51651 => x"FF",
		51652 => x"FF",
		51653 => x"FF",
		51654 => x"FF",
		51655 => x"FF",
		51656 => x"FF",
		51657 => x"FF",
		51658 => x"FF",
		51659 => x"FF",
		51660 => x"FF",
		51661 => x"FF",
		51662 => x"FF",
		51663 => x"FF",
		51664 => x"FF",
		51665 => x"FF",
		51666 => x"FF",
		51667 => x"FF",
		51668 => x"FF",
		51669 => x"FF",
		51670 => x"FF",
		51671 => x"FF",
		51672 => x"FF",
		51673 => x"FF",
		51674 => x"FF",
		51675 => x"FF",
		51676 => x"FF",
		51677 => x"FF",
		51678 => x"FF",
		51679 => x"FF",
		51680 => x"FF",
		51681 => x"FF",
		51682 => x"FF",
		51683 => x"FF",
		51684 => x"FF",
		51685 => x"FF",
		51686 => x"FF",
		51687 => x"FF",
		51688 => x"FF",
		51689 => x"FF",
		51690 => x"FF",
		51691 => x"FF",
		51692 => x"FF",
		51693 => x"FF",
		51694 => x"FF",
		51695 => x"FF",
		51696 => x"FF",
		51697 => x"FF",
		52342 => x"FF",
		52343 => x"FF",
		52344 => x"FF",
		52345 => x"FF",
		52346 => x"FF",
		52347 => x"FF",
		52348 => x"FF",
		52349 => x"FF",
		52350 => x"FF",
		52351 => x"FF",
		52352 => x"FF",
		52353 => x"FF",
		52354 => x"FF",
		52355 => x"FF",
		52356 => x"FF",
		52357 => x"FF",
		52358 => x"FF",
		52359 => x"FF",
		52360 => x"FF",
		52361 => x"FF",
		52362 => x"FF",
		52363 => x"FF",
		52364 => x"FF",
		52365 => x"FF",
		52366 => x"FF",
		52367 => x"FF",
		52368 => x"FF",
		52369 => x"FF",
		52370 => x"FF",
		52371 => x"FF",
		52372 => x"FF",
		52373 => x"FF",
		52374 => x"FF",
		52375 => x"FF",
		52376 => x"FF",
		52377 => x"FF",
		52378 => x"FF",
		52379 => x"FF",
		52380 => x"FF",
		52381 => x"FF",
		52382 => x"FF",
		52383 => x"FF",
		52384 => x"FF",
		52385 => x"FF",
		52386 => x"FF",
		52387 => x"FF",
		52388 => x"FF",
		52389 => x"FF",
		52390 => x"FF",
		52391 => x"FF",
		52392 => x"FF",
		52393 => x"FF",
		52394 => x"FF",
		52395 => x"FF",
		52396 => x"FF",
		52397 => x"FF",
		52398 => x"FF",
		52399 => x"FF",
		52400 => x"FF",
		52401 => x"FF",
		52402 => x"FF",
		52403 => x"FF",
		52404 => x"FF",
		52405 => x"FF",
		52406 => x"FF",
		52407 => x"FF",
		52408 => x"FF",
		52409 => x"FF",
		52410 => x"FF",
		52411 => x"FF",
		52412 => x"FF",
		52413 => x"FF",
		52414 => x"FF",
		52415 => x"FF",
		52416 => x"FF",
		52417 => x"FF",
		52418 => x"FF",
		52419 => x"FF",
		52420 => x"FF",
		52421 => x"FF",
		52422 => x"FF",
		52423 => x"FF",
		52424 => x"FF",
		52425 => x"FF",
		52426 => x"FF",
		52427 => x"FF",
		52428 => x"FF",
		52429 => x"FF",
		52430 => x"FF",
		52431 => x"FF",
		52432 => x"FF",
		52433 => x"FF",
		52434 => x"FF",
		52435 => x"FF",
		52436 => x"FF",
		52437 => x"FF",
		52438 => x"FF",
		52439 => x"FF",
		52440 => x"FF",
		52441 => x"FF",
		52442 => x"FF",
		52443 => x"FF",
		52444 => x"FF",
		52445 => x"FF",
		52446 => x"FF",
		52447 => x"FF",
		52448 => x"FF",
		52449 => x"FF",
		52450 => x"FF",
		52451 => x"FF",
		52452 => x"FF",
		52453 => x"FF",
		52454 => x"FF",
		52455 => x"FF",
		52456 => x"FF",
		52457 => x"FF",
		52458 => x"FF",
		52459 => x"FF",
		52460 => x"FF",
		52461 => x"FF",
		52462 => x"FF",
		52463 => x"FF",
		52464 => x"FF",
		52465 => x"FF",
		52466 => x"FF",
		52467 => x"FF",
		52468 => x"FF",
		52469 => x"FF",
		52470 => x"FF",
		52471 => x"FF",
		52472 => x"FF",
		52473 => x"FF",
		52474 => x"FF",
		52475 => x"FF",
		52476 => x"FF",
		52477 => x"FF",
		52478 => x"FF",
		52479 => x"FF",
		52480 => x"FF",
		52481 => x"FF",
		52482 => x"FF",
		52483 => x"FF",
		52484 => x"FF",
		52485 => x"FF",
		52486 => x"FF",
		52487 => x"FF",
		52488 => x"FF",
		52489 => x"FF",
		52490 => x"FF",
		52491 => x"FF",
		52492 => x"FF",
		52493 => x"FF",
		52494 => x"FF",
		52495 => x"FF",
		52496 => x"FF",
		52497 => x"FF",
		52498 => x"FF",
		52499 => x"FF",
		52500 => x"FF",
		52501 => x"FF",
		52502 => x"FF",
		52503 => x"FF",
		52504 => x"FF",
		52505 => x"FF",
		52506 => x"FF",
		52507 => x"FF",
		52508 => x"FF",
		52509 => x"FF",
		52510 => x"FF",
		52511 => x"FF",
		52512 => x"FF",
		52513 => x"FF",
		52514 => x"FF",
		52515 => x"FF",
		52516 => x"FF",
		52517 => x"FF",
		52518 => x"FF",
		52519 => x"FF",
		52520 => x"FF",
		52521 => x"FF",
		52522 => x"FF",
		52523 => x"FF",
		52524 => x"FF",
		52525 => x"FF",
		52526 => x"FF",
		52527 => x"FF",
		52528 => x"FF",
		52529 => x"FF",
		52530 => x"FF",
		52531 => x"FF",
		52532 => x"FF",
		52533 => x"FF",
		52534 => x"FF",
		52535 => x"FF",
		52536 => x"FF",
		52537 => x"FF",
		52538 => x"FF",
		52539 => x"FF",
		52540 => x"FF",
		52541 => x"FF",
		52542 => x"FF",
		52543 => x"FF",
		52544 => x"FF",
		52545 => x"FF",
		52546 => x"FF",
		52547 => x"FF",
		52548 => x"FF",
		52549 => x"FF",
		52550 => x"FF",
		52551 => x"FF",
		52552 => x"FF",
		52553 => x"FF",
		52554 => x"FF",
		52555 => x"FF",
		52556 => x"FF",
		52557 => x"FF",
		52558 => x"FF",
		52559 => x"FF",
		52560 => x"FF",
		52561 => x"FF",
		52562 => x"FF",
		52563 => x"FF",
		52564 => x"FF",
		52565 => x"FF",
		52566 => x"FF",
		52567 => x"FF",
		52568 => x"FF",
		52569 => x"FF",
		52570 => x"FF",
		52571 => x"FF",
		52572 => x"FF",
		52573 => x"FF",
		52574 => x"FF",
		52575 => x"FF",
		52576 => x"FF",
		52577 => x"FF",
		52578 => x"FF",
		52579 => x"FF",
		52580 => x"FF",
		52581 => x"FF",
		52582 => x"FF",
		52583 => x"FF",
		52584 => x"FF",
		52585 => x"FF",
		52586 => x"FF",
		52587 => x"FF",
		52588 => x"FF",
		52589 => x"FF",
		52590 => x"FF",
		52591 => x"FF",
		52592 => x"FF",
		52593 => x"FF",
		52594 => x"FF",
		52595 => x"FF",
		52596 => x"FF",
		52597 => x"FF",
		52598 => x"FF",
		52599 => x"FF",
		52600 => x"FF",
		52601 => x"FF",
		52602 => x"FF",
		52603 => x"FF",
		52604 => x"FF",
		52605 => x"FF",
		52606 => x"FF",
		52607 => x"FF",
		52608 => x"FF",
		52609 => x"FF",
		52610 => x"FF",
		52611 => x"FF",
		52612 => x"FF",
		52613 => x"FF",
		52614 => x"FF",
		52615 => x"FF",
		52616 => x"FF",
		52617 => x"FF",
		52618 => x"FF",
		52619 => x"FF",
		52620 => x"FF",
		52621 => x"FF",
		52622 => x"FF",
		52623 => x"FF",
		52624 => x"FF",
		52625 => x"FF",
		52626 => x"FF",
		52627 => x"FF",
		52628 => x"FF",
		52629 => x"FF",
		52630 => x"FF",
		52631 => x"FF",
		52632 => x"FF",
		52633 => x"FF",
		52634 => x"FF",
		52635 => x"FF",
		52636 => x"FF",
		52637 => x"FF",
		52638 => x"FF",
		52639 => x"FF",
		52640 => x"FF",
		52641 => x"FF",
		52642 => x"FF",
		52643 => x"FF",
		52644 => x"FF",
		52645 => x"FF",
		52646 => x"FF",
		52647 => x"FF",
		52648 => x"FF",
		52649 => x"FF",
		52650 => x"FF",
		52651 => x"FF",
		52652 => x"FF",
		52653 => x"FF",
		52654 => x"FF",
		52655 => x"FF",
		52656 => x"FF",
		52657 => x"FF",
		52658 => x"FF",
		52659 => x"FF",
		52660 => x"FF",
		52661 => x"FF",
		52662 => x"FF",
		52663 => x"FF",
		52664 => x"FF",
		52665 => x"FF",
		52666 => x"FF",
		52667 => x"FF",
		52668 => x"FF",
		52669 => x"FF",
		52670 => x"FF",
		52671 => x"FF",
		52672 => x"FF",
		52673 => x"FF",
		52674 => x"FF",
		52675 => x"FF",
		52676 => x"FF",
		52677 => x"FF",
		52678 => x"FF",
		52679 => x"FF",
		52680 => x"FF",
		52681 => x"FF",
		52682 => x"FF",
		52683 => x"FF",
		52684 => x"FF",
		52685 => x"FF",
		52686 => x"FF",
		52687 => x"FF",
		52688 => x"FF",
		52689 => x"FF",
		52690 => x"FF",
		52691 => x"FF",
		52692 => x"FF",
		52693 => x"FF",
		52694 => x"FF",
		52695 => x"FF",
		52696 => x"FF",
		52697 => x"FF",
		52698 => x"FF",
		52699 => x"FF",
		52700 => x"FF",
		52701 => x"FF",
		52702 => x"FF",
		52703 => x"FF",
		52704 => x"FF",
		52705 => x"FF",
		52706 => x"FF",
		52707 => x"FF",
		52708 => x"FF",
		52709 => x"FF",
		52710 => x"FF",
		52711 => x"FF",
		52712 => x"FF",
		52713 => x"FF",
		52714 => x"FF",
		52715 => x"FF",
		52716 => x"FF",
		52717 => x"FF",
		52718 => x"FF",
		52719 => x"FF",
		52720 => x"FF",
		52721 => x"FF",
		53366 => x"FF",
		53367 => x"FF",
		53368 => x"FF",
		53369 => x"FF",
		53370 => x"FF",
		53371 => x"FF",
		53372 => x"FF",
		53373 => x"FF",
		53374 => x"FF",
		53375 => x"FF",
		53376 => x"FF",
		53377 => x"FF",
		53378 => x"FF",
		53379 => x"FF",
		53380 => x"FF",
		53381 => x"FF",
		53382 => x"FF",
		53383 => x"FF",
		53384 => x"FF",
		53385 => x"FF",
		53386 => x"FF",
		53387 => x"FF",
		53388 => x"FF",
		53389 => x"FF",
		53390 => x"FF",
		53391 => x"FF",
		53392 => x"FF",
		53393 => x"FF",
		53394 => x"FF",
		53395 => x"FF",
		53396 => x"FF",
		53397 => x"FF",
		53398 => x"FF",
		53399 => x"FF",
		53400 => x"FF",
		53401 => x"FF",
		53402 => x"FF",
		53403 => x"FF",
		53404 => x"FF",
		53405 => x"FF",
		53406 => x"FF",
		53407 => x"FF",
		53408 => x"FF",
		53409 => x"FF",
		53410 => x"FF",
		53411 => x"FF",
		53412 => x"FF",
		53413 => x"FF",
		53414 => x"FF",
		53415 => x"FF",
		53416 => x"FF",
		53417 => x"FF",
		53418 => x"FF",
		53419 => x"FF",
		53420 => x"FF",
		53421 => x"FF",
		53422 => x"FF",
		53423 => x"FF",
		53424 => x"FF",
		53425 => x"FF",
		53426 => x"FF",
		53427 => x"FF",
		53428 => x"FF",
		53429 => x"FF",
		53430 => x"FF",
		53431 => x"FF",
		53432 => x"FF",
		53433 => x"FF",
		53434 => x"FF",
		53435 => x"FF",
		53436 => x"FF",
		53437 => x"FF",
		53438 => x"FF",
		53439 => x"FF",
		53440 => x"FF",
		53441 => x"FF",
		53442 => x"FF",
		53443 => x"FF",
		53444 => x"FF",
		53445 => x"FF",
		53446 => x"FF",
		53447 => x"FF",
		53448 => x"FF",
		53449 => x"FF",
		53450 => x"FF",
		53451 => x"FF",
		53452 => x"FF",
		53453 => x"FF",
		53454 => x"FF",
		53455 => x"FF",
		53456 => x"FF",
		53457 => x"FF",
		53458 => x"FF",
		53459 => x"FF",
		53460 => x"FF",
		53461 => x"FF",
		53462 => x"FF",
		53463 => x"FF",
		53464 => x"FF",
		53465 => x"FF",
		53466 => x"FF",
		53467 => x"FF",
		53468 => x"FF",
		53469 => x"FF",
		53470 => x"FF",
		53471 => x"FF",
		53472 => x"FF",
		53473 => x"FF",
		53474 => x"FF",
		53475 => x"FF",
		53476 => x"FF",
		53477 => x"FF",
		53478 => x"FF",
		53479 => x"FF",
		53480 => x"FF",
		53481 => x"FF",
		53482 => x"FF",
		53483 => x"FF",
		53484 => x"FF",
		53485 => x"FF",
		53486 => x"FF",
		53487 => x"FF",
		53488 => x"FF",
		53489 => x"FF",
		53490 => x"FF",
		53491 => x"FF",
		53492 => x"FF",
		53493 => x"FF",
		53494 => x"FF",
		53495 => x"FF",
		53496 => x"FF",
		53497 => x"FF",
		53498 => x"FF",
		53499 => x"FF",
		53500 => x"FF",
		53501 => x"FF",
		53502 => x"FF",
		53503 => x"FF",
		53504 => x"FF",
		53505 => x"FF",
		53506 => x"FF",
		53507 => x"FF",
		53508 => x"FF",
		53509 => x"FF",
		53510 => x"FF",
		53511 => x"FF",
		53512 => x"FF",
		53513 => x"FF",
		53514 => x"FF",
		53515 => x"FF",
		53516 => x"FF",
		53517 => x"FF",
		53518 => x"FF",
		53519 => x"FF",
		53520 => x"FF",
		53521 => x"FF",
		53522 => x"FF",
		53523 => x"FF",
		53524 => x"FF",
		53525 => x"FF",
		53526 => x"FF",
		53527 => x"FF",
		53528 => x"FF",
		53529 => x"FF",
		53530 => x"FF",
		53531 => x"FF",
		53532 => x"FF",
		53533 => x"FF",
		53534 => x"FF",
		53535 => x"FF",
		53536 => x"FF",
		53537 => x"FF",
		53538 => x"FF",
		53539 => x"FF",
		53540 => x"FF",
		53541 => x"FF",
		53542 => x"FF",
		53543 => x"FF",
		53544 => x"FF",
		53545 => x"FF",
		53546 => x"FF",
		53547 => x"FF",
		53548 => x"FF",
		53549 => x"FF",
		53550 => x"FF",
		53551 => x"FF",
		53552 => x"FF",
		53553 => x"FF",
		53554 => x"FF",
		53555 => x"FF",
		53556 => x"FF",
		53557 => x"FF",
		53558 => x"FF",
		53559 => x"FF",
		53560 => x"FF",
		53561 => x"FF",
		53562 => x"FF",
		53563 => x"FF",
		53564 => x"FF",
		53565 => x"FF",
		53566 => x"FF",
		53567 => x"FF",
		53568 => x"FF",
		53569 => x"FF",
		53570 => x"FF",
		53571 => x"FF",
		53572 => x"FF",
		53573 => x"FF",
		53574 => x"FF",
		53575 => x"FF",
		53576 => x"FF",
		53577 => x"FF",
		53578 => x"FF",
		53579 => x"FF",
		53580 => x"FF",
		53581 => x"FF",
		53582 => x"FF",
		53583 => x"FF",
		53584 => x"FF",
		53585 => x"FF",
		53586 => x"FF",
		53587 => x"FF",
		53588 => x"FF",
		53589 => x"FF",
		53590 => x"FF",
		53591 => x"FF",
		53592 => x"FF",
		53593 => x"FF",
		53594 => x"FF",
		53595 => x"FF",
		53596 => x"FF",
		53597 => x"FF",
		53598 => x"FF",
		53599 => x"FF",
		53600 => x"FF",
		53601 => x"FF",
		53602 => x"FF",
		53603 => x"FF",
		53604 => x"FF",
		53605 => x"FF",
		53606 => x"FF",
		53607 => x"FF",
		53608 => x"FF",
		53609 => x"FF",
		53610 => x"FF",
		53611 => x"FF",
		53612 => x"FF",
		53613 => x"FF",
		53614 => x"FF",
		53615 => x"FF",
		53616 => x"FF",
		53617 => x"FF",
		53618 => x"FF",
		53619 => x"FF",
		53620 => x"FF",
		53621 => x"FF",
		53622 => x"FF",
		53623 => x"FF",
		53624 => x"FF",
		53625 => x"FF",
		53626 => x"FF",
		53627 => x"FF",
		53628 => x"FF",
		53629 => x"FF",
		53630 => x"FF",
		53631 => x"FF",
		53632 => x"FF",
		53633 => x"FF",
		53634 => x"FF",
		53635 => x"FF",
		53636 => x"FF",
		53637 => x"FF",
		53638 => x"FF",
		53639 => x"FF",
		53640 => x"FF",
		53641 => x"FF",
		53642 => x"FF",
		53643 => x"FF",
		53644 => x"FF",
		53645 => x"FF",
		53646 => x"FF",
		53647 => x"FF",
		53648 => x"FF",
		53649 => x"FF",
		53650 => x"FF",
		53651 => x"FF",
		53652 => x"FF",
		53653 => x"FF",
		53654 => x"FF",
		53655 => x"FF",
		53656 => x"FF",
		53657 => x"FF",
		53658 => x"FF",
		53659 => x"FF",
		53660 => x"FF",
		53661 => x"FF",
		53662 => x"FF",
		53663 => x"FF",
		53664 => x"FF",
		53665 => x"FF",
		53666 => x"FF",
		53667 => x"FF",
		53668 => x"FF",
		53669 => x"FF",
		53670 => x"FF",
		53671 => x"FF",
		53672 => x"FF",
		53673 => x"FF",
		53674 => x"FF",
		53675 => x"FF",
		53676 => x"FF",
		53677 => x"FF",
		53678 => x"FF",
		53679 => x"FF",
		53680 => x"FF",
		53681 => x"FF",
		53682 => x"FF",
		53683 => x"FF",
		53684 => x"FF",
		53685 => x"FF",
		53686 => x"FF",
		53687 => x"FF",
		53688 => x"FF",
		53689 => x"FF",
		53690 => x"FF",
		53691 => x"FF",
		53692 => x"FF",
		53693 => x"FF",
		53694 => x"FF",
		53695 => x"FF",
		53696 => x"FF",
		53697 => x"FF",
		53698 => x"FF",
		53699 => x"FF",
		53700 => x"FF",
		53701 => x"FF",
		53702 => x"FF",
		53703 => x"FF",
		53704 => x"FF",
		53705 => x"FF",
		53706 => x"FF",
		53707 => x"FF",
		53708 => x"FF",
		53709 => x"FF",
		53710 => x"FF",
		53711 => x"FF",
		53712 => x"FF",
		53713 => x"FF",
		53714 => x"FF",
		53715 => x"FF",
		53716 => x"FF",
		53717 => x"FF",
		53718 => x"FF",
		53719 => x"FF",
		53720 => x"FF",
		53721 => x"FF",
		53722 => x"FF",
		53723 => x"FF",
		53724 => x"FF",
		53725 => x"FF",
		53726 => x"FF",
		53727 => x"FF",
		53728 => x"FF",
		53729 => x"FF",
		53730 => x"FF",
		53731 => x"FF",
		53732 => x"FF",
		53733 => x"FF",
		53734 => x"FF",
		53735 => x"FF",
		53736 => x"FF",
		53737 => x"FF",
		53738 => x"FF",
		53739 => x"FF",
		53740 => x"FF",
		53741 => x"FF",
		53742 => x"FF",
		53743 => x"FF",
		53744 => x"FF",
		53745 => x"FF",
		54390 => x"FF",
		54391 => x"FF",
		54392 => x"FF",
		54393 => x"FF",
		54394 => x"FF",
		54515 => x"FF",
		54516 => x"FF",
		54517 => x"FF",
		54518 => x"FF",
		54519 => x"FF",
		54640 => x"FF",
		54641 => x"FF",
		54642 => x"FF",
		54643 => x"FF",
		54644 => x"FF",
		54765 => x"FF",
		54766 => x"FF",
		54767 => x"FF",
		54768 => x"FF",
		54769 => x"FF",
		55414 => x"FF",
		55415 => x"FF",
		55416 => x"FF",
		55417 => x"FF",
		55418 => x"FF",
		55539 => x"FF",
		55540 => x"FF",
		55541 => x"FF",
		55542 => x"FF",
		55543 => x"FF",
		55664 => x"FF",
		55665 => x"FF",
		55666 => x"FF",
		55667 => x"FF",
		55668 => x"FF",
		55789 => x"FF",
		55790 => x"FF",
		55791 => x"FF",
		55792 => x"FF",
		55793 => x"FF",
		56438 => x"FF",
		56439 => x"FF",
		56440 => x"FF",
		56441 => x"FF",
		56442 => x"FF",
		56563 => x"FF",
		56564 => x"FF",
		56565 => x"FF",
		56566 => x"FF",
		56567 => x"FF",
		56688 => x"FF",
		56689 => x"FF",
		56690 => x"FF",
		56691 => x"FF",
		56692 => x"FF",
		56813 => x"FF",
		56814 => x"FF",
		56815 => x"FF",
		56816 => x"FF",
		56817 => x"FF",
		57462 => x"FF",
		57463 => x"FF",
		57464 => x"FF",
		57465 => x"FF",
		57466 => x"FF",
		57587 => x"FF",
		57588 => x"FF",
		57589 => x"FF",
		57590 => x"FF",
		57591 => x"FF",
		57712 => x"FF",
		57713 => x"FF",
		57714 => x"FF",
		57715 => x"FF",
		57716 => x"FF",
		57837 => x"FF",
		57838 => x"FF",
		57839 => x"FF",
		57840 => x"FF",
		57841 => x"FF",
		58486 => x"FF",
		58487 => x"FF",
		58488 => x"FF",
		58489 => x"FF",
		58490 => x"FF",
		58611 => x"FF",
		58612 => x"FF",
		58613 => x"FF",
		58614 => x"FF",
		58615 => x"FF",
		58736 => x"FF",
		58737 => x"FF",
		58738 => x"FF",
		58739 => x"FF",
		58740 => x"FF",
		58861 => x"FF",
		58862 => x"FF",
		58863 => x"FF",
		58864 => x"FF",
		58865 => x"FF",
		59510 => x"FF",
		59511 => x"FF",
		59512 => x"FF",
		59513 => x"FF",
		59514 => x"FF",
		59635 => x"FF",
		59636 => x"FF",
		59637 => x"FF",
		59638 => x"FF",
		59639 => x"FF",
		59760 => x"FF",
		59761 => x"FF",
		59762 => x"FF",
		59763 => x"FF",
		59764 => x"FF",
		59885 => x"FF",
		59886 => x"FF",
		59887 => x"FF",
		59888 => x"FF",
		59889 => x"FF",
		60534 => x"FF",
		60535 => x"FF",
		60536 => x"FF",
		60537 => x"FF",
		60538 => x"FF",
		60659 => x"FF",
		60660 => x"FF",
		60661 => x"FF",
		60662 => x"FF",
		60663 => x"FF",
		60784 => x"FF",
		60785 => x"FF",
		60786 => x"FF",
		60787 => x"FF",
		60788 => x"FF",
		60909 => x"FF",
		60910 => x"FF",
		60911 => x"FF",
		60912 => x"FF",
		60913 => x"FF",
		61558 => x"FF",
		61559 => x"FF",
		61560 => x"FF",
		61561 => x"FF",
		61562 => x"FF",
		61683 => x"FF",
		61684 => x"FF",
		61685 => x"FF",
		61686 => x"FF",
		61687 => x"FF",
		61808 => x"FF",
		61809 => x"FF",
		61810 => x"FF",
		61811 => x"FF",
		61812 => x"FF",
		61933 => x"FF",
		61934 => x"FF",
		61935 => x"FF",
		61936 => x"FF",
		61937 => x"FF",
		62582 => x"FF",
		62583 => x"FF",
		62584 => x"FF",
		62585 => x"FF",
		62586 => x"FF",
		62707 => x"FF",
		62708 => x"FF",
		62709 => x"FF",
		62710 => x"FF",
		62711 => x"FF",
		62832 => x"FF",
		62833 => x"FF",
		62834 => x"FF",
		62835 => x"FF",
		62836 => x"FF",
		62957 => x"FF",
		62958 => x"FF",
		62959 => x"FF",
		62960 => x"FF",
		62961 => x"FF",
		63606 => x"FF",
		63607 => x"FF",
		63608 => x"FF",
		63609 => x"FF",
		63610 => x"FF",
		63731 => x"FF",
		63732 => x"FF",
		63733 => x"FF",
		63734 => x"FF",
		63735 => x"FF",
		63856 => x"FF",
		63857 => x"FF",
		63858 => x"FF",
		63859 => x"FF",
		63860 => x"FF",
		63981 => x"FF",
		63982 => x"FF",
		63983 => x"FF",
		63984 => x"FF",
		63985 => x"FF",
		64630 => x"FF",
		64631 => x"FF",
		64632 => x"FF",
		64633 => x"FF",
		64634 => x"FF",
		64755 => x"FF",
		64756 => x"FF",
		64757 => x"FF",
		64758 => x"FF",
		64759 => x"FF",
		64880 => x"FF",
		64881 => x"FF",
		64882 => x"FF",
		64883 => x"FF",
		64884 => x"FF",
		65005 => x"FF",
		65006 => x"FF",
		65007 => x"FF",
		65008 => x"FF",
		65009 => x"FF",
		65654 => x"FF",
		65655 => x"FF",
		65656 => x"FF",
		65657 => x"FF",
		65658 => x"FF",
		65779 => x"FF",
		65780 => x"FF",
		65781 => x"FF",
		65782 => x"FF",
		65783 => x"FF",
		65904 => x"FF",
		65905 => x"FF",
		65906 => x"FF",
		65907 => x"FF",
		65908 => x"FF",
		66029 => x"FF",
		66030 => x"FF",
		66031 => x"FF",
		66032 => x"FF",
		66033 => x"FF",
		66678 => x"FF",
		66679 => x"FF",
		66680 => x"FF",
		66681 => x"FF",
		66682 => x"FF",
		66803 => x"FF",
		66804 => x"FF",
		66805 => x"FF",
		66806 => x"FF",
		66807 => x"FF",
		66928 => x"FF",
		66929 => x"FF",
		66930 => x"FF",
		66931 => x"FF",
		66932 => x"FF",
		67053 => x"FF",
		67054 => x"FF",
		67055 => x"FF",
		67056 => x"FF",
		67057 => x"FF",
		67702 => x"FF",
		67703 => x"FF",
		67704 => x"FF",
		67705 => x"FF",
		67706 => x"FF",
		67827 => x"FF",
		67828 => x"FF",
		67829 => x"FF",
		67830 => x"FF",
		67831 => x"FF",
		67952 => x"FF",
		67953 => x"FF",
		67954 => x"FF",
		67955 => x"FF",
		67956 => x"FF",
		68077 => x"FF",
		68078 => x"FF",
		68079 => x"FF",
		68080 => x"FF",
		68081 => x"FF",
		68726 => x"FF",
		68727 => x"FF",
		68728 => x"FF",
		68729 => x"FF",
		68730 => x"FF",
		68851 => x"FF",
		68852 => x"FF",
		68853 => x"FF",
		68854 => x"FF",
		68855 => x"FF",
		68976 => x"FF",
		68977 => x"FF",
		68978 => x"FF",
		68979 => x"FF",
		68980 => x"FF",
		69101 => x"FF",
		69102 => x"FF",
		69103 => x"FF",
		69104 => x"FF",
		69105 => x"FF",
		69750 => x"FF",
		69751 => x"FF",
		69752 => x"FF",
		69753 => x"FF",
		69754 => x"FF",
		69875 => x"FF",
		69876 => x"FF",
		69877 => x"FF",
		69878 => x"FF",
		69879 => x"FF",
		70000 => x"FF",
		70001 => x"FF",
		70002 => x"FF",
		70003 => x"FF",
		70004 => x"FF",
		70125 => x"FF",
		70126 => x"FF",
		70127 => x"FF",
		70128 => x"FF",
		70129 => x"FF",
		70774 => x"FF",
		70775 => x"FF",
		70776 => x"FF",
		70777 => x"FF",
		70778 => x"FF",
		70899 => x"FF",
		70900 => x"FF",
		70901 => x"FF",
		70902 => x"FF",
		70903 => x"FF",
		71024 => x"FF",
		71025 => x"FF",
		71026 => x"FF",
		71027 => x"FF",
		71028 => x"FF",
		71149 => x"FF",
		71150 => x"FF",
		71151 => x"FF",
		71152 => x"FF",
		71153 => x"FF",
		71798 => x"FF",
		71799 => x"FF",
		71800 => x"FF",
		71801 => x"FF",
		71802 => x"FF",
		71923 => x"FF",
		71924 => x"FF",
		71925 => x"FF",
		71926 => x"FF",
		71927 => x"FF",
		72048 => x"FF",
		72049 => x"FF",
		72050 => x"FF",
		72051 => x"FF",
		72052 => x"FF",
		72173 => x"FF",
		72174 => x"FF",
		72175 => x"FF",
		72176 => x"FF",
		72177 => x"FF",
		72822 => x"FF",
		72823 => x"FF",
		72824 => x"FF",
		72825 => x"FF",
		72826 => x"FF",
		72947 => x"FF",
		72948 => x"FF",
		72949 => x"FF",
		72950 => x"FF",
		72951 => x"FF",
		73072 => x"FF",
		73073 => x"FF",
		73074 => x"FF",
		73075 => x"FF",
		73076 => x"FF",
		73197 => x"FF",
		73198 => x"FF",
		73199 => x"FF",
		73200 => x"FF",
		73201 => x"FF",
		73846 => x"FF",
		73847 => x"FF",
		73848 => x"FF",
		73849 => x"FF",
		73850 => x"FF",
		73971 => x"FF",
		73972 => x"FF",
		73973 => x"FF",
		73974 => x"FF",
		73975 => x"FF",
		74096 => x"FF",
		74097 => x"FF",
		74098 => x"FF",
		74099 => x"FF",
		74100 => x"FF",
		74221 => x"FF",
		74222 => x"FF",
		74223 => x"FF",
		74224 => x"FF",
		74225 => x"FF",
		74870 => x"FF",
		74871 => x"FF",
		74872 => x"FF",
		74873 => x"FF",
		74874 => x"FF",
		74995 => x"FF",
		74996 => x"FF",
		74997 => x"FF",
		74998 => x"FF",
		74999 => x"FF",
		75120 => x"FF",
		75121 => x"FF",
		75122 => x"FF",
		75123 => x"FF",
		75124 => x"FF",
		75245 => x"FF",
		75246 => x"FF",
		75247 => x"FF",
		75248 => x"FF",
		75249 => x"FF",
		75894 => x"FF",
		75895 => x"FF",
		75896 => x"FF",
		75897 => x"FF",
		75898 => x"FF",
		76019 => x"FF",
		76020 => x"FF",
		76021 => x"FF",
		76022 => x"FF",
		76023 => x"FF",
		76144 => x"FF",
		76145 => x"FF",
		76146 => x"FF",
		76147 => x"FF",
		76148 => x"FF",
		76269 => x"FF",
		76270 => x"FF",
		76271 => x"FF",
		76272 => x"FF",
		76273 => x"FF",
		76918 => x"FF",
		76919 => x"FF",
		76920 => x"FF",
		76921 => x"FF",
		76922 => x"FF",
		77043 => x"FF",
		77044 => x"FF",
		77045 => x"FF",
		77046 => x"FF",
		77047 => x"FF",
		77168 => x"FF",
		77169 => x"FF",
		77170 => x"FF",
		77171 => x"FF",
		77172 => x"FF",
		77293 => x"FF",
		77294 => x"FF",
		77295 => x"FF",
		77296 => x"FF",
		77297 => x"FF",
		77942 => x"FF",
		77943 => x"FF",
		77944 => x"FF",
		77945 => x"FF",
		77946 => x"FF",
		78067 => x"FF",
		78068 => x"FF",
		78069 => x"FF",
		78070 => x"FF",
		78071 => x"FF",
		78192 => x"FF",
		78193 => x"FF",
		78194 => x"FF",
		78195 => x"FF",
		78196 => x"FF",
		78317 => x"FF",
		78318 => x"FF",
		78319 => x"FF",
		78320 => x"FF",
		78321 => x"FF",
		78966 => x"FF",
		78967 => x"FF",
		78968 => x"FF",
		78969 => x"FF",
		78970 => x"FF",
		79091 => x"FF",
		79092 => x"FF",
		79093 => x"FF",
		79094 => x"FF",
		79095 => x"FF",
		79216 => x"FF",
		79217 => x"FF",
		79218 => x"FF",
		79219 => x"FF",
		79220 => x"FF",
		79341 => x"FF",
		79342 => x"FF",
		79343 => x"FF",
		79344 => x"FF",
		79345 => x"FF",
		79990 => x"FF",
		79991 => x"FF",
		79992 => x"FF",
		79993 => x"FF",
		79994 => x"FF",
		80115 => x"FF",
		80116 => x"FF",
		80117 => x"FF",
		80118 => x"FF",
		80119 => x"FF",
		80240 => x"FF",
		80241 => x"FF",
		80242 => x"FF",
		80243 => x"FF",
		80244 => x"FF",
		80365 => x"FF",
		80366 => x"FF",
		80367 => x"FF",
		80368 => x"FF",
		80369 => x"FF",
		81014 => x"FF",
		81015 => x"FF",
		81016 => x"FF",
		81017 => x"FF",
		81018 => x"FF",
		81139 => x"FF",
		81140 => x"FF",
		81141 => x"FF",
		81142 => x"FF",
		81143 => x"FF",
		81264 => x"FF",
		81265 => x"FF",
		81266 => x"FF",
		81267 => x"FF",
		81268 => x"FF",
		81389 => x"FF",
		81390 => x"FF",
		81391 => x"FF",
		81392 => x"FF",
		81393 => x"FF",
		82038 => x"FF",
		82039 => x"FF",
		82040 => x"FF",
		82041 => x"FF",
		82042 => x"FF",
		82163 => x"FF",
		82164 => x"FF",
		82165 => x"FF",
		82166 => x"FF",
		82167 => x"FF",
		82288 => x"FF",
		82289 => x"FF",
		82290 => x"FF",
		82291 => x"FF",
		82292 => x"FF",
		82413 => x"FF",
		82414 => x"FF",
		82415 => x"FF",
		82416 => x"FF",
		82417 => x"FF",
		83062 => x"FF",
		83063 => x"FF",
		83064 => x"FF",
		83065 => x"FF",
		83066 => x"FF",
		83187 => x"FF",
		83188 => x"FF",
		83189 => x"FF",
		83190 => x"FF",
		83191 => x"FF",
		83312 => x"FF",
		83313 => x"FF",
		83314 => x"FF",
		83315 => x"FF",
		83316 => x"FF",
		83437 => x"FF",
		83438 => x"FF",
		83439 => x"FF",
		83440 => x"FF",
		83441 => x"FF",
		84086 => x"FF",
		84087 => x"FF",
		84088 => x"FF",
		84089 => x"FF",
		84090 => x"FF",
		84211 => x"FF",
		84212 => x"FF",
		84213 => x"FF",
		84214 => x"FF",
		84215 => x"FF",
		84336 => x"FF",
		84337 => x"FF",
		84338 => x"FF",
		84339 => x"FF",
		84340 => x"FF",
		84461 => x"FF",
		84462 => x"FF",
		84463 => x"FF",
		84464 => x"FF",
		84465 => x"FF",
		85110 => x"FF",
		85111 => x"FF",
		85112 => x"FF",
		85113 => x"FF",
		85114 => x"FF",
		85235 => x"FF",
		85236 => x"FF",
		85237 => x"FF",
		85238 => x"FF",
		85239 => x"FF",
		85360 => x"FF",
		85361 => x"FF",
		85362 => x"FF",
		85363 => x"FF",
		85364 => x"FF",
		85485 => x"FF",
		85486 => x"FF",
		85487 => x"FF",
		85488 => x"FF",
		85489 => x"FF",
		86134 => x"FF",
		86135 => x"FF",
		86136 => x"FF",
		86137 => x"FF",
		86138 => x"FF",
		86259 => x"FF",
		86260 => x"FF",
		86261 => x"FF",
		86262 => x"FF",
		86263 => x"FF",
		86384 => x"FF",
		86385 => x"FF",
		86386 => x"FF",
		86387 => x"FF",
		86388 => x"FF",
		86509 => x"FF",
		86510 => x"FF",
		86511 => x"FF",
		86512 => x"FF",
		86513 => x"FF",
		87158 => x"FF",
		87159 => x"FF",
		87160 => x"FF",
		87161 => x"FF",
		87162 => x"FF",
		87283 => x"FF",
		87284 => x"FF",
		87285 => x"FF",
		87286 => x"FF",
		87287 => x"FF",
		87408 => x"FF",
		87409 => x"FF",
		87410 => x"FF",
		87411 => x"FF",
		87412 => x"FF",
		87533 => x"FF",
		87534 => x"FF",
		87535 => x"FF",
		87536 => x"FF",
		87537 => x"FF",
		88182 => x"FF",
		88183 => x"FF",
		88184 => x"FF",
		88185 => x"FF",
		88186 => x"FF",
		88307 => x"FF",
		88308 => x"FF",
		88309 => x"FF",
		88310 => x"FF",
		88311 => x"FF",
		88432 => x"FF",
		88433 => x"FF",
		88434 => x"FF",
		88435 => x"FF",
		88436 => x"FF",
		88557 => x"FF",
		88558 => x"FF",
		88559 => x"FF",
		88560 => x"FF",
		88561 => x"FF",
		89206 => x"FF",
		89207 => x"FF",
		89208 => x"FF",
		89209 => x"FF",
		89210 => x"FF",
		89331 => x"FF",
		89332 => x"FF",
		89333 => x"FF",
		89334 => x"FF",
		89335 => x"FF",
		89456 => x"FF",
		89457 => x"FF",
		89458 => x"FF",
		89459 => x"FF",
		89460 => x"FF",
		89581 => x"FF",
		89582 => x"FF",
		89583 => x"FF",
		89584 => x"FF",
		89585 => x"FF",
		90230 => x"FF",
		90231 => x"FF",
		90232 => x"FF",
		90233 => x"FF",
		90234 => x"FF",
		90355 => x"FF",
		90356 => x"FF",
		90357 => x"FF",
		90358 => x"FF",
		90359 => x"FF",
		90480 => x"FF",
		90481 => x"FF",
		90482 => x"FF",
		90483 => x"FF",
		90484 => x"FF",
		90605 => x"FF",
		90606 => x"FF",
		90607 => x"FF",
		90608 => x"FF",
		90609 => x"FF",
		91254 => x"FF",
		91255 => x"FF",
		91256 => x"FF",
		91257 => x"FF",
		91258 => x"FF",
		91379 => x"FF",
		91380 => x"FF",
		91381 => x"FF",
		91382 => x"FF",
		91383 => x"FF",
		91504 => x"FF",
		91505 => x"FF",
		91506 => x"FF",
		91507 => x"FF",
		91508 => x"FF",
		91629 => x"FF",
		91630 => x"FF",
		91631 => x"FF",
		91632 => x"FF",
		91633 => x"FF",
		92278 => x"FF",
		92279 => x"FF",
		92280 => x"FF",
		92281 => x"FF",
		92282 => x"FF",
		92403 => x"FF",
		92404 => x"FF",
		92405 => x"FF",
		92406 => x"FF",
		92407 => x"FF",
		92528 => x"FF",
		92529 => x"FF",
		92530 => x"FF",
		92531 => x"FF",
		92532 => x"FF",
		92653 => x"FF",
		92654 => x"FF",
		92655 => x"FF",
		92656 => x"FF",
		92657 => x"FF",
		93302 => x"FF",
		93303 => x"FF",
		93304 => x"FF",
		93305 => x"FF",
		93306 => x"FF",
		93427 => x"FF",
		93428 => x"FF",
		93429 => x"FF",
		93430 => x"FF",
		93431 => x"FF",
		93552 => x"FF",
		93553 => x"FF",
		93554 => x"FF",
		93555 => x"FF",
		93556 => x"FF",
		93677 => x"FF",
		93678 => x"FF",
		93679 => x"FF",
		93680 => x"FF",
		93681 => x"FF",
		94326 => x"FF",
		94327 => x"FF",
		94328 => x"FF",
		94329 => x"FF",
		94330 => x"FF",
		94451 => x"FF",
		94452 => x"FF",
		94453 => x"FF",
		94454 => x"FF",
		94455 => x"FF",
		94576 => x"FF",
		94577 => x"FF",
		94578 => x"FF",
		94579 => x"FF",
		94580 => x"FF",
		94701 => x"FF",
		94702 => x"FF",
		94703 => x"FF",
		94704 => x"FF",
		94705 => x"FF",
		95350 => x"FF",
		95351 => x"FF",
		95352 => x"FF",
		95353 => x"FF",
		95354 => x"FF",
		95475 => x"FF",
		95476 => x"FF",
		95477 => x"FF",
		95478 => x"FF",
		95479 => x"FF",
		95600 => x"FF",
		95601 => x"FF",
		95602 => x"FF",
		95603 => x"FF",
		95604 => x"FF",
		95725 => x"FF",
		95726 => x"FF",
		95727 => x"FF",
		95728 => x"FF",
		95729 => x"FF",
		96374 => x"FF",
		96375 => x"FF",
		96376 => x"FF",
		96377 => x"FF",
		96378 => x"FF",
		96499 => x"FF",
		96500 => x"FF",
		96501 => x"FF",
		96502 => x"FF",
		96503 => x"FF",
		96624 => x"FF",
		96625 => x"FF",
		96626 => x"FF",
		96627 => x"FF",
		96628 => x"FF",
		96749 => x"FF",
		96750 => x"FF",
		96751 => x"FF",
		96752 => x"FF",
		96753 => x"FF",
		97398 => x"FF",
		97399 => x"FF",
		97400 => x"FF",
		97401 => x"FF",
		97402 => x"FF",
		97523 => x"FF",
		97524 => x"FF",
		97525 => x"FF",
		97526 => x"FF",
		97527 => x"FF",
		97648 => x"FF",
		97649 => x"FF",
		97650 => x"FF",
		97651 => x"FF",
		97652 => x"FF",
		97773 => x"FF",
		97774 => x"FF",
		97775 => x"FF",
		97776 => x"FF",
		97777 => x"FF",
		98422 => x"FF",
		98423 => x"FF",
		98424 => x"FF",
		98425 => x"FF",
		98426 => x"FF",
		98547 => x"FF",
		98548 => x"FF",
		98549 => x"FF",
		98550 => x"FF",
		98551 => x"FF",
		98672 => x"FF",
		98673 => x"FF",
		98674 => x"FF",
		98675 => x"FF",
		98676 => x"FF",
		98797 => x"FF",
		98798 => x"FF",
		98799 => x"FF",
		98800 => x"FF",
		98801 => x"FF",
		99446 => x"FF",
		99447 => x"FF",
		99448 => x"FF",
		99449 => x"FF",
		99450 => x"FF",
		99571 => x"FF",
		99572 => x"FF",
		99573 => x"FF",
		99574 => x"FF",
		99575 => x"FF",
		99696 => x"FF",
		99697 => x"FF",
		99698 => x"FF",
		99699 => x"FF",
		99700 => x"FF",
		99821 => x"FF",
		99822 => x"FF",
		99823 => x"FF",
		99824 => x"FF",
		99825 => x"FF",
		100470 => x"FF",
		100471 => x"FF",
		100472 => x"FF",
		100473 => x"FF",
		100474 => x"FF",
		100595 => x"FF",
		100596 => x"FF",
		100597 => x"FF",
		100598 => x"FF",
		100599 => x"FF",
		100720 => x"FF",
		100721 => x"FF",
		100722 => x"FF",
		100723 => x"FF",
		100724 => x"FF",
		100845 => x"FF",
		100846 => x"FF",
		100847 => x"FF",
		100848 => x"FF",
		100849 => x"FF",
		101494 => x"FF",
		101495 => x"FF",
		101496 => x"FF",
		101497 => x"FF",
		101498 => x"FF",
		101619 => x"FF",
		101620 => x"FF",
		101621 => x"FF",
		101622 => x"FF",
		101623 => x"FF",
		101744 => x"FF",
		101745 => x"FF",
		101746 => x"FF",
		101747 => x"FF",
		101748 => x"FF",
		101869 => x"FF",
		101870 => x"FF",
		101871 => x"FF",
		101872 => x"FF",
		101873 => x"FF",
		102518 => x"FF",
		102519 => x"FF",
		102520 => x"FF",
		102521 => x"FF",
		102522 => x"FF",
		102643 => x"FF",
		102644 => x"FF",
		102645 => x"FF",
		102646 => x"FF",
		102647 => x"FF",
		102768 => x"FF",
		102769 => x"FF",
		102770 => x"FF",
		102771 => x"FF",
		102772 => x"FF",
		102893 => x"FF",
		102894 => x"FF",
		102895 => x"FF",
		102896 => x"FF",
		102897 => x"FF",
		103542 => x"FF",
		103543 => x"FF",
		103544 => x"FF",
		103545 => x"FF",
		103546 => x"FF",
		103667 => x"FF",
		103668 => x"FF",
		103669 => x"FF",
		103670 => x"FF",
		103671 => x"FF",
		103792 => x"FF",
		103793 => x"FF",
		103794 => x"FF",
		103795 => x"FF",
		103796 => x"FF",
		103917 => x"FF",
		103918 => x"FF",
		103919 => x"FF",
		103920 => x"FF",
		103921 => x"FF",
		104566 => x"FF",
		104567 => x"FF",
		104568 => x"FF",
		104569 => x"FF",
		104570 => x"FF",
		104691 => x"FF",
		104692 => x"FF",
		104693 => x"FF",
		104694 => x"FF",
		104695 => x"FF",
		104816 => x"FF",
		104817 => x"FF",
		104818 => x"FF",
		104819 => x"FF",
		104820 => x"FF",
		104941 => x"FF",
		104942 => x"FF",
		104943 => x"FF",
		104944 => x"FF",
		104945 => x"FF",
		105590 => x"FF",
		105591 => x"FF",
		105592 => x"FF",
		105593 => x"FF",
		105594 => x"FF",
		105715 => x"FF",
		105716 => x"FF",
		105717 => x"FF",
		105718 => x"FF",
		105719 => x"FF",
		105840 => x"FF",
		105841 => x"FF",
		105842 => x"FF",
		105843 => x"FF",
		105844 => x"FF",
		105965 => x"FF",
		105966 => x"FF",
		105967 => x"FF",
		105968 => x"FF",
		105969 => x"FF",
		106614 => x"FF",
		106615 => x"FF",
		106616 => x"FF",
		106617 => x"FF",
		106618 => x"FF",
		106739 => x"FF",
		106740 => x"FF",
		106741 => x"FF",
		106742 => x"FF",
		106743 => x"FF",
		106864 => x"FF",
		106865 => x"FF",
		106866 => x"FF",
		106867 => x"FF",
		106868 => x"FF",
		106989 => x"FF",
		106990 => x"FF",
		106991 => x"FF",
		106992 => x"FF",
		106993 => x"FF",
		107638 => x"FF",
		107639 => x"FF",
		107640 => x"FF",
		107641 => x"FF",
		107642 => x"FF",
		107763 => x"FF",
		107764 => x"FF",
		107765 => x"FF",
		107766 => x"FF",
		107767 => x"FF",
		107888 => x"FF",
		107889 => x"FF",
		107890 => x"FF",
		107891 => x"FF",
		107892 => x"FF",
		108013 => x"FF",
		108014 => x"FF",
		108015 => x"FF",
		108016 => x"FF",
		108017 => x"FF",
		108662 => x"FF",
		108663 => x"FF",
		108664 => x"FF",
		108665 => x"FF",
		108666 => x"FF",
		108787 => x"FF",
		108788 => x"FF",
		108789 => x"FF",
		108790 => x"FF",
		108791 => x"FF",
		108912 => x"FF",
		108913 => x"FF",
		108914 => x"FF",
		108915 => x"FF",
		108916 => x"FF",
		109037 => x"FF",
		109038 => x"FF",
		109039 => x"FF",
		109040 => x"FF",
		109041 => x"FF",
		109686 => x"FF",
		109687 => x"FF",
		109688 => x"FF",
		109689 => x"FF",
		109690 => x"FF",
		109811 => x"FF",
		109812 => x"FF",
		109813 => x"FF",
		109814 => x"FF",
		109815 => x"FF",
		109936 => x"FF",
		109937 => x"FF",
		109938 => x"FF",
		109939 => x"FF",
		109940 => x"FF",
		110061 => x"FF",
		110062 => x"FF",
		110063 => x"FF",
		110064 => x"FF",
		110065 => x"FF",
		110710 => x"FF",
		110711 => x"FF",
		110712 => x"FF",
		110713 => x"FF",
		110714 => x"FF",
		110835 => x"FF",
		110836 => x"FF",
		110837 => x"FF",
		110838 => x"FF",
		110839 => x"FF",
		110960 => x"FF",
		110961 => x"FF",
		110962 => x"FF",
		110963 => x"FF",
		110964 => x"FF",
		111085 => x"FF",
		111086 => x"FF",
		111087 => x"FF",
		111088 => x"FF",
		111089 => x"FF",
		111734 => x"FF",
		111735 => x"FF",
		111736 => x"FF",
		111737 => x"FF",
		111738 => x"FF",
		111859 => x"FF",
		111860 => x"FF",
		111861 => x"FF",
		111862 => x"FF",
		111863 => x"FF",
		111984 => x"FF",
		111985 => x"FF",
		111986 => x"FF",
		111987 => x"FF",
		111988 => x"FF",
		112109 => x"FF",
		112110 => x"FF",
		112111 => x"FF",
		112112 => x"FF",
		112113 => x"FF",
		112758 => x"FF",
		112759 => x"FF",
		112760 => x"FF",
		112761 => x"FF",
		112762 => x"FF",
		112883 => x"FF",
		112884 => x"FF",
		112885 => x"FF",
		112886 => x"FF",
		112887 => x"FF",
		113008 => x"FF",
		113009 => x"FF",
		113010 => x"FF",
		113011 => x"FF",
		113012 => x"FF",
		113133 => x"FF",
		113134 => x"FF",
		113135 => x"FF",
		113136 => x"FF",
		113137 => x"FF",
		113782 => x"FF",
		113783 => x"FF",
		113784 => x"FF",
		113785 => x"FF",
		113786 => x"FF",
		113907 => x"FF",
		113908 => x"FF",
		113909 => x"FF",
		113910 => x"FF",
		113911 => x"FF",
		114032 => x"FF",
		114033 => x"FF",
		114034 => x"FF",
		114035 => x"FF",
		114036 => x"FF",
		114157 => x"FF",
		114158 => x"FF",
		114159 => x"FF",
		114160 => x"FF",
		114161 => x"FF",
		114806 => x"FF",
		114807 => x"FF",
		114808 => x"FF",
		114809 => x"FF",
		114810 => x"FF",
		114931 => x"FF",
		114932 => x"FF",
		114933 => x"FF",
		114934 => x"FF",
		114935 => x"FF",
		115056 => x"FF",
		115057 => x"FF",
		115058 => x"FF",
		115059 => x"FF",
		115060 => x"FF",
		115181 => x"FF",
		115182 => x"FF",
		115183 => x"FF",
		115184 => x"FF",
		115185 => x"FF",
		115830 => x"FF",
		115831 => x"FF",
		115832 => x"FF",
		115833 => x"FF",
		115834 => x"FF",
		115955 => x"FF",
		115956 => x"FF",
		115957 => x"FF",
		115958 => x"FF",
		115959 => x"FF",
		116080 => x"FF",
		116081 => x"FF",
		116082 => x"FF",
		116083 => x"FF",
		116084 => x"FF",
		116205 => x"FF",
		116206 => x"FF",
		116207 => x"FF",
		116208 => x"FF",
		116209 => x"FF",
		116854 => x"FF",
		116855 => x"FF",
		116856 => x"FF",
		116857 => x"FF",
		116858 => x"FF",
		116979 => x"FF",
		116980 => x"FF",
		116981 => x"FF",
		116982 => x"FF",
		116983 => x"FF",
		117104 => x"FF",
		117105 => x"FF",
		117106 => x"FF",
		117107 => x"FF",
		117108 => x"FF",
		117229 => x"FF",
		117230 => x"FF",
		117231 => x"FF",
		117232 => x"FF",
		117233 => x"FF",
		117878 => x"FF",
		117879 => x"FF",
		117880 => x"FF",
		117881 => x"FF",
		117882 => x"FF",
		118003 => x"FF",
		118004 => x"FF",
		118005 => x"FF",
		118006 => x"FF",
		118007 => x"FF",
		118128 => x"FF",
		118129 => x"FF",
		118130 => x"FF",
		118131 => x"FF",
		118132 => x"FF",
		118253 => x"FF",
		118254 => x"FF",
		118255 => x"FF",
		118256 => x"FF",
		118257 => x"FF",
		118902 => x"FF",
		118903 => x"FF",
		118904 => x"FF",
		118905 => x"FF",
		118906 => x"FF",
		119027 => x"FF",
		119028 => x"FF",
		119029 => x"FF",
		119030 => x"FF",
		119031 => x"FF",
		119152 => x"FF",
		119153 => x"FF",
		119154 => x"FF",
		119155 => x"FF",
		119156 => x"FF",
		119277 => x"FF",
		119278 => x"FF",
		119279 => x"FF",
		119280 => x"FF",
		119281 => x"FF",
		119926 => x"FF",
		119927 => x"FF",
		119928 => x"FF",
		119929 => x"FF",
		119930 => x"FF",
		120051 => x"FF",
		120052 => x"FF",
		120053 => x"FF",
		120054 => x"FF",
		120055 => x"FF",
		120176 => x"FF",
		120177 => x"FF",
		120178 => x"FF",
		120179 => x"FF",
		120180 => x"FF",
		120301 => x"FF",
		120302 => x"FF",
		120303 => x"FF",
		120304 => x"FF",
		120305 => x"FF",
		120950 => x"FF",
		120951 => x"FF",
		120952 => x"FF",
		120953 => x"FF",
		120954 => x"FF",
		121075 => x"FF",
		121076 => x"FF",
		121077 => x"FF",
		121078 => x"FF",
		121079 => x"FF",
		121200 => x"FF",
		121201 => x"FF",
		121202 => x"FF",
		121203 => x"FF",
		121204 => x"FF",
		121325 => x"FF",
		121326 => x"FF",
		121327 => x"FF",
		121328 => x"FF",
		121329 => x"FF",
		121974 => x"FF",
		121975 => x"FF",
		121976 => x"FF",
		121977 => x"FF",
		121978 => x"FF",
		122099 => x"FF",
		122100 => x"FF",
		122101 => x"FF",
		122102 => x"FF",
		122103 => x"FF",
		122224 => x"FF",
		122225 => x"FF",
		122226 => x"FF",
		122227 => x"FF",
		122228 => x"FF",
		122349 => x"FF",
		122350 => x"FF",
		122351 => x"FF",
		122352 => x"FF",
		122353 => x"FF",
		122998 => x"FF",
		122999 => x"FF",
		123000 => x"FF",
		123001 => x"FF",
		123002 => x"FF",
		123123 => x"FF",
		123124 => x"FF",
		123125 => x"FF",
		123126 => x"FF",
		123127 => x"FF",
		123248 => x"FF",
		123249 => x"FF",
		123250 => x"FF",
		123251 => x"FF",
		123252 => x"FF",
		123373 => x"FF",
		123374 => x"FF",
		123375 => x"FF",
		123376 => x"FF",
		123377 => x"FF",
		124022 => x"FF",
		124023 => x"FF",
		124024 => x"FF",
		124025 => x"FF",
		124026 => x"FF",
		124147 => x"FF",
		124148 => x"FF",
		124149 => x"FF",
		124150 => x"FF",
		124151 => x"FF",
		124272 => x"FF",
		124273 => x"FF",
		124274 => x"FF",
		124275 => x"FF",
		124276 => x"FF",
		124397 => x"FF",
		124398 => x"FF",
		124399 => x"FF",
		124400 => x"FF",
		124401 => x"FF",
		125046 => x"FF",
		125047 => x"FF",
		125048 => x"FF",
		125049 => x"FF",
		125050 => x"FF",
		125171 => x"FF",
		125172 => x"FF",
		125173 => x"FF",
		125174 => x"FF",
		125175 => x"FF",
		125296 => x"FF",
		125297 => x"FF",
		125298 => x"FF",
		125299 => x"FF",
		125300 => x"FF",
		125421 => x"FF",
		125422 => x"FF",
		125423 => x"FF",
		125424 => x"FF",
		125425 => x"FF",
		126070 => x"FF",
		126071 => x"FF",
		126072 => x"FF",
		126073 => x"FF",
		126074 => x"FF",
		126195 => x"FF",
		126196 => x"FF",
		126197 => x"FF",
		126198 => x"FF",
		126199 => x"FF",
		126320 => x"FF",
		126321 => x"FF",
		126322 => x"FF",
		126323 => x"FF",
		126324 => x"FF",
		126445 => x"FF",
		126446 => x"FF",
		126447 => x"FF",
		126448 => x"FF",
		126449 => x"FF",
		127094 => x"FF",
		127095 => x"FF",
		127096 => x"FF",
		127097 => x"FF",
		127098 => x"FF",
		127219 => x"FF",
		127220 => x"FF",
		127221 => x"FF",
		127222 => x"FF",
		127223 => x"FF",
		127344 => x"FF",
		127345 => x"FF",
		127346 => x"FF",
		127347 => x"FF",
		127348 => x"FF",
		127469 => x"FF",
		127470 => x"FF",
		127471 => x"FF",
		127472 => x"FF",
		127473 => x"FF",
		128118 => x"FF",
		128119 => x"FF",
		128120 => x"FF",
		128121 => x"FF",
		128122 => x"FF",
		128243 => x"FF",
		128244 => x"FF",
		128245 => x"FF",
		128246 => x"FF",
		128247 => x"FF",
		128368 => x"FF",
		128369 => x"FF",
		128370 => x"FF",
		128371 => x"FF",
		128372 => x"FF",
		128493 => x"FF",
		128494 => x"FF",
		128495 => x"FF",
		128496 => x"FF",
		128497 => x"FF",
		129142 => x"FF",
		129143 => x"FF",
		129144 => x"FF",
		129145 => x"FF",
		129146 => x"FF",
		129267 => x"FF",
		129268 => x"FF",
		129269 => x"FF",
		129270 => x"FF",
		129271 => x"FF",
		129392 => x"FF",
		129393 => x"FF",
		129394 => x"FF",
		129395 => x"FF",
		129396 => x"FF",
		129517 => x"FF",
		129518 => x"FF",
		129519 => x"FF",
		129520 => x"FF",
		129521 => x"FF",
		130166 => x"FF",
		130167 => x"FF",
		130168 => x"FF",
		130169 => x"FF",
		130170 => x"FF",
		130291 => x"FF",
		130292 => x"FF",
		130293 => x"FF",
		130294 => x"FF",
		130295 => x"FF",
		130416 => x"FF",
		130417 => x"FF",
		130418 => x"FF",
		130419 => x"FF",
		130420 => x"FF",
		130541 => x"FF",
		130542 => x"FF",
		130543 => x"FF",
		130544 => x"FF",
		130545 => x"FF",
		131190 => x"FF",
		131191 => x"FF",
		131192 => x"FF",
		131193 => x"FF",
		131194 => x"FF",
		131315 => x"FF",
		131316 => x"FF",
		131317 => x"FF",
		131318 => x"FF",
		131319 => x"FF",
		131440 => x"FF",
		131441 => x"FF",
		131442 => x"FF",
		131443 => x"FF",
		131444 => x"FF",
		131565 => x"FF",
		131566 => x"FF",
		131567 => x"FF",
		131568 => x"FF",
		131569 => x"FF",
		132214 => x"FF",
		132215 => x"FF",
		132216 => x"FF",
		132217 => x"FF",
		132218 => x"FF",
		132339 => x"FF",
		132340 => x"FF",
		132341 => x"FF",
		132342 => x"FF",
		132343 => x"FF",
		132464 => x"FF",
		132465 => x"FF",
		132466 => x"FF",
		132467 => x"FF",
		132468 => x"FF",
		132589 => x"FF",
		132590 => x"FF",
		132591 => x"FF",
		132592 => x"FF",
		132593 => x"FF",
		133238 => x"FF",
		133239 => x"FF",
		133240 => x"FF",
		133241 => x"FF",
		133242 => x"FF",
		133363 => x"FF",
		133364 => x"FF",
		133365 => x"FF",
		133366 => x"FF",
		133367 => x"FF",
		133488 => x"FF",
		133489 => x"FF",
		133490 => x"FF",
		133491 => x"FF",
		133492 => x"FF",
		133613 => x"FF",
		133614 => x"FF",
		133615 => x"FF",
		133616 => x"FF",
		133617 => x"FF",
		134262 => x"FF",
		134263 => x"FF",
		134264 => x"FF",
		134265 => x"FF",
		134266 => x"FF",
		134387 => x"FF",
		134388 => x"FF",
		134389 => x"FF",
		134390 => x"FF",
		134391 => x"FF",
		134512 => x"FF",
		134513 => x"FF",
		134514 => x"FF",
		134515 => x"FF",
		134516 => x"FF",
		134637 => x"FF",
		134638 => x"FF",
		134639 => x"FF",
		134640 => x"FF",
		134641 => x"FF",
		135286 => x"FF",
		135287 => x"FF",
		135288 => x"FF",
		135289 => x"FF",
		135290 => x"FF",
		135411 => x"FF",
		135412 => x"FF",
		135413 => x"FF",
		135414 => x"FF",
		135415 => x"FF",
		135536 => x"FF",
		135537 => x"FF",
		135538 => x"FF",
		135539 => x"FF",
		135540 => x"FF",
		135661 => x"FF",
		135662 => x"FF",
		135663 => x"FF",
		135664 => x"FF",
		135665 => x"FF",
		136310 => x"FF",
		136311 => x"FF",
		136312 => x"FF",
		136313 => x"FF",
		136314 => x"FF",
		136435 => x"FF",
		136436 => x"FF",
		136437 => x"FF",
		136438 => x"FF",
		136439 => x"FF",
		136560 => x"FF",
		136561 => x"FF",
		136562 => x"FF",
		136563 => x"FF",
		136564 => x"FF",
		136685 => x"FF",
		136686 => x"FF",
		136687 => x"FF",
		136688 => x"FF",
		136689 => x"FF",
		137334 => x"FF",
		137335 => x"FF",
		137336 => x"FF",
		137337 => x"FF",
		137338 => x"FF",
		137459 => x"FF",
		137460 => x"FF",
		137461 => x"FF",
		137462 => x"FF",
		137463 => x"FF",
		137584 => x"FF",
		137585 => x"FF",
		137586 => x"FF",
		137587 => x"FF",
		137588 => x"FF",
		137709 => x"FF",
		137710 => x"FF",
		137711 => x"FF",
		137712 => x"FF",
		137713 => x"FF",
		138358 => x"FF",
		138359 => x"FF",
		138360 => x"FF",
		138361 => x"FF",
		138362 => x"FF",
		138483 => x"FF",
		138484 => x"FF",
		138485 => x"FF",
		138486 => x"FF",
		138487 => x"FF",
		138608 => x"FF",
		138609 => x"FF",
		138610 => x"FF",
		138611 => x"FF",
		138612 => x"FF",
		138733 => x"FF",
		138734 => x"FF",
		138735 => x"FF",
		138736 => x"FF",
		138737 => x"FF",
		139382 => x"FF",
		139383 => x"FF",
		139384 => x"FF",
		139385 => x"FF",
		139386 => x"FF",
		139507 => x"FF",
		139508 => x"FF",
		139509 => x"FF",
		139510 => x"FF",
		139511 => x"FF",
		139632 => x"FF",
		139633 => x"FF",
		139634 => x"FF",
		139635 => x"FF",
		139636 => x"FF",
		139757 => x"FF",
		139758 => x"FF",
		139759 => x"FF",
		139760 => x"FF",
		139761 => x"FF",
		140406 => x"FF",
		140407 => x"FF",
		140408 => x"FF",
		140409 => x"FF",
		140410 => x"FF",
		140531 => x"FF",
		140532 => x"FF",
		140533 => x"FF",
		140534 => x"FF",
		140535 => x"FF",
		140656 => x"FF",
		140657 => x"FF",
		140658 => x"FF",
		140659 => x"FF",
		140660 => x"FF",
		140781 => x"FF",
		140782 => x"FF",
		140783 => x"FF",
		140784 => x"FF",
		140785 => x"FF",
		141430 => x"FF",
		141431 => x"FF",
		141432 => x"FF",
		141433 => x"FF",
		141434 => x"FF",
		141555 => x"FF",
		141556 => x"FF",
		141557 => x"FF",
		141558 => x"FF",
		141559 => x"FF",
		141680 => x"FF",
		141681 => x"FF",
		141682 => x"FF",
		141683 => x"FF",
		141684 => x"FF",
		141805 => x"FF",
		141806 => x"FF",
		141807 => x"FF",
		141808 => x"FF",
		141809 => x"FF",
		142454 => x"FF",
		142455 => x"FF",
		142456 => x"FF",
		142457 => x"FF",
		142458 => x"FF",
		142579 => x"FF",
		142580 => x"FF",
		142581 => x"FF",
		142582 => x"FF",
		142583 => x"FF",
		142704 => x"FF",
		142705 => x"FF",
		142706 => x"FF",
		142707 => x"FF",
		142708 => x"FF",
		142829 => x"FF",
		142830 => x"FF",
		142831 => x"FF",
		142832 => x"FF",
		142833 => x"FF",
		143478 => x"FF",
		143479 => x"FF",
		143480 => x"FF",
		143481 => x"FF",
		143482 => x"FF",
		143603 => x"FF",
		143604 => x"FF",
		143605 => x"FF",
		143606 => x"FF",
		143607 => x"FF",
		143728 => x"FF",
		143729 => x"FF",
		143730 => x"FF",
		143731 => x"FF",
		143732 => x"FF",
		143853 => x"FF",
		143854 => x"FF",
		143855 => x"FF",
		143856 => x"FF",
		143857 => x"FF",
		144502 => x"FF",
		144503 => x"FF",
		144504 => x"FF",
		144505 => x"FF",
		144506 => x"FF",
		144627 => x"FF",
		144628 => x"FF",
		144629 => x"FF",
		144630 => x"FF",
		144631 => x"FF",
		144752 => x"FF",
		144753 => x"FF",
		144754 => x"FF",
		144755 => x"FF",
		144756 => x"FF",
		144877 => x"FF",
		144878 => x"FF",
		144879 => x"FF",
		144880 => x"FF",
		144881 => x"FF",
		145526 => x"FF",
		145527 => x"FF",
		145528 => x"FF",
		145529 => x"FF",
		145530 => x"FF",
		145651 => x"FF",
		145652 => x"FF",
		145653 => x"FF",
		145654 => x"FF",
		145655 => x"FF",
		145776 => x"FF",
		145777 => x"FF",
		145778 => x"FF",
		145779 => x"FF",
		145780 => x"FF",
		145901 => x"FF",
		145902 => x"FF",
		145903 => x"FF",
		145904 => x"FF",
		145905 => x"FF",
		146550 => x"FF",
		146551 => x"FF",
		146552 => x"FF",
		146553 => x"FF",
		146554 => x"FF",
		146675 => x"FF",
		146676 => x"FF",
		146677 => x"FF",
		146678 => x"FF",
		146679 => x"FF",
		146800 => x"FF",
		146801 => x"FF",
		146802 => x"FF",
		146803 => x"FF",
		146804 => x"FF",
		146925 => x"FF",
		146926 => x"FF",
		146927 => x"FF",
		146928 => x"FF",
		146929 => x"FF",
		147574 => x"FF",
		147575 => x"FF",
		147576 => x"FF",
		147577 => x"FF",
		147578 => x"FF",
		147699 => x"FF",
		147700 => x"FF",
		147701 => x"FF",
		147702 => x"FF",
		147703 => x"FF",
		147824 => x"FF",
		147825 => x"FF",
		147826 => x"FF",
		147827 => x"FF",
		147828 => x"FF",
		147949 => x"FF",
		147950 => x"FF",
		147951 => x"FF",
		147952 => x"FF",
		147953 => x"FF",
		148598 => x"FF",
		148599 => x"FF",
		148600 => x"FF",
		148601 => x"FF",
		148602 => x"FF",
		148723 => x"FF",
		148724 => x"FF",
		148725 => x"FF",
		148726 => x"FF",
		148727 => x"FF",
		148848 => x"FF",
		148849 => x"FF",
		148850 => x"FF",
		148851 => x"FF",
		148852 => x"FF",
		148973 => x"FF",
		148974 => x"FF",
		148975 => x"FF",
		148976 => x"FF",
		148977 => x"FF",
		149622 => x"FF",
		149623 => x"FF",
		149624 => x"FF",
		149625 => x"FF",
		149626 => x"FF",
		149747 => x"FF",
		149748 => x"FF",
		149749 => x"FF",
		149750 => x"FF",
		149751 => x"FF",
		149872 => x"FF",
		149873 => x"FF",
		149874 => x"FF",
		149875 => x"FF",
		149876 => x"FF",
		149997 => x"FF",
		149998 => x"FF",
		149999 => x"FF",
		150000 => x"FF",
		150001 => x"FF",
		150646 => x"FF",
		150647 => x"FF",
		150648 => x"FF",
		150649 => x"FF",
		150650 => x"FF",
		150771 => x"FF",
		150772 => x"FF",
		150773 => x"FF",
		150774 => x"FF",
		150775 => x"FF",
		150896 => x"FF",
		150897 => x"FF",
		150898 => x"FF",
		150899 => x"FF",
		150900 => x"FF",
		151021 => x"FF",
		151022 => x"FF",
		151023 => x"FF",
		151024 => x"FF",
		151025 => x"FF",
		151670 => x"FF",
		151671 => x"FF",
		151672 => x"FF",
		151673 => x"FF",
		151674 => x"FF",
		151795 => x"FF",
		151796 => x"FF",
		151797 => x"FF",
		151798 => x"FF",
		151799 => x"FF",
		151920 => x"FF",
		151921 => x"FF",
		151922 => x"FF",
		151923 => x"FF",
		151924 => x"FF",
		152045 => x"FF",
		152046 => x"FF",
		152047 => x"FF",
		152048 => x"FF",
		152049 => x"FF",
		152694 => x"FF",
		152695 => x"FF",
		152696 => x"FF",
		152697 => x"FF",
		152698 => x"FF",
		152819 => x"FF",
		152820 => x"FF",
		152821 => x"FF",
		152822 => x"FF",
		152823 => x"FF",
		152944 => x"FF",
		152945 => x"FF",
		152946 => x"FF",
		152947 => x"FF",
		152948 => x"FF",
		153069 => x"FF",
		153070 => x"FF",
		153071 => x"FF",
		153072 => x"FF",
		153073 => x"FF",
		153718 => x"FF",
		153719 => x"FF",
		153720 => x"FF",
		153721 => x"FF",
		153722 => x"FF",
		153843 => x"FF",
		153844 => x"FF",
		153845 => x"FF",
		153846 => x"FF",
		153847 => x"FF",
		153968 => x"FF",
		153969 => x"FF",
		153970 => x"FF",
		153971 => x"FF",
		153972 => x"FF",
		154093 => x"FF",
		154094 => x"FF",
		154095 => x"FF",
		154096 => x"FF",
		154097 => x"FF",
		154742 => x"FF",
		154743 => x"FF",
		154744 => x"FF",
		154745 => x"FF",
		154746 => x"FF",
		154867 => x"FF",
		154868 => x"FF",
		154869 => x"FF",
		154870 => x"FF",
		154871 => x"FF",
		154992 => x"FF",
		154993 => x"FF",
		154994 => x"FF",
		154995 => x"FF",
		154996 => x"FF",
		155117 => x"FF",
		155118 => x"FF",
		155119 => x"FF",
		155120 => x"FF",
		155121 => x"FF",
		155766 => x"FF",
		155767 => x"FF",
		155768 => x"FF",
		155769 => x"FF",
		155770 => x"FF",
		155891 => x"FF",
		155892 => x"FF",
		155893 => x"FF",
		155894 => x"FF",
		155895 => x"FF",
		156016 => x"FF",
		156017 => x"FF",
		156018 => x"FF",
		156019 => x"FF",
		156020 => x"FF",
		156141 => x"FF",
		156142 => x"FF",
		156143 => x"FF",
		156144 => x"FF",
		156145 => x"FF",
		156790 => x"FF",
		156791 => x"FF",
		156792 => x"FF",
		156793 => x"FF",
		156794 => x"FF",
		156915 => x"FF",
		156916 => x"FF",
		156917 => x"FF",
		156918 => x"FF",
		156919 => x"FF",
		157040 => x"FF",
		157041 => x"FF",
		157042 => x"FF",
		157043 => x"FF",
		157044 => x"FF",
		157165 => x"FF",
		157166 => x"FF",
		157167 => x"FF",
		157168 => x"FF",
		157169 => x"FF",
		157814 => x"FF",
		157815 => x"FF",
		157816 => x"FF",
		157817 => x"FF",
		157818 => x"FF",
		157939 => x"FF",
		157940 => x"FF",
		157941 => x"FF",
		157942 => x"FF",
		157943 => x"FF",
		158064 => x"FF",
		158065 => x"FF",
		158066 => x"FF",
		158067 => x"FF",
		158068 => x"FF",
		158189 => x"FF",
		158190 => x"FF",
		158191 => x"FF",
		158192 => x"FF",
		158193 => x"FF",
		158838 => x"FF",
		158839 => x"FF",
		158840 => x"FF",
		158841 => x"FF",
		158842 => x"FF",
		158963 => x"FF",
		158964 => x"FF",
		158965 => x"FF",
		158966 => x"FF",
		158967 => x"FF",
		159088 => x"FF",
		159089 => x"FF",
		159090 => x"FF",
		159091 => x"FF",
		159092 => x"FF",
		159213 => x"FF",
		159214 => x"FF",
		159215 => x"FF",
		159216 => x"FF",
		159217 => x"FF",
		159862 => x"FF",
		159863 => x"FF",
		159864 => x"FF",
		159865 => x"FF",
		159866 => x"FF",
		159987 => x"FF",
		159988 => x"FF",
		159989 => x"FF",
		159990 => x"FF",
		159991 => x"FF",
		160112 => x"FF",
		160113 => x"FF",
		160114 => x"FF",
		160115 => x"FF",
		160116 => x"FF",
		160237 => x"FF",
		160238 => x"FF",
		160239 => x"FF",
		160240 => x"FF",
		160241 => x"FF",
		160886 => x"FF",
		160887 => x"FF",
		160888 => x"FF",
		160889 => x"FF",
		160890 => x"FF",
		161011 => x"FF",
		161012 => x"FF",
		161013 => x"FF",
		161014 => x"FF",
		161015 => x"FF",
		161136 => x"FF",
		161137 => x"FF",
		161138 => x"FF",
		161139 => x"FF",
		161140 => x"FF",
		161261 => x"FF",
		161262 => x"FF",
		161263 => x"FF",
		161264 => x"FF",
		161265 => x"FF",
		161910 => x"FF",
		161911 => x"FF",
		161912 => x"FF",
		161913 => x"FF",
		161914 => x"FF",
		162035 => x"FF",
		162036 => x"FF",
		162037 => x"FF",
		162038 => x"FF",
		162039 => x"FF",
		162160 => x"FF",
		162161 => x"FF",
		162162 => x"FF",
		162163 => x"FF",
		162164 => x"FF",
		162285 => x"FF",
		162286 => x"FF",
		162287 => x"FF",
		162288 => x"FF",
		162289 => x"FF",
		162934 => x"FF",
		162935 => x"FF",
		162936 => x"FF",
		162937 => x"FF",
		162938 => x"FF",
		163059 => x"FF",
		163060 => x"FF",
		163061 => x"FF",
		163062 => x"FF",
		163063 => x"FF",
		163184 => x"FF",
		163185 => x"FF",
		163186 => x"FF",
		163187 => x"FF",
		163188 => x"FF",
		163309 => x"FF",
		163310 => x"FF",
		163311 => x"FF",
		163312 => x"FF",
		163313 => x"FF",
		163958 => x"FF",
		163959 => x"FF",
		163960 => x"FF",
		163961 => x"FF",
		163962 => x"FF",
		164083 => x"FF",
		164084 => x"FF",
		164085 => x"FF",
		164086 => x"FF",
		164087 => x"FF",
		164208 => x"FF",
		164209 => x"FF",
		164210 => x"FF",
		164211 => x"FF",
		164212 => x"FF",
		164333 => x"FF",
		164334 => x"FF",
		164335 => x"FF",
		164336 => x"FF",
		164337 => x"FF",
		164982 => x"FF",
		164983 => x"FF",
		164984 => x"FF",
		164985 => x"FF",
		164986 => x"FF",
		165107 => x"FF",
		165108 => x"FF",
		165109 => x"FF",
		165110 => x"FF",
		165111 => x"FF",
		165232 => x"FF",
		165233 => x"FF",
		165234 => x"FF",
		165235 => x"FF",
		165236 => x"FF",
		165357 => x"FF",
		165358 => x"FF",
		165359 => x"FF",
		165360 => x"FF",
		165361 => x"FF",
		166006 => x"FF",
		166007 => x"FF",
		166008 => x"FF",
		166009 => x"FF",
		166010 => x"FF",
		166131 => x"FF",
		166132 => x"FF",
		166133 => x"FF",
		166134 => x"FF",
		166135 => x"FF",
		166256 => x"FF",
		166257 => x"FF",
		166258 => x"FF",
		166259 => x"FF",
		166260 => x"FF",
		166381 => x"FF",
		166382 => x"FF",
		166383 => x"FF",
		166384 => x"FF",
		166385 => x"FF",
		167030 => x"FF",
		167031 => x"FF",
		167032 => x"FF",
		167033 => x"FF",
		167034 => x"FF",
		167155 => x"FF",
		167156 => x"FF",
		167157 => x"FF",
		167158 => x"FF",
		167159 => x"FF",
		167280 => x"FF",
		167281 => x"FF",
		167282 => x"FF",
		167283 => x"FF",
		167284 => x"FF",
		167405 => x"FF",
		167406 => x"FF",
		167407 => x"FF",
		167408 => x"FF",
		167409 => x"FF",
		168054 => x"FF",
		168055 => x"FF",
		168056 => x"FF",
		168057 => x"FF",
		168058 => x"FF",
		168179 => x"FF",
		168180 => x"FF",
		168181 => x"FF",
		168182 => x"FF",
		168183 => x"FF",
		168304 => x"FF",
		168305 => x"FF",
		168306 => x"FF",
		168307 => x"FF",
		168308 => x"FF",
		168429 => x"FF",
		168430 => x"FF",
		168431 => x"FF",
		168432 => x"FF",
		168433 => x"FF",
		169078 => x"FF",
		169079 => x"FF",
		169080 => x"FF",
		169081 => x"FF",
		169082 => x"FF",
		169203 => x"FF",
		169204 => x"FF",
		169205 => x"FF",
		169206 => x"FF",
		169207 => x"FF",
		169328 => x"FF",
		169329 => x"FF",
		169330 => x"FF",
		169331 => x"FF",
		169332 => x"FF",
		169453 => x"FF",
		169454 => x"FF",
		169455 => x"FF",
		169456 => x"FF",
		169457 => x"FF",
		170102 => x"FF",
		170103 => x"FF",
		170104 => x"FF",
		170105 => x"FF",
		170106 => x"FF",
		170227 => x"FF",
		170228 => x"FF",
		170229 => x"FF",
		170230 => x"FF",
		170231 => x"FF",
		170352 => x"FF",
		170353 => x"FF",
		170354 => x"FF",
		170355 => x"FF",
		170356 => x"FF",
		170477 => x"FF",
		170478 => x"FF",
		170479 => x"FF",
		170480 => x"FF",
		170481 => x"FF",
		171126 => x"FF",
		171127 => x"FF",
		171128 => x"FF",
		171129 => x"FF",
		171130 => x"FF",
		171251 => x"FF",
		171252 => x"FF",
		171253 => x"FF",
		171254 => x"FF",
		171255 => x"FF",
		171376 => x"FF",
		171377 => x"FF",
		171378 => x"FF",
		171379 => x"FF",
		171380 => x"FF",
		171501 => x"FF",
		171502 => x"FF",
		171503 => x"FF",
		171504 => x"FF",
		171505 => x"FF",
		172150 => x"FF",
		172151 => x"FF",
		172152 => x"FF",
		172153 => x"FF",
		172154 => x"FF",
		172275 => x"FF",
		172276 => x"FF",
		172277 => x"FF",
		172278 => x"FF",
		172279 => x"FF",
		172400 => x"FF",
		172401 => x"FF",
		172402 => x"FF",
		172403 => x"FF",
		172404 => x"FF",
		172525 => x"FF",
		172526 => x"FF",
		172527 => x"FF",
		172528 => x"FF",
		172529 => x"FF",
		173174 => x"FF",
		173175 => x"FF",
		173176 => x"FF",
		173177 => x"FF",
		173178 => x"FF",
		173299 => x"FF",
		173300 => x"FF",
		173301 => x"FF",
		173302 => x"FF",
		173303 => x"FF",
		173424 => x"FF",
		173425 => x"FF",
		173426 => x"FF",
		173427 => x"FF",
		173428 => x"FF",
		173549 => x"FF",
		173550 => x"FF",
		173551 => x"FF",
		173552 => x"FF",
		173553 => x"FF",
		174198 => x"FF",
		174199 => x"FF",
		174200 => x"FF",
		174201 => x"FF",
		174202 => x"FF",
		174323 => x"FF",
		174324 => x"FF",
		174325 => x"FF",
		174326 => x"FF",
		174327 => x"FF",
		174448 => x"FF",
		174449 => x"FF",
		174450 => x"FF",
		174451 => x"FF",
		174452 => x"FF",
		174573 => x"FF",
		174574 => x"FF",
		174575 => x"FF",
		174576 => x"FF",
		174577 => x"FF",
		175222 => x"FF",
		175223 => x"FF",
		175224 => x"FF",
		175225 => x"FF",
		175226 => x"FF",
		175347 => x"FF",
		175348 => x"FF",
		175349 => x"FF",
		175350 => x"FF",
		175351 => x"FF",
		175472 => x"FF",
		175473 => x"FF",
		175474 => x"FF",
		175475 => x"FF",
		175476 => x"FF",
		175597 => x"FF",
		175598 => x"FF",
		175599 => x"FF",
		175600 => x"FF",
		175601 => x"FF",
		176246 => x"FF",
		176247 => x"FF",
		176248 => x"FF",
		176249 => x"FF",
		176250 => x"FF",
		176371 => x"FF",
		176372 => x"FF",
		176373 => x"FF",
		176374 => x"FF",
		176375 => x"FF",
		176496 => x"FF",
		176497 => x"FF",
		176498 => x"FF",
		176499 => x"FF",
		176500 => x"FF",
		176621 => x"FF",
		176622 => x"FF",
		176623 => x"FF",
		176624 => x"FF",
		176625 => x"FF",
		177270 => x"FF",
		177271 => x"FF",
		177272 => x"FF",
		177273 => x"FF",
		177274 => x"FF",
		177275 => x"FF",
		177276 => x"FF",
		177277 => x"FF",
		177278 => x"FF",
		177279 => x"FF",
		177280 => x"FF",
		177281 => x"FF",
		177282 => x"FF",
		177283 => x"FF",
		177284 => x"FF",
		177285 => x"FF",
		177286 => x"FF",
		177287 => x"FF",
		177288 => x"FF",
		177289 => x"FF",
		177290 => x"FF",
		177291 => x"FF",
		177292 => x"FF",
		177293 => x"FF",
		177294 => x"FF",
		177295 => x"FF",
		177296 => x"FF",
		177297 => x"FF",
		177298 => x"FF",
		177299 => x"FF",
		177300 => x"FF",
		177301 => x"FF",
		177302 => x"FF",
		177303 => x"FF",
		177304 => x"FF",
		177305 => x"FF",
		177306 => x"FF",
		177307 => x"FF",
		177308 => x"FF",
		177309 => x"FF",
		177310 => x"FF",
		177311 => x"FF",
		177312 => x"FF",
		177313 => x"FF",
		177314 => x"FF",
		177315 => x"FF",
		177316 => x"FF",
		177317 => x"FF",
		177318 => x"FF",
		177319 => x"FF",
		177320 => x"FF",
		177321 => x"FF",
		177322 => x"FF",
		177323 => x"FF",
		177324 => x"FF",
		177325 => x"FF",
		177326 => x"FF",
		177327 => x"FF",
		177328 => x"FF",
		177329 => x"FF",
		177330 => x"FF",
		177331 => x"FF",
		177332 => x"FF",
		177333 => x"FF",
		177334 => x"FF",
		177335 => x"FF",
		177336 => x"FF",
		177337 => x"FF",
		177338 => x"FF",
		177339 => x"FF",
		177340 => x"FF",
		177341 => x"FF",
		177342 => x"FF",
		177343 => x"FF",
		177344 => x"FF",
		177345 => x"FF",
		177346 => x"FF",
		177347 => x"FF",
		177348 => x"FF",
		177349 => x"FF",
		177350 => x"FF",
		177351 => x"FF",
		177352 => x"FF",
		177353 => x"FF",
		177354 => x"FF",
		177355 => x"FF",
		177356 => x"FF",
		177357 => x"FF",
		177358 => x"FF",
		177359 => x"FF",
		177360 => x"FF",
		177361 => x"FF",
		177362 => x"FF",
		177363 => x"FF",
		177364 => x"FF",
		177365 => x"FF",
		177366 => x"FF",
		177367 => x"FF",
		177368 => x"FF",
		177369 => x"FF",
		177370 => x"FF",
		177371 => x"FF",
		177372 => x"FF",
		177373 => x"FF",
		177374 => x"FF",
		177375 => x"FF",
		177376 => x"FF",
		177377 => x"FF",
		177378 => x"FF",
		177379 => x"FF",
		177380 => x"FF",
		177381 => x"FF",
		177382 => x"FF",
		177383 => x"FF",
		177384 => x"FF",
		177385 => x"FF",
		177386 => x"FF",
		177387 => x"FF",
		177388 => x"FF",
		177389 => x"FF",
		177390 => x"FF",
		177391 => x"FF",
		177392 => x"FF",
		177393 => x"FF",
		177394 => x"FF",
		177395 => x"FF",
		177396 => x"FF",
		177397 => x"FF",
		177398 => x"FF",
		177399 => x"FF",
		177400 => x"FF",
		177401 => x"FF",
		177402 => x"FF",
		177403 => x"FF",
		177404 => x"FF",
		177405 => x"FF",
		177406 => x"FF",
		177407 => x"FF",
		177408 => x"FF",
		177409 => x"FF",
		177410 => x"FF",
		177411 => x"FF",
		177412 => x"FF",
		177413 => x"FF",
		177414 => x"FF",
		177415 => x"FF",
		177416 => x"FF",
		177417 => x"FF",
		177418 => x"FF",
		177419 => x"FF",
		177420 => x"FF",
		177421 => x"FF",
		177422 => x"FF",
		177423 => x"FF",
		177424 => x"FF",
		177425 => x"FF",
		177426 => x"FF",
		177427 => x"FF",
		177428 => x"FF",
		177429 => x"FF",
		177430 => x"FF",
		177431 => x"FF",
		177432 => x"FF",
		177433 => x"FF",
		177434 => x"FF",
		177435 => x"FF",
		177436 => x"FF",
		177437 => x"FF",
		177438 => x"FF",
		177439 => x"FF",
		177440 => x"FF",
		177441 => x"FF",
		177442 => x"FF",
		177443 => x"FF",
		177444 => x"FF",
		177445 => x"FF",
		177446 => x"FF",
		177447 => x"FF",
		177448 => x"FF",
		177449 => x"FF",
		177450 => x"FF",
		177451 => x"FF",
		177452 => x"FF",
		177453 => x"FF",
		177454 => x"FF",
		177455 => x"FF",
		177456 => x"FF",
		177457 => x"FF",
		177458 => x"FF",
		177459 => x"FF",
		177460 => x"FF",
		177461 => x"FF",
		177462 => x"FF",
		177463 => x"FF",
		177464 => x"FF",
		177465 => x"FF",
		177466 => x"FF",
		177467 => x"FF",
		177468 => x"FF",
		177469 => x"FF",
		177470 => x"FF",
		177471 => x"FF",
		177472 => x"FF",
		177473 => x"FF",
		177474 => x"FF",
		177475 => x"FF",
		177476 => x"FF",
		177477 => x"FF",
		177478 => x"FF",
		177479 => x"FF",
		177480 => x"FF",
		177481 => x"FF",
		177482 => x"FF",
		177483 => x"FF",
		177484 => x"FF",
		177485 => x"FF",
		177486 => x"FF",
		177487 => x"FF",
		177488 => x"FF",
		177489 => x"FF",
		177490 => x"FF",
		177491 => x"FF",
		177492 => x"FF",
		177493 => x"FF",
		177494 => x"FF",
		177495 => x"FF",
		177496 => x"FF",
		177497 => x"FF",
		177498 => x"FF",
		177499 => x"FF",
		177500 => x"FF",
		177501 => x"FF",
		177502 => x"FF",
		177503 => x"FF",
		177504 => x"FF",
		177505 => x"FF",
		177506 => x"FF",
		177507 => x"FF",
		177508 => x"FF",
		177509 => x"FF",
		177510 => x"FF",
		177511 => x"FF",
		177512 => x"FF",
		177513 => x"FF",
		177514 => x"FF",
		177515 => x"FF",
		177516 => x"FF",
		177517 => x"FF",
		177518 => x"FF",
		177519 => x"FF",
		177520 => x"FF",
		177521 => x"FF",
		177522 => x"FF",
		177523 => x"FF",
		177524 => x"FF",
		177525 => x"FF",
		177526 => x"FF",
		177527 => x"FF",
		177528 => x"FF",
		177529 => x"FF",
		177530 => x"FF",
		177531 => x"FF",
		177532 => x"FF",
		177533 => x"FF",
		177534 => x"FF",
		177535 => x"FF",
		177536 => x"FF",
		177537 => x"FF",
		177538 => x"FF",
		177539 => x"FF",
		177540 => x"FF",
		177541 => x"FF",
		177542 => x"FF",
		177543 => x"FF",
		177544 => x"FF",
		177545 => x"FF",
		177546 => x"FF",
		177547 => x"FF",
		177548 => x"FF",
		177549 => x"FF",
		177550 => x"FF",
		177551 => x"FF",
		177552 => x"FF",
		177553 => x"FF",
		177554 => x"FF",
		177555 => x"FF",
		177556 => x"FF",
		177557 => x"FF",
		177558 => x"FF",
		177559 => x"FF",
		177560 => x"FF",
		177561 => x"FF",
		177562 => x"FF",
		177563 => x"FF",
		177564 => x"FF",
		177565 => x"FF",
		177566 => x"FF",
		177567 => x"FF",
		177568 => x"FF",
		177569 => x"FF",
		177570 => x"FF",
		177571 => x"FF",
		177572 => x"FF",
		177573 => x"FF",
		177574 => x"FF",
		177575 => x"FF",
		177576 => x"FF",
		177577 => x"FF",
		177578 => x"FF",
		177579 => x"FF",
		177580 => x"FF",
		177581 => x"FF",
		177582 => x"FF",
		177583 => x"FF",
		177584 => x"FF",
		177585 => x"FF",
		177586 => x"FF",
		177587 => x"FF",
		177588 => x"FF",
		177589 => x"FF",
		177590 => x"FF",
		177591 => x"FF",
		177592 => x"FF",
		177593 => x"FF",
		177594 => x"FF",
		177595 => x"FF",
		177596 => x"FF",
		177597 => x"FF",
		177598 => x"FF",
		177599 => x"FF",
		177600 => x"FF",
		177601 => x"FF",
		177602 => x"FF",
		177603 => x"FF",
		177604 => x"FF",
		177605 => x"FF",
		177606 => x"FF",
		177607 => x"FF",
		177608 => x"FF",
		177609 => x"FF",
		177610 => x"FF",
		177611 => x"FF",
		177612 => x"FF",
		177613 => x"FF",
		177614 => x"FF",
		177615 => x"FF",
		177616 => x"FF",
		177617 => x"FF",
		177618 => x"FF",
		177619 => x"FF",
		177620 => x"FF",
		177621 => x"FF",
		177622 => x"FF",
		177623 => x"FF",
		177624 => x"FF",
		177625 => x"FF",
		177626 => x"FF",
		177627 => x"FF",
		177628 => x"FF",
		177629 => x"FF",
		177630 => x"FF",
		177631 => x"FF",
		177632 => x"FF",
		177633 => x"FF",
		177634 => x"FF",
		177635 => x"FF",
		177636 => x"FF",
		177637 => x"FF",
		177638 => x"FF",
		177639 => x"FF",
		177640 => x"FF",
		177641 => x"FF",
		177642 => x"FF",
		177643 => x"FF",
		177644 => x"FF",
		177645 => x"FF",
		177646 => x"FF",
		177647 => x"FF",
		177648 => x"FF",
		177649 => x"FF",
		178294 => x"FF",
		178295 => x"FF",
		178296 => x"FF",
		178297 => x"FF",
		178298 => x"FF",
		178299 => x"FF",
		178300 => x"FF",
		178301 => x"FF",
		178302 => x"FF",
		178303 => x"FF",
		178304 => x"FF",
		178305 => x"FF",
		178306 => x"FF",
		178307 => x"FF",
		178308 => x"FF",
		178309 => x"FF",
		178310 => x"FF",
		178311 => x"FF",
		178312 => x"FF",
		178313 => x"FF",
		178314 => x"FF",
		178315 => x"FF",
		178316 => x"FF",
		178317 => x"FF",
		178318 => x"FF",
		178319 => x"FF",
		178320 => x"FF",
		178321 => x"FF",
		178322 => x"FF",
		178323 => x"FF",
		178324 => x"FF",
		178325 => x"FF",
		178326 => x"FF",
		178327 => x"FF",
		178328 => x"FF",
		178329 => x"FF",
		178330 => x"FF",
		178331 => x"FF",
		178332 => x"FF",
		178333 => x"FF",
		178334 => x"FF",
		178335 => x"FF",
		178336 => x"FF",
		178337 => x"FF",
		178338 => x"FF",
		178339 => x"FF",
		178340 => x"FF",
		178341 => x"FF",
		178342 => x"FF",
		178343 => x"FF",
		178344 => x"FF",
		178345 => x"FF",
		178346 => x"FF",
		178347 => x"FF",
		178348 => x"FF",
		178349 => x"FF",
		178350 => x"FF",
		178351 => x"FF",
		178352 => x"FF",
		178353 => x"FF",
		178354 => x"FF",
		178355 => x"FF",
		178356 => x"FF",
		178357 => x"FF",
		178358 => x"FF",
		178359 => x"FF",
		178360 => x"FF",
		178361 => x"FF",
		178362 => x"FF",
		178363 => x"FF",
		178364 => x"FF",
		178365 => x"FF",
		178366 => x"FF",
		178367 => x"FF",
		178368 => x"FF",
		178369 => x"FF",
		178370 => x"FF",
		178371 => x"FF",
		178372 => x"FF",
		178373 => x"FF",
		178374 => x"FF",
		178375 => x"FF",
		178376 => x"FF",
		178377 => x"FF",
		178378 => x"FF",
		178379 => x"FF",
		178380 => x"FF",
		178381 => x"FF",
		178382 => x"FF",
		178383 => x"FF",
		178384 => x"FF",
		178385 => x"FF",
		178386 => x"FF",
		178387 => x"FF",
		178388 => x"FF",
		178389 => x"FF",
		178390 => x"FF",
		178391 => x"FF",
		178392 => x"FF",
		178393 => x"FF",
		178394 => x"FF",
		178395 => x"FF",
		178396 => x"FF",
		178397 => x"FF",
		178398 => x"FF",
		178399 => x"FF",
		178400 => x"FF",
		178401 => x"FF",
		178402 => x"FF",
		178403 => x"FF",
		178404 => x"FF",
		178405 => x"FF",
		178406 => x"FF",
		178407 => x"FF",
		178408 => x"FF",
		178409 => x"FF",
		178410 => x"FF",
		178411 => x"FF",
		178412 => x"FF",
		178413 => x"FF",
		178414 => x"FF",
		178415 => x"FF",
		178416 => x"FF",
		178417 => x"FF",
		178418 => x"FF",
		178419 => x"FF",
		178420 => x"FF",
		178421 => x"FF",
		178422 => x"FF",
		178423 => x"FF",
		178424 => x"FF",
		178425 => x"FF",
		178426 => x"FF",
		178427 => x"FF",
		178428 => x"FF",
		178429 => x"FF",
		178430 => x"FF",
		178431 => x"FF",
		178432 => x"FF",
		178433 => x"FF",
		178434 => x"FF",
		178435 => x"FF",
		178436 => x"FF",
		178437 => x"FF",
		178438 => x"FF",
		178439 => x"FF",
		178440 => x"FF",
		178441 => x"FF",
		178442 => x"FF",
		178443 => x"FF",
		178444 => x"FF",
		178445 => x"FF",
		178446 => x"FF",
		178447 => x"FF",
		178448 => x"FF",
		178449 => x"FF",
		178450 => x"FF",
		178451 => x"FF",
		178452 => x"FF",
		178453 => x"FF",
		178454 => x"FF",
		178455 => x"FF",
		178456 => x"FF",
		178457 => x"FF",
		178458 => x"FF",
		178459 => x"FF",
		178460 => x"FF",
		178461 => x"FF",
		178462 => x"FF",
		178463 => x"FF",
		178464 => x"FF",
		178465 => x"FF",
		178466 => x"FF",
		178467 => x"FF",
		178468 => x"FF",
		178469 => x"FF",
		178470 => x"FF",
		178471 => x"FF",
		178472 => x"FF",
		178473 => x"FF",
		178474 => x"FF",
		178475 => x"FF",
		178476 => x"FF",
		178477 => x"FF",
		178478 => x"FF",
		178479 => x"FF",
		178480 => x"FF",
		178481 => x"FF",
		178482 => x"FF",
		178483 => x"FF",
		178484 => x"FF",
		178485 => x"FF",
		178486 => x"FF",
		178487 => x"FF",
		178488 => x"FF",
		178489 => x"FF",
		178490 => x"FF",
		178491 => x"FF",
		178492 => x"FF",
		178493 => x"FF",
		178494 => x"FF",
		178495 => x"FF",
		178496 => x"FF",
		178497 => x"FF",
		178498 => x"FF",
		178499 => x"FF",
		178500 => x"FF",
		178501 => x"FF",
		178502 => x"FF",
		178503 => x"FF",
		178504 => x"FF",
		178505 => x"FF",
		178506 => x"FF",
		178507 => x"FF",
		178508 => x"FF",
		178509 => x"FF",
		178510 => x"FF",
		178511 => x"FF",
		178512 => x"FF",
		178513 => x"FF",
		178514 => x"FF",
		178515 => x"FF",
		178516 => x"FF",
		178517 => x"FF",
		178518 => x"FF",
		178519 => x"FF",
		178520 => x"FF",
		178521 => x"FF",
		178522 => x"FF",
		178523 => x"FF",
		178524 => x"FF",
		178525 => x"FF",
		178526 => x"FF",
		178527 => x"FF",
		178528 => x"FF",
		178529 => x"FF",
		178530 => x"FF",
		178531 => x"FF",
		178532 => x"FF",
		178533 => x"FF",
		178534 => x"FF",
		178535 => x"FF",
		178536 => x"FF",
		178537 => x"FF",
		178538 => x"FF",
		178539 => x"FF",
		178540 => x"FF",
		178541 => x"FF",
		178542 => x"FF",
		178543 => x"FF",
		178544 => x"FF",
		178545 => x"FF",
		178546 => x"FF",
		178547 => x"FF",
		178548 => x"FF",
		178549 => x"FF",
		178550 => x"FF",
		178551 => x"FF",
		178552 => x"FF",
		178553 => x"FF",
		178554 => x"FF",
		178555 => x"FF",
		178556 => x"FF",
		178557 => x"FF",
		178558 => x"FF",
		178559 => x"FF",
		178560 => x"FF",
		178561 => x"FF",
		178562 => x"FF",
		178563 => x"FF",
		178564 => x"FF",
		178565 => x"FF",
		178566 => x"FF",
		178567 => x"FF",
		178568 => x"FF",
		178569 => x"FF",
		178570 => x"FF",
		178571 => x"FF",
		178572 => x"FF",
		178573 => x"FF",
		178574 => x"FF",
		178575 => x"FF",
		178576 => x"FF",
		178577 => x"FF",
		178578 => x"FF",
		178579 => x"FF",
		178580 => x"FF",
		178581 => x"FF",
		178582 => x"FF",
		178583 => x"FF",
		178584 => x"FF",
		178585 => x"FF",
		178586 => x"FF",
		178587 => x"FF",
		178588 => x"FF",
		178589 => x"FF",
		178590 => x"FF",
		178591 => x"FF",
		178592 => x"FF",
		178593 => x"FF",
		178594 => x"FF",
		178595 => x"FF",
		178596 => x"FF",
		178597 => x"FF",
		178598 => x"FF",
		178599 => x"FF",
		178600 => x"FF",
		178601 => x"FF",
		178602 => x"FF",
		178603 => x"FF",
		178604 => x"FF",
		178605 => x"FF",
		178606 => x"FF",
		178607 => x"FF",
		178608 => x"FF",
		178609 => x"FF",
		178610 => x"FF",
		178611 => x"FF",
		178612 => x"FF",
		178613 => x"FF",
		178614 => x"FF",
		178615 => x"FF",
		178616 => x"FF",
		178617 => x"FF",
		178618 => x"FF",
		178619 => x"FF",
		178620 => x"FF",
		178621 => x"FF",
		178622 => x"FF",
		178623 => x"FF",
		178624 => x"FF",
		178625 => x"FF",
		178626 => x"FF",
		178627 => x"FF",
		178628 => x"FF",
		178629 => x"FF",
		178630 => x"FF",
		178631 => x"FF",
		178632 => x"FF",
		178633 => x"FF",
		178634 => x"FF",
		178635 => x"FF",
		178636 => x"FF",
		178637 => x"FF",
		178638 => x"FF",
		178639 => x"FF",
		178640 => x"FF",
		178641 => x"FF",
		178642 => x"FF",
		178643 => x"FF",
		178644 => x"FF",
		178645 => x"FF",
		178646 => x"FF",
		178647 => x"FF",
		178648 => x"FF",
		178649 => x"FF",
		178650 => x"FF",
		178651 => x"FF",
		178652 => x"FF",
		178653 => x"FF",
		178654 => x"FF",
		178655 => x"FF",
		178656 => x"FF",
		178657 => x"FF",
		178658 => x"FF",
		178659 => x"FF",
		178660 => x"FF",
		178661 => x"FF",
		178662 => x"FF",
		178663 => x"FF",
		178664 => x"FF",
		178665 => x"FF",
		178666 => x"FF",
		178667 => x"FF",
		178668 => x"FF",
		178669 => x"FF",
		178670 => x"FF",
		178671 => x"FF",
		178672 => x"FF",
		178673 => x"FF",
		179318 => x"FF",
		179319 => x"FF",
		179320 => x"FF",
		179321 => x"FF",
		179322 => x"FF",
		179323 => x"FF",
		179324 => x"FF",
		179325 => x"FF",
		179326 => x"FF",
		179327 => x"FF",
		179328 => x"FF",
		179329 => x"FF",
		179330 => x"FF",
		179331 => x"FF",
		179332 => x"FF",
		179333 => x"FF",
		179334 => x"FF",
		179335 => x"FF",
		179336 => x"FF",
		179337 => x"FF",
		179338 => x"FF",
		179339 => x"FF",
		179340 => x"FF",
		179341 => x"FF",
		179342 => x"FF",
		179343 => x"FF",
		179344 => x"FF",
		179345 => x"FF",
		179346 => x"FF",
		179347 => x"FF",
		179348 => x"FF",
		179349 => x"FF",
		179350 => x"FF",
		179351 => x"FF",
		179352 => x"FF",
		179353 => x"FF",
		179354 => x"FF",
		179355 => x"FF",
		179356 => x"FF",
		179357 => x"FF",
		179358 => x"FF",
		179359 => x"FF",
		179360 => x"FF",
		179361 => x"FF",
		179362 => x"FF",
		179363 => x"FF",
		179364 => x"FF",
		179365 => x"FF",
		179366 => x"FF",
		179367 => x"FF",
		179368 => x"FF",
		179369 => x"FF",
		179370 => x"FF",
		179371 => x"FF",
		179372 => x"FF",
		179373 => x"FF",
		179374 => x"FF",
		179375 => x"FF",
		179376 => x"FF",
		179377 => x"FF",
		179378 => x"FF",
		179379 => x"FF",
		179380 => x"FF",
		179381 => x"FF",
		179382 => x"FF",
		179383 => x"FF",
		179384 => x"FF",
		179385 => x"FF",
		179386 => x"FF",
		179387 => x"FF",
		179388 => x"FF",
		179389 => x"FF",
		179390 => x"FF",
		179391 => x"FF",
		179392 => x"FF",
		179393 => x"FF",
		179394 => x"FF",
		179395 => x"FF",
		179396 => x"FF",
		179397 => x"FF",
		179398 => x"FF",
		179399 => x"FF",
		179400 => x"FF",
		179401 => x"FF",
		179402 => x"FF",
		179403 => x"FF",
		179404 => x"FF",
		179405 => x"FF",
		179406 => x"FF",
		179407 => x"FF",
		179408 => x"FF",
		179409 => x"FF",
		179410 => x"FF",
		179411 => x"FF",
		179412 => x"FF",
		179413 => x"FF",
		179414 => x"FF",
		179415 => x"FF",
		179416 => x"FF",
		179417 => x"FF",
		179418 => x"FF",
		179419 => x"FF",
		179420 => x"FF",
		179421 => x"FF",
		179422 => x"FF",
		179423 => x"FF",
		179424 => x"FF",
		179425 => x"FF",
		179426 => x"FF",
		179427 => x"FF",
		179428 => x"FF",
		179429 => x"FF",
		179430 => x"FF",
		179431 => x"FF",
		179432 => x"FF",
		179433 => x"FF",
		179434 => x"FF",
		179435 => x"FF",
		179436 => x"FF",
		179437 => x"FF",
		179438 => x"FF",
		179439 => x"FF",
		179440 => x"FF",
		179441 => x"FF",
		179442 => x"FF",
		179443 => x"FF",
		179444 => x"FF",
		179445 => x"FF",
		179446 => x"FF",
		179447 => x"FF",
		179448 => x"FF",
		179449 => x"FF",
		179450 => x"FF",
		179451 => x"FF",
		179452 => x"FF",
		179453 => x"FF",
		179454 => x"FF",
		179455 => x"FF",
		179456 => x"FF",
		179457 => x"FF",
		179458 => x"FF",
		179459 => x"FF",
		179460 => x"FF",
		179461 => x"FF",
		179462 => x"FF",
		179463 => x"FF",
		179464 => x"FF",
		179465 => x"FF",
		179466 => x"FF",
		179467 => x"FF",
		179468 => x"FF",
		179469 => x"FF",
		179470 => x"FF",
		179471 => x"FF",
		179472 => x"FF",
		179473 => x"FF",
		179474 => x"FF",
		179475 => x"FF",
		179476 => x"FF",
		179477 => x"FF",
		179478 => x"FF",
		179479 => x"FF",
		179480 => x"FF",
		179481 => x"FF",
		179482 => x"FF",
		179483 => x"FF",
		179484 => x"FF",
		179485 => x"FF",
		179486 => x"FF",
		179487 => x"FF",
		179488 => x"FF",
		179489 => x"FF",
		179490 => x"FF",
		179491 => x"FF",
		179492 => x"FF",
		179493 => x"FF",
		179494 => x"FF",
		179495 => x"FF",
		179496 => x"FF",
		179497 => x"FF",
		179498 => x"FF",
		179499 => x"FF",
		179500 => x"FF",
		179501 => x"FF",
		179502 => x"FF",
		179503 => x"FF",
		179504 => x"FF",
		179505 => x"FF",
		179506 => x"FF",
		179507 => x"FF",
		179508 => x"FF",
		179509 => x"FF",
		179510 => x"FF",
		179511 => x"FF",
		179512 => x"FF",
		179513 => x"FF",
		179514 => x"FF",
		179515 => x"FF",
		179516 => x"FF",
		179517 => x"FF",
		179518 => x"FF",
		179519 => x"FF",
		179520 => x"FF",
		179521 => x"FF",
		179522 => x"FF",
		179523 => x"FF",
		179524 => x"FF",
		179525 => x"FF",
		179526 => x"FF",
		179527 => x"FF",
		179528 => x"FF",
		179529 => x"FF",
		179530 => x"FF",
		179531 => x"FF",
		179532 => x"FF",
		179533 => x"FF",
		179534 => x"FF",
		179535 => x"FF",
		179536 => x"FF",
		179537 => x"FF",
		179538 => x"FF",
		179539 => x"FF",
		179540 => x"FF",
		179541 => x"FF",
		179542 => x"FF",
		179543 => x"FF",
		179544 => x"FF",
		179545 => x"FF",
		179546 => x"FF",
		179547 => x"FF",
		179548 => x"FF",
		179549 => x"FF",
		179550 => x"FF",
		179551 => x"FF",
		179552 => x"FF",
		179553 => x"FF",
		179554 => x"FF",
		179555 => x"FF",
		179556 => x"FF",
		179557 => x"FF",
		179558 => x"FF",
		179559 => x"FF",
		179560 => x"FF",
		179561 => x"FF",
		179562 => x"FF",
		179563 => x"FF",
		179564 => x"FF",
		179565 => x"FF",
		179566 => x"FF",
		179567 => x"FF",
		179568 => x"FF",
		179569 => x"FF",
		179570 => x"FF",
		179571 => x"FF",
		179572 => x"FF",
		179573 => x"FF",
		179574 => x"FF",
		179575 => x"FF",
		179576 => x"FF",
		179577 => x"FF",
		179578 => x"FF",
		179579 => x"FF",
		179580 => x"FF",
		179581 => x"FF",
		179582 => x"FF",
		179583 => x"FF",
		179584 => x"FF",
		179585 => x"FF",
		179586 => x"FF",
		179587 => x"FF",
		179588 => x"FF",
		179589 => x"FF",
		179590 => x"FF",
		179591 => x"FF",
		179592 => x"FF",
		179593 => x"FF",
		179594 => x"FF",
		179595 => x"FF",
		179596 => x"FF",
		179597 => x"FF",
		179598 => x"FF",
		179599 => x"FF",
		179600 => x"FF",
		179601 => x"FF",
		179602 => x"FF",
		179603 => x"FF",
		179604 => x"FF",
		179605 => x"FF",
		179606 => x"FF",
		179607 => x"FF",
		179608 => x"FF",
		179609 => x"FF",
		179610 => x"FF",
		179611 => x"FF",
		179612 => x"FF",
		179613 => x"FF",
		179614 => x"FF",
		179615 => x"FF",
		179616 => x"FF",
		179617 => x"FF",
		179618 => x"FF",
		179619 => x"FF",
		179620 => x"FF",
		179621 => x"FF",
		179622 => x"FF",
		179623 => x"FF",
		179624 => x"FF",
		179625 => x"FF",
		179626 => x"FF",
		179627 => x"FF",
		179628 => x"FF",
		179629 => x"FF",
		179630 => x"FF",
		179631 => x"FF",
		179632 => x"FF",
		179633 => x"FF",
		179634 => x"FF",
		179635 => x"FF",
		179636 => x"FF",
		179637 => x"FF",
		179638 => x"FF",
		179639 => x"FF",
		179640 => x"FF",
		179641 => x"FF",
		179642 => x"FF",
		179643 => x"FF",
		179644 => x"FF",
		179645 => x"FF",
		179646 => x"FF",
		179647 => x"FF",
		179648 => x"FF",
		179649 => x"FF",
		179650 => x"FF",
		179651 => x"FF",
		179652 => x"FF",
		179653 => x"FF",
		179654 => x"FF",
		179655 => x"FF",
		179656 => x"FF",
		179657 => x"FF",
		179658 => x"FF",
		179659 => x"FF",
		179660 => x"FF",
		179661 => x"FF",
		179662 => x"FF",
		179663 => x"FF",
		179664 => x"FF",
		179665 => x"FF",
		179666 => x"FF",
		179667 => x"FF",
		179668 => x"FF",
		179669 => x"FF",
		179670 => x"FF",
		179671 => x"FF",
		179672 => x"FF",
		179673 => x"FF",
		179674 => x"FF",
		179675 => x"FF",
		179676 => x"FF",
		179677 => x"FF",
		179678 => x"FF",
		179679 => x"FF",
		179680 => x"FF",
		179681 => x"FF",
		179682 => x"FF",
		179683 => x"FF",
		179684 => x"FF",
		179685 => x"FF",
		179686 => x"FF",
		179687 => x"FF",
		179688 => x"FF",
		179689 => x"FF",
		179690 => x"FF",
		179691 => x"FF",
		179692 => x"FF",
		179693 => x"FF",
		179694 => x"FF",
		179695 => x"FF",
		179696 => x"FF",
		179697 => x"FF",
		180342 => x"FF",
		180343 => x"FF",
		180344 => x"FF",
		180345 => x"FF",
		180346 => x"FF",
		180347 => x"FF",
		180348 => x"FF",
		180349 => x"FF",
		180350 => x"FF",
		180351 => x"FF",
		180352 => x"FF",
		180353 => x"FF",
		180354 => x"FF",
		180355 => x"FF",
		180356 => x"FF",
		180357 => x"FF",
		180358 => x"FF",
		180359 => x"FF",
		180360 => x"FF",
		180361 => x"FF",
		180362 => x"FF",
		180363 => x"FF",
		180364 => x"FF",
		180365 => x"FF",
		180366 => x"FF",
		180367 => x"FF",
		180368 => x"FF",
		180369 => x"FF",
		180370 => x"FF",
		180371 => x"FF",
		180372 => x"FF",
		180373 => x"FF",
		180374 => x"FF",
		180375 => x"FF",
		180376 => x"FF",
		180377 => x"FF",
		180378 => x"FF",
		180379 => x"FF",
		180380 => x"FF",
		180381 => x"FF",
		180382 => x"FF",
		180383 => x"FF",
		180384 => x"FF",
		180385 => x"FF",
		180386 => x"FF",
		180387 => x"FF",
		180388 => x"FF",
		180389 => x"FF",
		180390 => x"FF",
		180391 => x"FF",
		180392 => x"FF",
		180393 => x"FF",
		180394 => x"FF",
		180395 => x"FF",
		180396 => x"FF",
		180397 => x"FF",
		180398 => x"FF",
		180399 => x"FF",
		180400 => x"FF",
		180401 => x"FF",
		180402 => x"FF",
		180403 => x"FF",
		180404 => x"FF",
		180405 => x"FF",
		180406 => x"FF",
		180407 => x"FF",
		180408 => x"FF",
		180409 => x"FF",
		180410 => x"FF",
		180411 => x"FF",
		180412 => x"FF",
		180413 => x"FF",
		180414 => x"FF",
		180415 => x"FF",
		180416 => x"FF",
		180417 => x"FF",
		180418 => x"FF",
		180419 => x"FF",
		180420 => x"FF",
		180421 => x"FF",
		180422 => x"FF",
		180423 => x"FF",
		180424 => x"FF",
		180425 => x"FF",
		180426 => x"FF",
		180427 => x"FF",
		180428 => x"FF",
		180429 => x"FF",
		180430 => x"FF",
		180431 => x"FF",
		180432 => x"FF",
		180433 => x"FF",
		180434 => x"FF",
		180435 => x"FF",
		180436 => x"FF",
		180437 => x"FF",
		180438 => x"FF",
		180439 => x"FF",
		180440 => x"FF",
		180441 => x"FF",
		180442 => x"FF",
		180443 => x"FF",
		180444 => x"FF",
		180445 => x"FF",
		180446 => x"FF",
		180447 => x"FF",
		180448 => x"FF",
		180449 => x"FF",
		180450 => x"FF",
		180451 => x"FF",
		180452 => x"FF",
		180453 => x"FF",
		180454 => x"FF",
		180455 => x"FF",
		180456 => x"FF",
		180457 => x"FF",
		180458 => x"FF",
		180459 => x"FF",
		180460 => x"FF",
		180461 => x"FF",
		180462 => x"FF",
		180463 => x"FF",
		180464 => x"FF",
		180465 => x"FF",
		180466 => x"FF",
		180467 => x"FF",
		180468 => x"FF",
		180469 => x"FF",
		180470 => x"FF",
		180471 => x"FF",
		180472 => x"FF",
		180473 => x"FF",
		180474 => x"FF",
		180475 => x"FF",
		180476 => x"FF",
		180477 => x"FF",
		180478 => x"FF",
		180479 => x"FF",
		180480 => x"FF",
		180481 => x"FF",
		180482 => x"FF",
		180483 => x"FF",
		180484 => x"FF",
		180485 => x"FF",
		180486 => x"FF",
		180487 => x"FF",
		180488 => x"FF",
		180489 => x"FF",
		180490 => x"FF",
		180491 => x"FF",
		180492 => x"FF",
		180493 => x"FF",
		180494 => x"FF",
		180495 => x"FF",
		180496 => x"FF",
		180497 => x"FF",
		180498 => x"FF",
		180499 => x"FF",
		180500 => x"FF",
		180501 => x"FF",
		180502 => x"FF",
		180503 => x"FF",
		180504 => x"FF",
		180505 => x"FF",
		180506 => x"FF",
		180507 => x"FF",
		180508 => x"FF",
		180509 => x"FF",
		180510 => x"FF",
		180511 => x"FF",
		180512 => x"FF",
		180513 => x"FF",
		180514 => x"FF",
		180515 => x"FF",
		180516 => x"FF",
		180517 => x"FF",
		180518 => x"FF",
		180519 => x"FF",
		180520 => x"FF",
		180521 => x"FF",
		180522 => x"FF",
		180523 => x"FF",
		180524 => x"FF",
		180525 => x"FF",
		180526 => x"FF",
		180527 => x"FF",
		180528 => x"FF",
		180529 => x"FF",
		180530 => x"FF",
		180531 => x"FF",
		180532 => x"FF",
		180533 => x"FF",
		180534 => x"FF",
		180535 => x"FF",
		180536 => x"FF",
		180537 => x"FF",
		180538 => x"FF",
		180539 => x"FF",
		180540 => x"FF",
		180541 => x"FF",
		180542 => x"FF",
		180543 => x"FF",
		180544 => x"FF",
		180545 => x"FF",
		180546 => x"FF",
		180547 => x"FF",
		180548 => x"FF",
		180549 => x"FF",
		180550 => x"FF",
		180551 => x"FF",
		180552 => x"FF",
		180553 => x"FF",
		180554 => x"FF",
		180555 => x"FF",
		180556 => x"FF",
		180557 => x"FF",
		180558 => x"FF",
		180559 => x"FF",
		180560 => x"FF",
		180561 => x"FF",
		180562 => x"FF",
		180563 => x"FF",
		180564 => x"FF",
		180565 => x"FF",
		180566 => x"FF",
		180567 => x"FF",
		180568 => x"FF",
		180569 => x"FF",
		180570 => x"FF",
		180571 => x"FF",
		180572 => x"FF",
		180573 => x"FF",
		180574 => x"FF",
		180575 => x"FF",
		180576 => x"FF",
		180577 => x"FF",
		180578 => x"FF",
		180579 => x"FF",
		180580 => x"FF",
		180581 => x"FF",
		180582 => x"FF",
		180583 => x"FF",
		180584 => x"FF",
		180585 => x"FF",
		180586 => x"FF",
		180587 => x"FF",
		180588 => x"FF",
		180589 => x"FF",
		180590 => x"FF",
		180591 => x"FF",
		180592 => x"FF",
		180593 => x"FF",
		180594 => x"FF",
		180595 => x"FF",
		180596 => x"FF",
		180597 => x"FF",
		180598 => x"FF",
		180599 => x"FF",
		180600 => x"FF",
		180601 => x"FF",
		180602 => x"FF",
		180603 => x"FF",
		180604 => x"FF",
		180605 => x"FF",
		180606 => x"FF",
		180607 => x"FF",
		180608 => x"FF",
		180609 => x"FF",
		180610 => x"FF",
		180611 => x"FF",
		180612 => x"FF",
		180613 => x"FF",
		180614 => x"FF",
		180615 => x"FF",
		180616 => x"FF",
		180617 => x"FF",
		180618 => x"FF",
		180619 => x"FF",
		180620 => x"FF",
		180621 => x"FF",
		180622 => x"FF",
		180623 => x"FF",
		180624 => x"FF",
		180625 => x"FF",
		180626 => x"FF",
		180627 => x"FF",
		180628 => x"FF",
		180629 => x"FF",
		180630 => x"FF",
		180631 => x"FF",
		180632 => x"FF",
		180633 => x"FF",
		180634 => x"FF",
		180635 => x"FF",
		180636 => x"FF",
		180637 => x"FF",
		180638 => x"FF",
		180639 => x"FF",
		180640 => x"FF",
		180641 => x"FF",
		180642 => x"FF",
		180643 => x"FF",
		180644 => x"FF",
		180645 => x"FF",
		180646 => x"FF",
		180647 => x"FF",
		180648 => x"FF",
		180649 => x"FF",
		180650 => x"FF",
		180651 => x"FF",
		180652 => x"FF",
		180653 => x"FF",
		180654 => x"FF",
		180655 => x"FF",
		180656 => x"FF",
		180657 => x"FF",
		180658 => x"FF",
		180659 => x"FF",
		180660 => x"FF",
		180661 => x"FF",
		180662 => x"FF",
		180663 => x"FF",
		180664 => x"FF",
		180665 => x"FF",
		180666 => x"FF",
		180667 => x"FF",
		180668 => x"FF",
		180669 => x"FF",
		180670 => x"FF",
		180671 => x"FF",
		180672 => x"FF",
		180673 => x"FF",
		180674 => x"FF",
		180675 => x"FF",
		180676 => x"FF",
		180677 => x"FF",
		180678 => x"FF",
		180679 => x"FF",
		180680 => x"FF",
		180681 => x"FF",
		180682 => x"FF",
		180683 => x"FF",
		180684 => x"FF",
		180685 => x"FF",
		180686 => x"FF",
		180687 => x"FF",
		180688 => x"FF",
		180689 => x"FF",
		180690 => x"FF",
		180691 => x"FF",
		180692 => x"FF",
		180693 => x"FF",
		180694 => x"FF",
		180695 => x"FF",
		180696 => x"FF",
		180697 => x"FF",
		180698 => x"FF",
		180699 => x"FF",
		180700 => x"FF",
		180701 => x"FF",
		180702 => x"FF",
		180703 => x"FF",
		180704 => x"FF",
		180705 => x"FF",
		180706 => x"FF",
		180707 => x"FF",
		180708 => x"FF",
		180709 => x"FF",
		180710 => x"FF",
		180711 => x"FF",
		180712 => x"FF",
		180713 => x"FF",
		180714 => x"FF",
		180715 => x"FF",
		180716 => x"FF",
		180717 => x"FF",
		180718 => x"FF",
		180719 => x"FF",
		180720 => x"FF",
		180721 => x"FF",
		181366 => x"FF",
		181367 => x"FF",
		181368 => x"FF",
		181369 => x"FF",
		181370 => x"FF",
		181371 => x"FF",
		181372 => x"FF",
		181373 => x"FF",
		181374 => x"FF",
		181375 => x"FF",
		181376 => x"FF",
		181377 => x"FF",
		181378 => x"FF",
		181379 => x"FF",
		181380 => x"FF",
		181381 => x"FF",
		181382 => x"FF",
		181383 => x"FF",
		181384 => x"FF",
		181385 => x"FF",
		181386 => x"FF",
		181387 => x"FF",
		181388 => x"FF",
		181389 => x"FF",
		181390 => x"FF",
		181391 => x"FF",
		181392 => x"FF",
		181393 => x"FF",
		181394 => x"FF",
		181395 => x"FF",
		181396 => x"FF",
		181397 => x"FF",
		181398 => x"FF",
		181399 => x"FF",
		181400 => x"FF",
		181401 => x"FF",
		181402 => x"FF",
		181403 => x"FF",
		181404 => x"FF",
		181405 => x"FF",
		181406 => x"FF",
		181407 => x"FF",
		181408 => x"FF",
		181409 => x"FF",
		181410 => x"FF",
		181411 => x"FF",
		181412 => x"FF",
		181413 => x"FF",
		181414 => x"FF",
		181415 => x"FF",
		181416 => x"FF",
		181417 => x"FF",
		181418 => x"FF",
		181419 => x"FF",
		181420 => x"FF",
		181421 => x"FF",
		181422 => x"FF",
		181423 => x"FF",
		181424 => x"FF",
		181425 => x"FF",
		181426 => x"FF",
		181427 => x"FF",
		181428 => x"FF",
		181429 => x"FF",
		181430 => x"FF",
		181431 => x"FF",
		181432 => x"FF",
		181433 => x"FF",
		181434 => x"FF",
		181435 => x"FF",
		181436 => x"FF",
		181437 => x"FF",
		181438 => x"FF",
		181439 => x"FF",
		181440 => x"FF",
		181441 => x"FF",
		181442 => x"FF",
		181443 => x"FF",
		181444 => x"FF",
		181445 => x"FF",
		181446 => x"FF",
		181447 => x"FF",
		181448 => x"FF",
		181449 => x"FF",
		181450 => x"FF",
		181451 => x"FF",
		181452 => x"FF",
		181453 => x"FF",
		181454 => x"FF",
		181455 => x"FF",
		181456 => x"FF",
		181457 => x"FF",
		181458 => x"FF",
		181459 => x"FF",
		181460 => x"FF",
		181461 => x"FF",
		181462 => x"FF",
		181463 => x"FF",
		181464 => x"FF",
		181465 => x"FF",
		181466 => x"FF",
		181467 => x"FF",
		181468 => x"FF",
		181469 => x"FF",
		181470 => x"FF",
		181471 => x"FF",
		181472 => x"FF",
		181473 => x"FF",
		181474 => x"FF",
		181475 => x"FF",
		181476 => x"FF",
		181477 => x"FF",
		181478 => x"FF",
		181479 => x"FF",
		181480 => x"FF",
		181481 => x"FF",
		181482 => x"FF",
		181483 => x"FF",
		181484 => x"FF",
		181485 => x"FF",
		181486 => x"FF",
		181487 => x"FF",
		181488 => x"FF",
		181489 => x"FF",
		181490 => x"FF",
		181491 => x"FF",
		181492 => x"FF",
		181493 => x"FF",
		181494 => x"FF",
		181495 => x"FF",
		181496 => x"FF",
		181497 => x"FF",
		181498 => x"FF",
		181499 => x"FF",
		181500 => x"FF",
		181501 => x"FF",
		181502 => x"FF",
		181503 => x"FF",
		181504 => x"FF",
		181505 => x"FF",
		181506 => x"FF",
		181507 => x"FF",
		181508 => x"FF",
		181509 => x"FF",
		181510 => x"FF",
		181511 => x"FF",
		181512 => x"FF",
		181513 => x"FF",
		181514 => x"FF",
		181515 => x"FF",
		181516 => x"FF",
		181517 => x"FF",
		181518 => x"FF",
		181519 => x"FF",
		181520 => x"FF",
		181521 => x"FF",
		181522 => x"FF",
		181523 => x"FF",
		181524 => x"FF",
		181525 => x"FF",
		181526 => x"FF",
		181527 => x"FF",
		181528 => x"FF",
		181529 => x"FF",
		181530 => x"FF",
		181531 => x"FF",
		181532 => x"FF",
		181533 => x"FF",
		181534 => x"FF",
		181535 => x"FF",
		181536 => x"FF",
		181537 => x"FF",
		181538 => x"FF",
		181539 => x"FF",
		181540 => x"FF",
		181541 => x"FF",
		181542 => x"FF",
		181543 => x"FF",
		181544 => x"FF",
		181545 => x"FF",
		181546 => x"FF",
		181547 => x"FF",
		181548 => x"FF",
		181549 => x"FF",
		181550 => x"FF",
		181551 => x"FF",
		181552 => x"FF",
		181553 => x"FF",
		181554 => x"FF",
		181555 => x"FF",
		181556 => x"FF",
		181557 => x"FF",
		181558 => x"FF",
		181559 => x"FF",
		181560 => x"FF",
		181561 => x"FF",
		181562 => x"FF",
		181563 => x"FF",
		181564 => x"FF",
		181565 => x"FF",
		181566 => x"FF",
		181567 => x"FF",
		181568 => x"FF",
		181569 => x"FF",
		181570 => x"FF",
		181571 => x"FF",
		181572 => x"FF",
		181573 => x"FF",
		181574 => x"FF",
		181575 => x"FF",
		181576 => x"FF",
		181577 => x"FF",
		181578 => x"FF",
		181579 => x"FF",
		181580 => x"FF",
		181581 => x"FF",
		181582 => x"FF",
		181583 => x"FF",
		181584 => x"FF",
		181585 => x"FF",
		181586 => x"FF",
		181587 => x"FF",
		181588 => x"FF",
		181589 => x"FF",
		181590 => x"FF",
		181591 => x"FF",
		181592 => x"FF",
		181593 => x"FF",
		181594 => x"FF",
		181595 => x"FF",
		181596 => x"FF",
		181597 => x"FF",
		181598 => x"FF",
		181599 => x"FF",
		181600 => x"FF",
		181601 => x"FF",
		181602 => x"FF",
		181603 => x"FF",
		181604 => x"FF",
		181605 => x"FF",
		181606 => x"FF",
		181607 => x"FF",
		181608 => x"FF",
		181609 => x"FF",
		181610 => x"FF",
		181611 => x"FF",
		181612 => x"FF",
		181613 => x"FF",
		181614 => x"FF",
		181615 => x"FF",
		181616 => x"FF",
		181617 => x"FF",
		181618 => x"FF",
		181619 => x"FF",
		181620 => x"FF",
		181621 => x"FF",
		181622 => x"FF",
		181623 => x"FF",
		181624 => x"FF",
		181625 => x"FF",
		181626 => x"FF",
		181627 => x"FF",
		181628 => x"FF",
		181629 => x"FF",
		181630 => x"FF",
		181631 => x"FF",
		181632 => x"FF",
		181633 => x"FF",
		181634 => x"FF",
		181635 => x"FF",
		181636 => x"FF",
		181637 => x"FF",
		181638 => x"FF",
		181639 => x"FF",
		181640 => x"FF",
		181641 => x"FF",
		181642 => x"FF",
		181643 => x"FF",
		181644 => x"FF",
		181645 => x"FF",
		181646 => x"FF",
		181647 => x"FF",
		181648 => x"FF",
		181649 => x"FF",
		181650 => x"FF",
		181651 => x"FF",
		181652 => x"FF",
		181653 => x"FF",
		181654 => x"FF",
		181655 => x"FF",
		181656 => x"FF",
		181657 => x"FF",
		181658 => x"FF",
		181659 => x"FF",
		181660 => x"FF",
		181661 => x"FF",
		181662 => x"FF",
		181663 => x"FF",
		181664 => x"FF",
		181665 => x"FF",
		181666 => x"FF",
		181667 => x"FF",
		181668 => x"FF",
		181669 => x"FF",
		181670 => x"FF",
		181671 => x"FF",
		181672 => x"FF",
		181673 => x"FF",
		181674 => x"FF",
		181675 => x"FF",
		181676 => x"FF",
		181677 => x"FF",
		181678 => x"FF",
		181679 => x"FF",
		181680 => x"FF",
		181681 => x"FF",
		181682 => x"FF",
		181683 => x"FF",
		181684 => x"FF",
		181685 => x"FF",
		181686 => x"FF",
		181687 => x"FF",
		181688 => x"FF",
		181689 => x"FF",
		181690 => x"FF",
		181691 => x"FF",
		181692 => x"FF",
		181693 => x"FF",
		181694 => x"FF",
		181695 => x"FF",
		181696 => x"FF",
		181697 => x"FF",
		181698 => x"FF",
		181699 => x"FF",
		181700 => x"FF",
		181701 => x"FF",
		181702 => x"FF",
		181703 => x"FF",
		181704 => x"FF",
		181705 => x"FF",
		181706 => x"FF",
		181707 => x"FF",
		181708 => x"FF",
		181709 => x"FF",
		181710 => x"FF",
		181711 => x"FF",
		181712 => x"FF",
		181713 => x"FF",
		181714 => x"FF",
		181715 => x"FF",
		181716 => x"FF",
		181717 => x"FF",
		181718 => x"FF",
		181719 => x"FF",
		181720 => x"FF",
		181721 => x"FF",
		181722 => x"FF",
		181723 => x"FF",
		181724 => x"FF",
		181725 => x"FF",
		181726 => x"FF",
		181727 => x"FF",
		181728 => x"FF",
		181729 => x"FF",
		181730 => x"FF",
		181731 => x"FF",
		181732 => x"FF",
		181733 => x"FF",
		181734 => x"FF",
		181735 => x"FF",
		181736 => x"FF",
		181737 => x"FF",
		181738 => x"FF",
		181739 => x"FF",
		181740 => x"FF",
		181741 => x"FF",
		181742 => x"FF",
		181743 => x"FF",
		181744 => x"FF",
		181745 => x"FF",
		182390 => x"FF",
		182391 => x"FF",
		182392 => x"FF",
		182393 => x"FF",
		182394 => x"FF",
		182515 => x"FF",
		182516 => x"FF",
		182517 => x"FF",
		182518 => x"FF",
		182519 => x"FF",
		182640 => x"FF",
		182641 => x"FF",
		182642 => x"FF",
		182643 => x"FF",
		182644 => x"FF",
		182765 => x"FF",
		182766 => x"FF",
		182767 => x"FF",
		182768 => x"FF",
		182769 => x"FF",
		183414 => x"FF",
		183415 => x"FF",
		183416 => x"FF",
		183417 => x"FF",
		183418 => x"FF",
		183539 => x"FF",
		183540 => x"FF",
		183541 => x"FF",
		183542 => x"FF",
		183543 => x"FF",
		183664 => x"FF",
		183665 => x"FF",
		183666 => x"FF",
		183667 => x"FF",
		183668 => x"FF",
		183789 => x"FF",
		183790 => x"FF",
		183791 => x"FF",
		183792 => x"FF",
		183793 => x"FF",
		184438 => x"FF",
		184439 => x"FF",
		184440 => x"FF",
		184441 => x"FF",
		184442 => x"FF",
		184563 => x"FF",
		184564 => x"FF",
		184565 => x"FF",
		184566 => x"FF",
		184567 => x"FF",
		184688 => x"FF",
		184689 => x"FF",
		184690 => x"FF",
		184691 => x"FF",
		184692 => x"FF",
		184813 => x"FF",
		184814 => x"FF",
		184815 => x"FF",
		184816 => x"FF",
		184817 => x"FF",
		185462 => x"FF",
		185463 => x"FF",
		185464 => x"FF",
		185465 => x"FF",
		185466 => x"FF",
		185587 => x"FF",
		185588 => x"FF",
		185589 => x"FF",
		185590 => x"FF",
		185591 => x"FF",
		185712 => x"FF",
		185713 => x"FF",
		185714 => x"FF",
		185715 => x"FF",
		185716 => x"FF",
		185837 => x"FF",
		185838 => x"FF",
		185839 => x"FF",
		185840 => x"FF",
		185841 => x"FF",
		186486 => x"FF",
		186487 => x"FF",
		186488 => x"FF",
		186489 => x"FF",
		186490 => x"FF",
		186611 => x"FF",
		186612 => x"FF",
		186613 => x"FF",
		186614 => x"FF",
		186615 => x"FF",
		186736 => x"FF",
		186737 => x"FF",
		186738 => x"FF",
		186739 => x"FF",
		186740 => x"FF",
		186861 => x"FF",
		186862 => x"FF",
		186863 => x"FF",
		186864 => x"FF",
		186865 => x"FF",
		187510 => x"FF",
		187511 => x"FF",
		187512 => x"FF",
		187513 => x"FF",
		187514 => x"FF",
		187635 => x"FF",
		187636 => x"FF",
		187637 => x"FF",
		187638 => x"FF",
		187639 => x"FF",
		187760 => x"FF",
		187761 => x"FF",
		187762 => x"FF",
		187763 => x"FF",
		187764 => x"FF",
		187885 => x"FF",
		187886 => x"FF",
		187887 => x"FF",
		187888 => x"FF",
		187889 => x"FF",
		188534 => x"FF",
		188535 => x"FF",
		188536 => x"FF",
		188537 => x"FF",
		188538 => x"FF",
		188659 => x"FF",
		188660 => x"FF",
		188661 => x"FF",
		188662 => x"FF",
		188663 => x"FF",
		188784 => x"FF",
		188785 => x"FF",
		188786 => x"FF",
		188787 => x"FF",
		188788 => x"FF",
		188909 => x"FF",
		188910 => x"FF",
		188911 => x"FF",
		188912 => x"FF",
		188913 => x"FF",
		189558 => x"FF",
		189559 => x"FF",
		189560 => x"FF",
		189561 => x"FF",
		189562 => x"FF",
		189683 => x"FF",
		189684 => x"FF",
		189685 => x"FF",
		189686 => x"FF",
		189687 => x"FF",
		189808 => x"FF",
		189809 => x"FF",
		189810 => x"FF",
		189811 => x"FF",
		189812 => x"FF",
		189933 => x"FF",
		189934 => x"FF",
		189935 => x"FF",
		189936 => x"FF",
		189937 => x"FF",
		190582 => x"FF",
		190583 => x"FF",
		190584 => x"FF",
		190585 => x"FF",
		190586 => x"FF",
		190707 => x"FF",
		190708 => x"FF",
		190709 => x"FF",
		190710 => x"FF",
		190711 => x"FF",
		190832 => x"FF",
		190833 => x"FF",
		190834 => x"FF",
		190835 => x"FF",
		190836 => x"FF",
		190957 => x"FF",
		190958 => x"FF",
		190959 => x"FF",
		190960 => x"FF",
		190961 => x"FF",
		191606 => x"FF",
		191607 => x"FF",
		191608 => x"FF",
		191609 => x"FF",
		191610 => x"FF",
		191731 => x"FF",
		191732 => x"FF",
		191733 => x"FF",
		191734 => x"FF",
		191735 => x"FF",
		191856 => x"FF",
		191857 => x"FF",
		191858 => x"FF",
		191859 => x"FF",
		191860 => x"FF",
		191981 => x"FF",
		191982 => x"FF",
		191983 => x"FF",
		191984 => x"FF",
		191985 => x"FF",
		192630 => x"FF",
		192631 => x"FF",
		192632 => x"FF",
		192633 => x"FF",
		192634 => x"FF",
		192755 => x"FF",
		192756 => x"FF",
		192757 => x"FF",
		192758 => x"FF",
		192759 => x"FF",
		192880 => x"FF",
		192881 => x"FF",
		192882 => x"FF",
		192883 => x"FF",
		192884 => x"FF",
		193005 => x"FF",
		193006 => x"FF",
		193007 => x"FF",
		193008 => x"FF",
		193009 => x"FF",
		193654 => x"FF",
		193655 => x"FF",
		193656 => x"FF",
		193657 => x"FF",
		193658 => x"FF",
		193779 => x"FF",
		193780 => x"FF",
		193781 => x"FF",
		193782 => x"FF",
		193783 => x"FF",
		193904 => x"FF",
		193905 => x"FF",
		193906 => x"FF",
		193907 => x"FF",
		193908 => x"FF",
		194029 => x"FF",
		194030 => x"FF",
		194031 => x"FF",
		194032 => x"FF",
		194033 => x"FF",
		194678 => x"FF",
		194679 => x"FF",
		194680 => x"FF",
		194681 => x"FF",
		194682 => x"FF",
		194803 => x"FF",
		194804 => x"FF",
		194805 => x"FF",
		194806 => x"FF",
		194807 => x"FF",
		194928 => x"FF",
		194929 => x"FF",
		194930 => x"FF",
		194931 => x"FF",
		194932 => x"FF",
		195053 => x"FF",
		195054 => x"FF",
		195055 => x"FF",
		195056 => x"FF",
		195057 => x"FF",
		195702 => x"FF",
		195703 => x"FF",
		195704 => x"FF",
		195705 => x"FF",
		195706 => x"FF",
		195827 => x"FF",
		195828 => x"FF",
		195829 => x"FF",
		195830 => x"FF",
		195831 => x"FF",
		195952 => x"FF",
		195953 => x"FF",
		195954 => x"FF",
		195955 => x"FF",
		195956 => x"FF",
		196077 => x"FF",
		196078 => x"FF",
		196079 => x"FF",
		196080 => x"FF",
		196081 => x"FF",
		196726 => x"FF",
		196727 => x"FF",
		196728 => x"FF",
		196729 => x"FF",
		196730 => x"FF",
		196851 => x"FF",
		196852 => x"FF",
		196853 => x"FF",
		196854 => x"FF",
		196855 => x"FF",
		196976 => x"FF",
		196977 => x"FF",
		196978 => x"FF",
		196979 => x"FF",
		196980 => x"FF",
		197101 => x"FF",
		197102 => x"FF",
		197103 => x"FF",
		197104 => x"FF",
		197105 => x"FF",
		197750 => x"FF",
		197751 => x"FF",
		197752 => x"FF",
		197753 => x"FF",
		197754 => x"FF",
		197875 => x"FF",
		197876 => x"FF",
		197877 => x"FF",
		197878 => x"FF",
		197879 => x"FF",
		198000 => x"FF",
		198001 => x"FF",
		198002 => x"FF",
		198003 => x"FF",
		198004 => x"FF",
		198125 => x"FF",
		198126 => x"FF",
		198127 => x"FF",
		198128 => x"FF",
		198129 => x"FF",
		198774 => x"FF",
		198775 => x"FF",
		198776 => x"FF",
		198777 => x"FF",
		198778 => x"FF",
		198899 => x"FF",
		198900 => x"FF",
		198901 => x"FF",
		198902 => x"FF",
		198903 => x"FF",
		199024 => x"FF",
		199025 => x"FF",
		199026 => x"FF",
		199027 => x"FF",
		199028 => x"FF",
		199149 => x"FF",
		199150 => x"FF",
		199151 => x"FF",
		199152 => x"FF",
		199153 => x"FF",
		199798 => x"FF",
		199799 => x"FF",
		199800 => x"FF",
		199801 => x"FF",
		199802 => x"FF",
		199923 => x"FF",
		199924 => x"FF",
		199925 => x"FF",
		199926 => x"FF",
		199927 => x"FF",
		200048 => x"FF",
		200049 => x"FF",
		200050 => x"FF",
		200051 => x"FF",
		200052 => x"FF",
		200173 => x"FF",
		200174 => x"FF",
		200175 => x"FF",
		200176 => x"FF",
		200177 => x"FF",
		200822 => x"FF",
		200823 => x"FF",
		200824 => x"FF",
		200825 => x"FF",
		200826 => x"FF",
		200947 => x"FF",
		200948 => x"FF",
		200949 => x"FF",
		200950 => x"FF",
		200951 => x"FF",
		201072 => x"FF",
		201073 => x"FF",
		201074 => x"FF",
		201075 => x"FF",
		201076 => x"FF",
		201197 => x"FF",
		201198 => x"FF",
		201199 => x"FF",
		201200 => x"FF",
		201201 => x"FF",
		201846 => x"FF",
		201847 => x"FF",
		201848 => x"FF",
		201849 => x"FF",
		201850 => x"FF",
		201971 => x"FF",
		201972 => x"FF",
		201973 => x"FF",
		201974 => x"FF",
		201975 => x"FF",
		202096 => x"FF",
		202097 => x"FF",
		202098 => x"FF",
		202099 => x"FF",
		202100 => x"FF",
		202221 => x"FF",
		202222 => x"FF",
		202223 => x"FF",
		202224 => x"FF",
		202225 => x"FF",
		202870 => x"FF",
		202871 => x"FF",
		202872 => x"FF",
		202873 => x"FF",
		202874 => x"FF",
		202995 => x"FF",
		202996 => x"FF",
		202997 => x"FF",
		202998 => x"FF",
		202999 => x"FF",
		203120 => x"FF",
		203121 => x"FF",
		203122 => x"FF",
		203123 => x"FF",
		203124 => x"FF",
		203245 => x"FF",
		203246 => x"FF",
		203247 => x"FF",
		203248 => x"FF",
		203249 => x"FF",
		203894 => x"FF",
		203895 => x"FF",
		203896 => x"FF",
		203897 => x"FF",
		203898 => x"FF",
		204019 => x"FF",
		204020 => x"FF",
		204021 => x"FF",
		204022 => x"FF",
		204023 => x"FF",
		204144 => x"FF",
		204145 => x"FF",
		204146 => x"FF",
		204147 => x"FF",
		204148 => x"FF",
		204269 => x"FF",
		204270 => x"FF",
		204271 => x"FF",
		204272 => x"FF",
		204273 => x"FF",
		204918 => x"FF",
		204919 => x"FF",
		204920 => x"FF",
		204921 => x"FF",
		204922 => x"FF",
		205043 => x"FF",
		205044 => x"FF",
		205045 => x"FF",
		205046 => x"FF",
		205047 => x"FF",
		205168 => x"FF",
		205169 => x"FF",
		205170 => x"FF",
		205171 => x"FF",
		205172 => x"FF",
		205293 => x"FF",
		205294 => x"FF",
		205295 => x"FF",
		205296 => x"FF",
		205297 => x"FF",
		205942 => x"FF",
		205943 => x"FF",
		205944 => x"FF",
		205945 => x"FF",
		205946 => x"FF",
		206067 => x"FF",
		206068 => x"FF",
		206069 => x"FF",
		206070 => x"FF",
		206071 => x"FF",
		206192 => x"FF",
		206193 => x"FF",
		206194 => x"FF",
		206195 => x"FF",
		206196 => x"FF",
		206317 => x"FF",
		206318 => x"FF",
		206319 => x"FF",
		206320 => x"FF",
		206321 => x"FF",
		206966 => x"FF",
		206967 => x"FF",
		206968 => x"FF",
		206969 => x"FF",
		206970 => x"FF",
		207091 => x"FF",
		207092 => x"FF",
		207093 => x"FF",
		207094 => x"FF",
		207095 => x"FF",
		207216 => x"FF",
		207217 => x"FF",
		207218 => x"FF",
		207219 => x"FF",
		207220 => x"FF",
		207341 => x"FF",
		207342 => x"FF",
		207343 => x"FF",
		207344 => x"FF",
		207345 => x"FF",
		207990 => x"FF",
		207991 => x"FF",
		207992 => x"FF",
		207993 => x"FF",
		207994 => x"FF",
		208115 => x"FF",
		208116 => x"FF",
		208117 => x"FF",
		208118 => x"FF",
		208119 => x"FF",
		208240 => x"FF",
		208241 => x"FF",
		208242 => x"FF",
		208243 => x"FF",
		208244 => x"FF",
		208365 => x"FF",
		208366 => x"FF",
		208367 => x"FF",
		208368 => x"FF",
		208369 => x"FF",
		209014 => x"FF",
		209015 => x"FF",
		209016 => x"FF",
		209017 => x"FF",
		209018 => x"FF",
		209139 => x"FF",
		209140 => x"FF",
		209141 => x"FF",
		209142 => x"FF",
		209143 => x"FF",
		209264 => x"FF",
		209265 => x"FF",
		209266 => x"FF",
		209267 => x"FF",
		209268 => x"FF",
		209389 => x"FF",
		209390 => x"FF",
		209391 => x"FF",
		209392 => x"FF",
		209393 => x"FF",
		210038 => x"FF",
		210039 => x"FF",
		210040 => x"FF",
		210041 => x"FF",
		210042 => x"FF",
		210163 => x"FF",
		210164 => x"FF",
		210165 => x"FF",
		210166 => x"FF",
		210167 => x"FF",
		210288 => x"FF",
		210289 => x"FF",
		210290 => x"FF",
		210291 => x"FF",
		210292 => x"FF",
		210413 => x"FF",
		210414 => x"FF",
		210415 => x"FF",
		210416 => x"FF",
		210417 => x"FF",
		211062 => x"FF",
		211063 => x"FF",
		211064 => x"FF",
		211065 => x"FF",
		211066 => x"FF",
		211187 => x"FF",
		211188 => x"FF",
		211189 => x"FF",
		211190 => x"FF",
		211191 => x"FF",
		211312 => x"FF",
		211313 => x"FF",
		211314 => x"FF",
		211315 => x"FF",
		211316 => x"FF",
		211437 => x"FF",
		211438 => x"FF",
		211439 => x"FF",
		211440 => x"FF",
		211441 => x"FF",
		212086 => x"FF",
		212087 => x"FF",
		212088 => x"FF",
		212089 => x"FF",
		212090 => x"FF",
		212211 => x"FF",
		212212 => x"FF",
		212213 => x"FF",
		212214 => x"FF",
		212215 => x"FF",
		212336 => x"FF",
		212337 => x"FF",
		212338 => x"FF",
		212339 => x"FF",
		212340 => x"FF",
		212461 => x"FF",
		212462 => x"FF",
		212463 => x"FF",
		212464 => x"FF",
		212465 => x"FF",
		213110 => x"FF",
		213111 => x"FF",
		213112 => x"FF",
		213113 => x"FF",
		213114 => x"FF",
		213235 => x"FF",
		213236 => x"FF",
		213237 => x"FF",
		213238 => x"FF",
		213239 => x"FF",
		213360 => x"FF",
		213361 => x"FF",
		213362 => x"FF",
		213363 => x"FF",
		213364 => x"FF",
		213485 => x"FF",
		213486 => x"FF",
		213487 => x"FF",
		213488 => x"FF",
		213489 => x"FF",
		214134 => x"FF",
		214135 => x"FF",
		214136 => x"FF",
		214137 => x"FF",
		214138 => x"FF",
		214259 => x"FF",
		214260 => x"FF",
		214261 => x"FF",
		214262 => x"FF",
		214263 => x"FF",
		214384 => x"FF",
		214385 => x"FF",
		214386 => x"FF",
		214387 => x"FF",
		214388 => x"FF",
		214509 => x"FF",
		214510 => x"FF",
		214511 => x"FF",
		214512 => x"FF",
		214513 => x"FF",
		215158 => x"FF",
		215159 => x"FF",
		215160 => x"FF",
		215161 => x"FF",
		215162 => x"FF",
		215283 => x"FF",
		215284 => x"FF",
		215285 => x"FF",
		215286 => x"FF",
		215287 => x"FF",
		215408 => x"FF",
		215409 => x"FF",
		215410 => x"FF",
		215411 => x"FF",
		215412 => x"FF",
		215533 => x"FF",
		215534 => x"FF",
		215535 => x"FF",
		215536 => x"FF",
		215537 => x"FF",
		216182 => x"FF",
		216183 => x"FF",
		216184 => x"FF",
		216185 => x"FF",
		216186 => x"FF",
		216307 => x"FF",
		216308 => x"FF",
		216309 => x"FF",
		216310 => x"FF",
		216311 => x"FF",
		216432 => x"FF",
		216433 => x"FF",
		216434 => x"FF",
		216435 => x"FF",
		216436 => x"FF",
		216557 => x"FF",
		216558 => x"FF",
		216559 => x"FF",
		216560 => x"FF",
		216561 => x"FF",
		217206 => x"FF",
		217207 => x"FF",
		217208 => x"FF",
		217209 => x"FF",
		217210 => x"FF",
		217331 => x"FF",
		217332 => x"FF",
		217333 => x"FF",
		217334 => x"FF",
		217335 => x"FF",
		217456 => x"FF",
		217457 => x"FF",
		217458 => x"FF",
		217459 => x"FF",
		217460 => x"FF",
		217581 => x"FF",
		217582 => x"FF",
		217583 => x"FF",
		217584 => x"FF",
		217585 => x"FF",
		218230 => x"FF",
		218231 => x"FF",
		218232 => x"FF",
		218233 => x"FF",
		218234 => x"FF",
		218355 => x"FF",
		218356 => x"FF",
		218357 => x"FF",
		218358 => x"FF",
		218359 => x"FF",
		218480 => x"FF",
		218481 => x"FF",
		218482 => x"FF",
		218483 => x"FF",
		218484 => x"FF",
		218605 => x"FF",
		218606 => x"FF",
		218607 => x"FF",
		218608 => x"FF",
		218609 => x"FF",
		219254 => x"FF",
		219255 => x"FF",
		219256 => x"FF",
		219257 => x"FF",
		219258 => x"FF",
		219379 => x"FF",
		219380 => x"FF",
		219381 => x"FF",
		219382 => x"FF",
		219383 => x"FF",
		219504 => x"FF",
		219505 => x"FF",
		219506 => x"FF",
		219507 => x"FF",
		219508 => x"FF",
		219629 => x"FF",
		219630 => x"FF",
		219631 => x"FF",
		219632 => x"FF",
		219633 => x"FF",
		220278 => x"FF",
		220279 => x"FF",
		220280 => x"FF",
		220281 => x"FF",
		220282 => x"FF",
		220403 => x"FF",
		220404 => x"FF",
		220405 => x"FF",
		220406 => x"FF",
		220407 => x"FF",
		220528 => x"FF",
		220529 => x"FF",
		220530 => x"FF",
		220531 => x"FF",
		220532 => x"FF",
		220653 => x"FF",
		220654 => x"FF",
		220655 => x"FF",
		220656 => x"FF",
		220657 => x"FF",
		221302 => x"FF",
		221303 => x"FF",
		221304 => x"FF",
		221305 => x"FF",
		221306 => x"FF",
		221427 => x"FF",
		221428 => x"FF",
		221429 => x"FF",
		221430 => x"FF",
		221431 => x"FF",
		221552 => x"FF",
		221553 => x"FF",
		221554 => x"FF",
		221555 => x"FF",
		221556 => x"FF",
		221677 => x"FF",
		221678 => x"FF",
		221679 => x"FF",
		221680 => x"FF",
		221681 => x"FF",
		222326 => x"FF",
		222327 => x"FF",
		222328 => x"FF",
		222329 => x"FF",
		222330 => x"FF",
		222451 => x"FF",
		222452 => x"FF",
		222453 => x"FF",
		222454 => x"FF",
		222455 => x"FF",
		222576 => x"FF",
		222577 => x"FF",
		222578 => x"FF",
		222579 => x"FF",
		222580 => x"FF",
		222701 => x"FF",
		222702 => x"FF",
		222703 => x"FF",
		222704 => x"FF",
		222705 => x"FF",
		223350 => x"FF",
		223351 => x"FF",
		223352 => x"FF",
		223353 => x"FF",
		223354 => x"FF",
		223475 => x"FF",
		223476 => x"FF",
		223477 => x"FF",
		223478 => x"FF",
		223479 => x"FF",
		223600 => x"FF",
		223601 => x"FF",
		223602 => x"FF",
		223603 => x"FF",
		223604 => x"FF",
		223725 => x"FF",
		223726 => x"FF",
		223727 => x"FF",
		223728 => x"FF",
		223729 => x"FF",
		224374 => x"FF",
		224375 => x"FF",
		224376 => x"FF",
		224377 => x"FF",
		224378 => x"FF",
		224499 => x"FF",
		224500 => x"FF",
		224501 => x"FF",
		224502 => x"FF",
		224503 => x"FF",
		224624 => x"FF",
		224625 => x"FF",
		224626 => x"FF",
		224627 => x"FF",
		224628 => x"FF",
		224749 => x"FF",
		224750 => x"FF",
		224751 => x"FF",
		224752 => x"FF",
		224753 => x"FF",
		225398 => x"FF",
		225399 => x"FF",
		225400 => x"FF",
		225401 => x"FF",
		225402 => x"FF",
		225523 => x"FF",
		225524 => x"FF",
		225525 => x"FF",
		225526 => x"FF",
		225527 => x"FF",
		225648 => x"FF",
		225649 => x"FF",
		225650 => x"FF",
		225651 => x"FF",
		225652 => x"FF",
		225773 => x"FF",
		225774 => x"FF",
		225775 => x"FF",
		225776 => x"FF",
		225777 => x"FF",
		226422 => x"FF",
		226423 => x"FF",
		226424 => x"FF",
		226425 => x"FF",
		226426 => x"FF",
		226547 => x"FF",
		226548 => x"FF",
		226549 => x"FF",
		226550 => x"FF",
		226551 => x"FF",
		226672 => x"FF",
		226673 => x"FF",
		226674 => x"FF",
		226675 => x"FF",
		226676 => x"FF",
		226797 => x"FF",
		226798 => x"FF",
		226799 => x"FF",
		226800 => x"FF",
		226801 => x"FF",
		227446 => x"FF",
		227447 => x"FF",
		227448 => x"FF",
		227449 => x"FF",
		227450 => x"FF",
		227571 => x"FF",
		227572 => x"FF",
		227573 => x"FF",
		227574 => x"FF",
		227575 => x"FF",
		227696 => x"FF",
		227697 => x"FF",
		227698 => x"FF",
		227699 => x"FF",
		227700 => x"FF",
		227821 => x"FF",
		227822 => x"FF",
		227823 => x"FF",
		227824 => x"FF",
		227825 => x"FF",
		228470 => x"FF",
		228471 => x"FF",
		228472 => x"FF",
		228473 => x"FF",
		228474 => x"FF",
		228595 => x"FF",
		228596 => x"FF",
		228597 => x"FF",
		228598 => x"FF",
		228599 => x"FF",
		228720 => x"FF",
		228721 => x"FF",
		228722 => x"FF",
		228723 => x"FF",
		228724 => x"FF",
		228845 => x"FF",
		228846 => x"FF",
		228847 => x"FF",
		228848 => x"FF",
		228849 => x"FF",
		229494 => x"FF",
		229495 => x"FF",
		229496 => x"FF",
		229497 => x"FF",
		229498 => x"FF",
		229619 => x"FF",
		229620 => x"FF",
		229621 => x"FF",
		229622 => x"FF",
		229623 => x"FF",
		229744 => x"FF",
		229745 => x"FF",
		229746 => x"FF",
		229747 => x"FF",
		229748 => x"FF",
		229869 => x"FF",
		229870 => x"FF",
		229871 => x"FF",
		229872 => x"FF",
		229873 => x"FF",
		230518 => x"FF",
		230519 => x"FF",
		230520 => x"FF",
		230521 => x"FF",
		230522 => x"FF",
		230643 => x"FF",
		230644 => x"FF",
		230645 => x"FF",
		230646 => x"FF",
		230647 => x"FF",
		230768 => x"FF",
		230769 => x"FF",
		230770 => x"FF",
		230771 => x"FF",
		230772 => x"FF",
		230893 => x"FF",
		230894 => x"FF",
		230895 => x"FF",
		230896 => x"FF",
		230897 => x"FF",
		231542 => x"FF",
		231543 => x"FF",
		231544 => x"FF",
		231545 => x"FF",
		231546 => x"FF",
		231667 => x"FF",
		231668 => x"FF",
		231669 => x"FF",
		231670 => x"FF",
		231671 => x"FF",
		231792 => x"FF",
		231793 => x"FF",
		231794 => x"FF",
		231795 => x"FF",
		231796 => x"FF",
		231917 => x"FF",
		231918 => x"FF",
		231919 => x"FF",
		231920 => x"FF",
		231921 => x"FF",
		232566 => x"FF",
		232567 => x"FF",
		232568 => x"FF",
		232569 => x"FF",
		232570 => x"FF",
		232691 => x"FF",
		232692 => x"FF",
		232693 => x"FF",
		232694 => x"FF",
		232695 => x"FF",
		232816 => x"FF",
		232817 => x"FF",
		232818 => x"FF",
		232819 => x"FF",
		232820 => x"FF",
		232941 => x"FF",
		232942 => x"FF",
		232943 => x"FF",
		232944 => x"FF",
		232945 => x"FF",
		233590 => x"FF",
		233591 => x"FF",
		233592 => x"FF",
		233593 => x"FF",
		233594 => x"FF",
		233715 => x"FF",
		233716 => x"FF",
		233717 => x"FF",
		233718 => x"FF",
		233719 => x"FF",
		233840 => x"FF",
		233841 => x"FF",
		233842 => x"FF",
		233843 => x"FF",
		233844 => x"FF",
		233965 => x"FF",
		233966 => x"FF",
		233967 => x"FF",
		233968 => x"FF",
		233969 => x"FF",
		234614 => x"FF",
		234615 => x"FF",
		234616 => x"FF",
		234617 => x"FF",
		234618 => x"FF",
		234739 => x"FF",
		234740 => x"FF",
		234741 => x"FF",
		234742 => x"FF",
		234743 => x"FF",
		234864 => x"FF",
		234865 => x"FF",
		234866 => x"FF",
		234867 => x"FF",
		234868 => x"FF",
		234989 => x"FF",
		234990 => x"FF",
		234991 => x"FF",
		234992 => x"FF",
		234993 => x"FF",
		235638 => x"FF",
		235639 => x"FF",
		235640 => x"FF",
		235641 => x"FF",
		235642 => x"FF",
		235763 => x"FF",
		235764 => x"FF",
		235765 => x"FF",
		235766 => x"FF",
		235767 => x"FF",
		235888 => x"FF",
		235889 => x"FF",
		235890 => x"FF",
		235891 => x"FF",
		235892 => x"FF",
		236013 => x"FF",
		236014 => x"FF",
		236015 => x"FF",
		236016 => x"FF",
		236017 => x"FF",
		236662 => x"FF",
		236663 => x"FF",
		236664 => x"FF",
		236665 => x"FF",
		236666 => x"FF",
		236787 => x"FF",
		236788 => x"FF",
		236789 => x"FF",
		236790 => x"FF",
		236791 => x"FF",
		236912 => x"FF",
		236913 => x"FF",
		236914 => x"FF",
		236915 => x"FF",
		236916 => x"FF",
		237037 => x"FF",
		237038 => x"FF",
		237039 => x"FF",
		237040 => x"FF",
		237041 => x"FF",
		237686 => x"FF",
		237687 => x"FF",
		237688 => x"FF",
		237689 => x"FF",
		237690 => x"FF",
		237811 => x"FF",
		237812 => x"FF",
		237813 => x"FF",
		237814 => x"FF",
		237815 => x"FF",
		237936 => x"FF",
		237937 => x"FF",
		237938 => x"FF",
		237939 => x"FF",
		237940 => x"FF",
		238061 => x"FF",
		238062 => x"FF",
		238063 => x"FF",
		238064 => x"FF",
		238065 => x"FF",
		238710 => x"FF",
		238711 => x"FF",
		238712 => x"FF",
		238713 => x"FF",
		238714 => x"FF",
		238835 => x"FF",
		238836 => x"FF",
		238837 => x"FF",
		238838 => x"FF",
		238839 => x"FF",
		238960 => x"FF",
		238961 => x"FF",
		238962 => x"FF",
		238963 => x"FF",
		238964 => x"FF",
		239085 => x"FF",
		239086 => x"FF",
		239087 => x"FF",
		239088 => x"FF",
		239089 => x"FF",
		239734 => x"FF",
		239735 => x"FF",
		239736 => x"FF",
		239737 => x"FF",
		239738 => x"FF",
		239859 => x"FF",
		239860 => x"FF",
		239861 => x"FF",
		239862 => x"FF",
		239863 => x"FF",
		239984 => x"FF",
		239985 => x"FF",
		239986 => x"FF",
		239987 => x"FF",
		239988 => x"FF",
		240109 => x"FF",
		240110 => x"FF",
		240111 => x"FF",
		240112 => x"FF",
		240113 => x"FF",
		240758 => x"FF",
		240759 => x"FF",
		240760 => x"FF",
		240761 => x"FF",
		240762 => x"FF",
		240883 => x"FF",
		240884 => x"FF",
		240885 => x"FF",
		240886 => x"FF",
		240887 => x"FF",
		241008 => x"FF",
		241009 => x"FF",
		241010 => x"FF",
		241011 => x"FF",
		241012 => x"FF",
		241133 => x"FF",
		241134 => x"FF",
		241135 => x"FF",
		241136 => x"FF",
		241137 => x"FF",
		241782 => x"FF",
		241783 => x"FF",
		241784 => x"FF",
		241785 => x"FF",
		241786 => x"FF",
		241907 => x"FF",
		241908 => x"FF",
		241909 => x"FF",
		241910 => x"FF",
		241911 => x"FF",
		242032 => x"FF",
		242033 => x"FF",
		242034 => x"FF",
		242035 => x"FF",
		242036 => x"FF",
		242157 => x"FF",
		242158 => x"FF",
		242159 => x"FF",
		242160 => x"FF",
		242161 => x"FF",
		242806 => x"FF",
		242807 => x"FF",
		242808 => x"FF",
		242809 => x"FF",
		242810 => x"FF",
		242931 => x"FF",
		242932 => x"FF",
		242933 => x"FF",
		242934 => x"FF",
		242935 => x"FF",
		243056 => x"FF",
		243057 => x"FF",
		243058 => x"FF",
		243059 => x"FF",
		243060 => x"FF",
		243181 => x"FF",
		243182 => x"FF",
		243183 => x"FF",
		243184 => x"FF",
		243185 => x"FF",
		243830 => x"FF",
		243831 => x"FF",
		243832 => x"FF",
		243833 => x"FF",
		243834 => x"FF",
		243955 => x"FF",
		243956 => x"FF",
		243957 => x"FF",
		243958 => x"FF",
		243959 => x"FF",
		244080 => x"FF",
		244081 => x"FF",
		244082 => x"FF",
		244083 => x"FF",
		244084 => x"FF",
		244205 => x"FF",
		244206 => x"FF",
		244207 => x"FF",
		244208 => x"FF",
		244209 => x"FF",
		244854 => x"FF",
		244855 => x"FF",
		244856 => x"FF",
		244857 => x"FF",
		244858 => x"FF",
		244979 => x"FF",
		244980 => x"FF",
		244981 => x"FF",
		244982 => x"FF",
		244983 => x"FF",
		245104 => x"FF",
		245105 => x"FF",
		245106 => x"FF",
		245107 => x"FF",
		245108 => x"FF",
		245229 => x"FF",
		245230 => x"FF",
		245231 => x"FF",
		245232 => x"FF",
		245233 => x"FF",
		245878 => x"FF",
		245879 => x"FF",
		245880 => x"FF",
		245881 => x"FF",
		245882 => x"FF",
		246003 => x"FF",
		246004 => x"FF",
		246005 => x"FF",
		246006 => x"FF",
		246007 => x"FF",
		246128 => x"FF",
		246129 => x"FF",
		246130 => x"FF",
		246131 => x"FF",
		246132 => x"FF",
		246253 => x"FF",
		246254 => x"FF",
		246255 => x"FF",
		246256 => x"FF",
		246257 => x"FF",
		246902 => x"FF",
		246903 => x"FF",
		246904 => x"FF",
		246905 => x"FF",
		246906 => x"FF",
		247027 => x"FF",
		247028 => x"FF",
		247029 => x"FF",
		247030 => x"FF",
		247031 => x"FF",
		247152 => x"FF",
		247153 => x"FF",
		247154 => x"FF",
		247155 => x"FF",
		247156 => x"FF",
		247277 => x"FF",
		247278 => x"FF",
		247279 => x"FF",
		247280 => x"FF",
		247281 => x"FF",
		247926 => x"FF",
		247927 => x"FF",
		247928 => x"FF",
		247929 => x"FF",
		247930 => x"FF",
		248051 => x"FF",
		248052 => x"FF",
		248053 => x"FF",
		248054 => x"FF",
		248055 => x"FF",
		248176 => x"FF",
		248177 => x"FF",
		248178 => x"FF",
		248179 => x"FF",
		248180 => x"FF",
		248301 => x"FF",
		248302 => x"FF",
		248303 => x"FF",
		248304 => x"FF",
		248305 => x"FF",
		248950 => x"FF",
		248951 => x"FF",
		248952 => x"FF",
		248953 => x"FF",
		248954 => x"FF",
		249075 => x"FF",
		249076 => x"FF",
		249077 => x"FF",
		249078 => x"FF",
		249079 => x"FF",
		249200 => x"FF",
		249201 => x"FF",
		249202 => x"FF",
		249203 => x"FF",
		249204 => x"FF",
		249325 => x"FF",
		249326 => x"FF",
		249327 => x"FF",
		249328 => x"FF",
		249329 => x"FF",
		249974 => x"FF",
		249975 => x"FF",
		249976 => x"FF",
		249977 => x"FF",
		249978 => x"FF",
		250099 => x"FF",
		250100 => x"FF",
		250101 => x"FF",
		250102 => x"FF",
		250103 => x"FF",
		250224 => x"FF",
		250225 => x"FF",
		250226 => x"FF",
		250227 => x"FF",
		250228 => x"FF",
		250349 => x"FF",
		250350 => x"FF",
		250351 => x"FF",
		250352 => x"FF",
		250353 => x"FF",
		250998 => x"FF",
		250999 => x"FF",
		251000 => x"FF",
		251001 => x"FF",
		251002 => x"FF",
		251123 => x"FF",
		251124 => x"FF",
		251125 => x"FF",
		251126 => x"FF",
		251127 => x"FF",
		251248 => x"FF",
		251249 => x"FF",
		251250 => x"FF",
		251251 => x"FF",
		251252 => x"FF",
		251373 => x"FF",
		251374 => x"FF",
		251375 => x"FF",
		251376 => x"FF",
		251377 => x"FF",
		252022 => x"FF",
		252023 => x"FF",
		252024 => x"FF",
		252025 => x"FF",
		252026 => x"FF",
		252147 => x"FF",
		252148 => x"FF",
		252149 => x"FF",
		252150 => x"FF",
		252151 => x"FF",
		252272 => x"FF",
		252273 => x"FF",
		252274 => x"FF",
		252275 => x"FF",
		252276 => x"FF",
		252397 => x"FF",
		252398 => x"FF",
		252399 => x"FF",
		252400 => x"FF",
		252401 => x"FF",
		253046 => x"FF",
		253047 => x"FF",
		253048 => x"FF",
		253049 => x"FF",
		253050 => x"FF",
		253171 => x"FF",
		253172 => x"FF",
		253173 => x"FF",
		253174 => x"FF",
		253175 => x"FF",
		253296 => x"FF",
		253297 => x"FF",
		253298 => x"FF",
		253299 => x"FF",
		253300 => x"FF",
		253421 => x"FF",
		253422 => x"FF",
		253423 => x"FF",
		253424 => x"FF",
		253425 => x"FF",
		254070 => x"FF",
		254071 => x"FF",
		254072 => x"FF",
		254073 => x"FF",
		254074 => x"FF",
		254195 => x"FF",
		254196 => x"FF",
		254197 => x"FF",
		254198 => x"FF",
		254199 => x"FF",
		254320 => x"FF",
		254321 => x"FF",
		254322 => x"FF",
		254323 => x"FF",
		254324 => x"FF",
		254445 => x"FF",
		254446 => x"FF",
		254447 => x"FF",
		254448 => x"FF",
		254449 => x"FF",
		255094 => x"FF",
		255095 => x"FF",
		255096 => x"FF",
		255097 => x"FF",
		255098 => x"FF",
		255219 => x"FF",
		255220 => x"FF",
		255221 => x"FF",
		255222 => x"FF",
		255223 => x"FF",
		255344 => x"FF",
		255345 => x"FF",
		255346 => x"FF",
		255347 => x"FF",
		255348 => x"FF",
		255469 => x"FF",
		255470 => x"FF",
		255471 => x"FF",
		255472 => x"FF",
		255473 => x"FF",
		256118 => x"FF",
		256119 => x"FF",
		256120 => x"FF",
		256121 => x"FF",
		256122 => x"FF",
		256243 => x"FF",
		256244 => x"FF",
		256245 => x"FF",
		256246 => x"FF",
		256247 => x"FF",
		256368 => x"FF",
		256369 => x"FF",
		256370 => x"FF",
		256371 => x"FF",
		256372 => x"FF",
		256493 => x"FF",
		256494 => x"FF",
		256495 => x"FF",
		256496 => x"FF",
		256497 => x"FF",
		257142 => x"FF",
		257143 => x"FF",
		257144 => x"FF",
		257145 => x"FF",
		257146 => x"FF",
		257267 => x"FF",
		257268 => x"FF",
		257269 => x"FF",
		257270 => x"FF",
		257271 => x"FF",
		257392 => x"FF",
		257393 => x"FF",
		257394 => x"FF",
		257395 => x"FF",
		257396 => x"FF",
		257517 => x"FF",
		257518 => x"FF",
		257519 => x"FF",
		257520 => x"FF",
		257521 => x"FF",
		258166 => x"FF",
		258167 => x"FF",
		258168 => x"FF",
		258169 => x"FF",
		258170 => x"FF",
		258291 => x"FF",
		258292 => x"FF",
		258293 => x"FF",
		258294 => x"FF",
		258295 => x"FF",
		258416 => x"FF",
		258417 => x"FF",
		258418 => x"FF",
		258419 => x"FF",
		258420 => x"FF",
		258541 => x"FF",
		258542 => x"FF",
		258543 => x"FF",
		258544 => x"FF",
		258545 => x"FF",
		259190 => x"FF",
		259191 => x"FF",
		259192 => x"FF",
		259193 => x"FF",
		259194 => x"FF",
		259315 => x"FF",
		259316 => x"FF",
		259317 => x"FF",
		259318 => x"FF",
		259319 => x"FF",
		259440 => x"FF",
		259441 => x"FF",
		259442 => x"FF",
		259443 => x"FF",
		259444 => x"FF",
		259565 => x"FF",
		259566 => x"FF",
		259567 => x"FF",
		259568 => x"FF",
		259569 => x"FF",
		260214 => x"FF",
		260215 => x"FF",
		260216 => x"FF",
		260217 => x"FF",
		260218 => x"FF",
		260339 => x"FF",
		260340 => x"FF",
		260341 => x"FF",
		260342 => x"FF",
		260343 => x"FF",
		260464 => x"FF",
		260465 => x"FF",
		260466 => x"FF",
		260467 => x"FF",
		260468 => x"FF",
		260589 => x"FF",
		260590 => x"FF",
		260591 => x"FF",
		260592 => x"FF",
		260593 => x"FF",
		261238 => x"FF",
		261239 => x"FF",
		261240 => x"FF",
		261241 => x"FF",
		261242 => x"FF",
		261363 => x"FF",
		261364 => x"FF",
		261365 => x"FF",
		261366 => x"FF",
		261367 => x"FF",
		261488 => x"FF",
		261489 => x"FF",
		261490 => x"FF",
		261491 => x"FF",
		261492 => x"FF",
		261613 => x"FF",
		261614 => x"FF",
		261615 => x"FF",
		261616 => x"FF",
		261617 => x"FF",
		262262 => x"FF",
		262263 => x"FF",
		262264 => x"FF",
		262265 => x"FF",
		262266 => x"FF",
		262387 => x"FF",
		262388 => x"FF",
		262389 => x"FF",
		262390 => x"FF",
		262391 => x"FF",
		262512 => x"FF",
		262513 => x"FF",
		262514 => x"FF",
		262515 => x"FF",
		262516 => x"FF",
		262637 => x"FF",
		262638 => x"FF",
		262639 => x"FF",
		262640 => x"FF",
		262641 => x"FF",
		263286 => x"FF",
		263287 => x"FF",
		263288 => x"FF",
		263289 => x"FF",
		263290 => x"FF",
		263411 => x"FF",
		263412 => x"FF",
		263413 => x"FF",
		263414 => x"FF",
		263415 => x"FF",
		263536 => x"FF",
		263537 => x"FF",
		263538 => x"FF",
		263539 => x"FF",
		263540 => x"FF",
		263661 => x"FF",
		263662 => x"FF",
		263663 => x"FF",
		263664 => x"FF",
		263665 => x"FF",
		264310 => x"FF",
		264311 => x"FF",
		264312 => x"FF",
		264313 => x"FF",
		264314 => x"FF",
		264435 => x"FF",
		264436 => x"FF",
		264437 => x"FF",
		264438 => x"FF",
		264439 => x"FF",
		264560 => x"FF",
		264561 => x"FF",
		264562 => x"FF",
		264563 => x"FF",
		264564 => x"FF",
		264685 => x"FF",
		264686 => x"FF",
		264687 => x"FF",
		264688 => x"FF",
		264689 => x"FF",
		265334 => x"FF",
		265335 => x"FF",
		265336 => x"FF",
		265337 => x"FF",
		265338 => x"FF",
		265459 => x"FF",
		265460 => x"FF",
		265461 => x"FF",
		265462 => x"FF",
		265463 => x"FF",
		265584 => x"FF",
		265585 => x"FF",
		265586 => x"FF",
		265587 => x"FF",
		265588 => x"FF",
		265709 => x"FF",
		265710 => x"FF",
		265711 => x"FF",
		265712 => x"FF",
		265713 => x"FF",
		266358 => x"FF",
		266359 => x"FF",
		266360 => x"FF",
		266361 => x"FF",
		266362 => x"FF",
		266483 => x"FF",
		266484 => x"FF",
		266485 => x"FF",
		266486 => x"FF",
		266487 => x"FF",
		266608 => x"FF",
		266609 => x"FF",
		266610 => x"FF",
		266611 => x"FF",
		266612 => x"FF",
		266733 => x"FF",
		266734 => x"FF",
		266735 => x"FF",
		266736 => x"FF",
		266737 => x"FF",
		267382 => x"FF",
		267383 => x"FF",
		267384 => x"FF",
		267385 => x"FF",
		267386 => x"FF",
		267507 => x"FF",
		267508 => x"FF",
		267509 => x"FF",
		267510 => x"FF",
		267511 => x"FF",
		267632 => x"FF",
		267633 => x"FF",
		267634 => x"FF",
		267635 => x"FF",
		267636 => x"FF",
		267757 => x"FF",
		267758 => x"FF",
		267759 => x"FF",
		267760 => x"FF",
		267761 => x"FF",
		268406 => x"FF",
		268407 => x"FF",
		268408 => x"FF",
		268409 => x"FF",
		268410 => x"FF",
		268531 => x"FF",
		268532 => x"FF",
		268533 => x"FF",
		268534 => x"FF",
		268535 => x"FF",
		268656 => x"FF",
		268657 => x"FF",
		268658 => x"FF",
		268659 => x"FF",
		268660 => x"FF",
		268781 => x"FF",
		268782 => x"FF",
		268783 => x"FF",
		268784 => x"FF",
		268785 => x"FF",
		269430 => x"FF",
		269431 => x"FF",
		269432 => x"FF",
		269433 => x"FF",
		269434 => x"FF",
		269555 => x"FF",
		269556 => x"FF",
		269557 => x"FF",
		269558 => x"FF",
		269559 => x"FF",
		269680 => x"FF",
		269681 => x"FF",
		269682 => x"FF",
		269683 => x"FF",
		269684 => x"FF",
		269805 => x"FF",
		269806 => x"FF",
		269807 => x"FF",
		269808 => x"FF",
		269809 => x"FF",
		270454 => x"FF",
		270455 => x"FF",
		270456 => x"FF",
		270457 => x"FF",
		270458 => x"FF",
		270579 => x"FF",
		270580 => x"FF",
		270581 => x"FF",
		270582 => x"FF",
		270583 => x"FF",
		270704 => x"FF",
		270705 => x"FF",
		270706 => x"FF",
		270707 => x"FF",
		270708 => x"FF",
		270829 => x"FF",
		270830 => x"FF",
		270831 => x"FF",
		270832 => x"FF",
		270833 => x"FF",
		271478 => x"FF",
		271479 => x"FF",
		271480 => x"FF",
		271481 => x"FF",
		271482 => x"FF",
		271603 => x"FF",
		271604 => x"FF",
		271605 => x"FF",
		271606 => x"FF",
		271607 => x"FF",
		271728 => x"FF",
		271729 => x"FF",
		271730 => x"FF",
		271731 => x"FF",
		271732 => x"FF",
		271853 => x"FF",
		271854 => x"FF",
		271855 => x"FF",
		271856 => x"FF",
		271857 => x"FF",
		272502 => x"FF",
		272503 => x"FF",
		272504 => x"FF",
		272505 => x"FF",
		272506 => x"FF",
		272627 => x"FF",
		272628 => x"FF",
		272629 => x"FF",
		272630 => x"FF",
		272631 => x"FF",
		272752 => x"FF",
		272753 => x"FF",
		272754 => x"FF",
		272755 => x"FF",
		272756 => x"FF",
		272877 => x"FF",
		272878 => x"FF",
		272879 => x"FF",
		272880 => x"FF",
		272881 => x"FF",
		273526 => x"FF",
		273527 => x"FF",
		273528 => x"FF",
		273529 => x"FF",
		273530 => x"FF",
		273651 => x"FF",
		273652 => x"FF",
		273653 => x"FF",
		273654 => x"FF",
		273655 => x"FF",
		273776 => x"FF",
		273777 => x"FF",
		273778 => x"FF",
		273779 => x"FF",
		273780 => x"FF",
		273901 => x"FF",
		273902 => x"FF",
		273903 => x"FF",
		273904 => x"FF",
		273905 => x"FF",
		274550 => x"FF",
		274551 => x"FF",
		274552 => x"FF",
		274553 => x"FF",
		274554 => x"FF",
		274675 => x"FF",
		274676 => x"FF",
		274677 => x"FF",
		274678 => x"FF",
		274679 => x"FF",
		274800 => x"FF",
		274801 => x"FF",
		274802 => x"FF",
		274803 => x"FF",
		274804 => x"FF",
		274925 => x"FF",
		274926 => x"FF",
		274927 => x"FF",
		274928 => x"FF",
		274929 => x"FF",
		275574 => x"FF",
		275575 => x"FF",
		275576 => x"FF",
		275577 => x"FF",
		275578 => x"FF",
		275699 => x"FF",
		275700 => x"FF",
		275701 => x"FF",
		275702 => x"FF",
		275703 => x"FF",
		275824 => x"FF",
		275825 => x"FF",
		275826 => x"FF",
		275827 => x"FF",
		275828 => x"FF",
		275949 => x"FF",
		275950 => x"FF",
		275951 => x"FF",
		275952 => x"FF",
		275953 => x"FF",
		276598 => x"FF",
		276599 => x"FF",
		276600 => x"FF",
		276601 => x"FF",
		276602 => x"FF",
		276723 => x"FF",
		276724 => x"FF",
		276725 => x"FF",
		276726 => x"FF",
		276727 => x"FF",
		276848 => x"FF",
		276849 => x"FF",
		276850 => x"FF",
		276851 => x"FF",
		276852 => x"FF",
		276973 => x"FF",
		276974 => x"FF",
		276975 => x"FF",
		276976 => x"FF",
		276977 => x"FF",
		277622 => x"FF",
		277623 => x"FF",
		277624 => x"FF",
		277625 => x"FF",
		277626 => x"FF",
		277747 => x"FF",
		277748 => x"FF",
		277749 => x"FF",
		277750 => x"FF",
		277751 => x"FF",
		277872 => x"FF",
		277873 => x"FF",
		277874 => x"FF",
		277875 => x"FF",
		277876 => x"FF",
		277997 => x"FF",
		277998 => x"FF",
		277999 => x"FF",
		278000 => x"FF",
		278001 => x"FF",
		278646 => x"FF",
		278647 => x"FF",
		278648 => x"FF",
		278649 => x"FF",
		278650 => x"FF",
		278771 => x"FF",
		278772 => x"FF",
		278773 => x"FF",
		278774 => x"FF",
		278775 => x"FF",
		278896 => x"FF",
		278897 => x"FF",
		278898 => x"FF",
		278899 => x"FF",
		278900 => x"FF",
		279021 => x"FF",
		279022 => x"FF",
		279023 => x"FF",
		279024 => x"FF",
		279025 => x"FF",
		279670 => x"FF",
		279671 => x"FF",
		279672 => x"FF",
		279673 => x"FF",
		279674 => x"FF",
		279795 => x"FF",
		279796 => x"FF",
		279797 => x"FF",
		279798 => x"FF",
		279799 => x"FF",
		279920 => x"FF",
		279921 => x"FF",
		279922 => x"FF",
		279923 => x"FF",
		279924 => x"FF",
		280045 => x"FF",
		280046 => x"FF",
		280047 => x"FF",
		280048 => x"FF",
		280049 => x"FF",
		280694 => x"FF",
		280695 => x"FF",
		280696 => x"FF",
		280697 => x"FF",
		280698 => x"FF",
		280819 => x"FF",
		280820 => x"FF",
		280821 => x"FF",
		280822 => x"FF",
		280823 => x"FF",
		280944 => x"FF",
		280945 => x"FF",
		280946 => x"FF",
		280947 => x"FF",
		280948 => x"FF",
		281069 => x"FF",
		281070 => x"FF",
		281071 => x"FF",
		281072 => x"FF",
		281073 => x"FF",
		281718 => x"FF",
		281719 => x"FF",
		281720 => x"FF",
		281721 => x"FF",
		281722 => x"FF",
		281843 => x"FF",
		281844 => x"FF",
		281845 => x"FF",
		281846 => x"FF",
		281847 => x"FF",
		281968 => x"FF",
		281969 => x"FF",
		281970 => x"FF",
		281971 => x"FF",
		281972 => x"FF",
		282093 => x"FF",
		282094 => x"FF",
		282095 => x"FF",
		282096 => x"FF",
		282097 => x"FF",
		282742 => x"FF",
		282743 => x"FF",
		282744 => x"FF",
		282745 => x"FF",
		282746 => x"FF",
		282867 => x"FF",
		282868 => x"FF",
		282869 => x"FF",
		282870 => x"FF",
		282871 => x"FF",
		282992 => x"FF",
		282993 => x"FF",
		282994 => x"FF",
		282995 => x"FF",
		282996 => x"FF",
		283117 => x"FF",
		283118 => x"FF",
		283119 => x"FF",
		283120 => x"FF",
		283121 => x"FF",
		283766 => x"FF",
		283767 => x"FF",
		283768 => x"FF",
		283769 => x"FF",
		283770 => x"FF",
		283891 => x"FF",
		283892 => x"FF",
		283893 => x"FF",
		283894 => x"FF",
		283895 => x"FF",
		284016 => x"FF",
		284017 => x"FF",
		284018 => x"FF",
		284019 => x"FF",
		284020 => x"FF",
		284141 => x"FF",
		284142 => x"FF",
		284143 => x"FF",
		284144 => x"FF",
		284145 => x"FF",
		284790 => x"FF",
		284791 => x"FF",
		284792 => x"FF",
		284793 => x"FF",
		284794 => x"FF",
		284915 => x"FF",
		284916 => x"FF",
		284917 => x"FF",
		284918 => x"FF",
		284919 => x"FF",
		285040 => x"FF",
		285041 => x"FF",
		285042 => x"FF",
		285043 => x"FF",
		285044 => x"FF",
		285165 => x"FF",
		285166 => x"FF",
		285167 => x"FF",
		285168 => x"FF",
		285169 => x"FF",
		285814 => x"FF",
		285815 => x"FF",
		285816 => x"FF",
		285817 => x"FF",
		285818 => x"FF",
		285939 => x"FF",
		285940 => x"FF",
		285941 => x"FF",
		285942 => x"FF",
		285943 => x"FF",
		286064 => x"FF",
		286065 => x"FF",
		286066 => x"FF",
		286067 => x"FF",
		286068 => x"FF",
		286189 => x"FF",
		286190 => x"FF",
		286191 => x"FF",
		286192 => x"FF",
		286193 => x"FF",
		286838 => x"FF",
		286839 => x"FF",
		286840 => x"FF",
		286841 => x"FF",
		286842 => x"FF",
		286963 => x"FF",
		286964 => x"FF",
		286965 => x"FF",
		286966 => x"FF",
		286967 => x"FF",
		287088 => x"FF",
		287089 => x"FF",
		287090 => x"FF",
		287091 => x"FF",
		287092 => x"FF",
		287213 => x"FF",
		287214 => x"FF",
		287215 => x"FF",
		287216 => x"FF",
		287217 => x"FF",
		287862 => x"FF",
		287863 => x"FF",
		287864 => x"FF",
		287865 => x"FF",
		287866 => x"FF",
		287987 => x"FF",
		287988 => x"FF",
		287989 => x"FF",
		287990 => x"FF",
		287991 => x"FF",
		288112 => x"FF",
		288113 => x"FF",
		288114 => x"FF",
		288115 => x"FF",
		288116 => x"FF",
		288237 => x"FF",
		288238 => x"FF",
		288239 => x"FF",
		288240 => x"FF",
		288241 => x"FF",
		288886 => x"FF",
		288887 => x"FF",
		288888 => x"FF",
		288889 => x"FF",
		288890 => x"FF",
		289011 => x"FF",
		289012 => x"FF",
		289013 => x"FF",
		289014 => x"FF",
		289015 => x"FF",
		289136 => x"FF",
		289137 => x"FF",
		289138 => x"FF",
		289139 => x"FF",
		289140 => x"FF",
		289261 => x"FF",
		289262 => x"FF",
		289263 => x"FF",
		289264 => x"FF",
		289265 => x"FF",
		289910 => x"FF",
		289911 => x"FF",
		289912 => x"FF",
		289913 => x"FF",
		289914 => x"FF",
		290035 => x"FF",
		290036 => x"FF",
		290037 => x"FF",
		290038 => x"FF",
		290039 => x"FF",
		290160 => x"FF",
		290161 => x"FF",
		290162 => x"FF",
		290163 => x"FF",
		290164 => x"FF",
		290285 => x"FF",
		290286 => x"FF",
		290287 => x"FF",
		290288 => x"FF",
		290289 => x"FF",
		290934 => x"FF",
		290935 => x"FF",
		290936 => x"FF",
		290937 => x"FF",
		290938 => x"FF",
		291059 => x"FF",
		291060 => x"FF",
		291061 => x"FF",
		291062 => x"FF",
		291063 => x"FF",
		291184 => x"FF",
		291185 => x"FF",
		291186 => x"FF",
		291187 => x"FF",
		291188 => x"FF",
		291309 => x"FF",
		291310 => x"FF",
		291311 => x"FF",
		291312 => x"FF",
		291313 => x"FF",
		291958 => x"FF",
		291959 => x"FF",
		291960 => x"FF",
		291961 => x"FF",
		291962 => x"FF",
		292083 => x"FF",
		292084 => x"FF",
		292085 => x"FF",
		292086 => x"FF",
		292087 => x"FF",
		292208 => x"FF",
		292209 => x"FF",
		292210 => x"FF",
		292211 => x"FF",
		292212 => x"FF",
		292333 => x"FF",
		292334 => x"FF",
		292335 => x"FF",
		292336 => x"FF",
		292337 => x"FF",
		292982 => x"FF",
		292983 => x"FF",
		292984 => x"FF",
		292985 => x"FF",
		292986 => x"FF",
		293107 => x"FF",
		293108 => x"FF",
		293109 => x"FF",
		293110 => x"FF",
		293111 => x"FF",
		293232 => x"FF",
		293233 => x"FF",
		293234 => x"FF",
		293235 => x"FF",
		293236 => x"FF",
		293357 => x"FF",
		293358 => x"FF",
		293359 => x"FF",
		293360 => x"FF",
		293361 => x"FF",
		294006 => x"FF",
		294007 => x"FF",
		294008 => x"FF",
		294009 => x"FF",
		294010 => x"FF",
		294131 => x"FF",
		294132 => x"FF",
		294133 => x"FF",
		294134 => x"FF",
		294135 => x"FF",
		294256 => x"FF",
		294257 => x"FF",
		294258 => x"FF",
		294259 => x"FF",
		294260 => x"FF",
		294381 => x"FF",
		294382 => x"FF",
		294383 => x"FF",
		294384 => x"FF",
		294385 => x"FF",
		295030 => x"FF",
		295031 => x"FF",
		295032 => x"FF",
		295033 => x"FF",
		295034 => x"FF",
		295155 => x"FF",
		295156 => x"FF",
		295157 => x"FF",
		295158 => x"FF",
		295159 => x"FF",
		295280 => x"FF",
		295281 => x"FF",
		295282 => x"FF",
		295283 => x"FF",
		295284 => x"FF",
		295405 => x"FF",
		295406 => x"FF",
		295407 => x"FF",
		295408 => x"FF",
		295409 => x"FF",
		296054 => x"FF",
		296055 => x"FF",
		296056 => x"FF",
		296057 => x"FF",
		296058 => x"FF",
		296179 => x"FF",
		296180 => x"FF",
		296181 => x"FF",
		296182 => x"FF",
		296183 => x"FF",
		296304 => x"FF",
		296305 => x"FF",
		296306 => x"FF",
		296307 => x"FF",
		296308 => x"FF",
		296429 => x"FF",
		296430 => x"FF",
		296431 => x"FF",
		296432 => x"FF",
		296433 => x"FF",
		297078 => x"FF",
		297079 => x"FF",
		297080 => x"FF",
		297081 => x"FF",
		297082 => x"FF",
		297203 => x"FF",
		297204 => x"FF",
		297205 => x"FF",
		297206 => x"FF",
		297207 => x"FF",
		297328 => x"FF",
		297329 => x"FF",
		297330 => x"FF",
		297331 => x"FF",
		297332 => x"FF",
		297453 => x"FF",
		297454 => x"FF",
		297455 => x"FF",
		297456 => x"FF",
		297457 => x"FF",
		298102 => x"FF",
		298103 => x"FF",
		298104 => x"FF",
		298105 => x"FF",
		298106 => x"FF",
		298227 => x"FF",
		298228 => x"FF",
		298229 => x"FF",
		298230 => x"FF",
		298231 => x"FF",
		298352 => x"FF",
		298353 => x"FF",
		298354 => x"FF",
		298355 => x"FF",
		298356 => x"FF",
		298477 => x"FF",
		298478 => x"FF",
		298479 => x"FF",
		298480 => x"FF",
		298481 => x"FF",
		299126 => x"FF",
		299127 => x"FF",
		299128 => x"FF",
		299129 => x"FF",
		299130 => x"FF",
		299251 => x"FF",
		299252 => x"FF",
		299253 => x"FF",
		299254 => x"FF",
		299255 => x"FF",
		299376 => x"FF",
		299377 => x"FF",
		299378 => x"FF",
		299379 => x"FF",
		299380 => x"FF",
		299501 => x"FF",
		299502 => x"FF",
		299503 => x"FF",
		299504 => x"FF",
		299505 => x"FF",
		300150 => x"FF",
		300151 => x"FF",
		300152 => x"FF",
		300153 => x"FF",
		300154 => x"FF",
		300275 => x"FF",
		300276 => x"FF",
		300277 => x"FF",
		300278 => x"FF",
		300279 => x"FF",
		300400 => x"FF",
		300401 => x"FF",
		300402 => x"FF",
		300403 => x"FF",
		300404 => x"FF",
		300525 => x"FF",
		300526 => x"FF",
		300527 => x"FF",
		300528 => x"FF",
		300529 => x"FF",
		301174 => x"FF",
		301175 => x"FF",
		301176 => x"FF",
		301177 => x"FF",
		301178 => x"FF",
		301299 => x"FF",
		301300 => x"FF",
		301301 => x"FF",
		301302 => x"FF",
		301303 => x"FF",
		301424 => x"FF",
		301425 => x"FF",
		301426 => x"FF",
		301427 => x"FF",
		301428 => x"FF",
		301549 => x"FF",
		301550 => x"FF",
		301551 => x"FF",
		301552 => x"FF",
		301553 => x"FF",
		302198 => x"FF",
		302199 => x"FF",
		302200 => x"FF",
		302201 => x"FF",
		302202 => x"FF",
		302323 => x"FF",
		302324 => x"FF",
		302325 => x"FF",
		302326 => x"FF",
		302327 => x"FF",
		302448 => x"FF",
		302449 => x"FF",
		302450 => x"FF",
		302451 => x"FF",
		302452 => x"FF",
		302573 => x"FF",
		302574 => x"FF",
		302575 => x"FF",
		302576 => x"FF",
		302577 => x"FF",
		303222 => x"FF",
		303223 => x"FF",
		303224 => x"FF",
		303225 => x"FF",
		303226 => x"FF",
		303347 => x"FF",
		303348 => x"FF",
		303349 => x"FF",
		303350 => x"FF",
		303351 => x"FF",
		303472 => x"FF",
		303473 => x"FF",
		303474 => x"FF",
		303475 => x"FF",
		303476 => x"FF",
		303597 => x"FF",
		303598 => x"FF",
		303599 => x"FF",
		303600 => x"FF",
		303601 => x"FF",
		304246 => x"FF",
		304247 => x"FF",
		304248 => x"FF",
		304249 => x"FF",
		304250 => x"FF",
		304371 => x"FF",
		304372 => x"FF",
		304373 => x"FF",
		304374 => x"FF",
		304375 => x"FF",
		304496 => x"FF",
		304497 => x"FF",
		304498 => x"FF",
		304499 => x"FF",
		304500 => x"FF",
		304621 => x"FF",
		304622 => x"FF",
		304623 => x"FF",
		304624 => x"FF",
		304625 => x"FF",
		305270 => x"FF",
		305271 => x"FF",
		305272 => x"FF",
		305273 => x"FF",
		305274 => x"FF",
		305275 => x"FF",
		305276 => x"FF",
		305277 => x"FF",
		305278 => x"FF",
		305279 => x"FF",
		305280 => x"FF",
		305281 => x"FF",
		305282 => x"FF",
		305283 => x"FF",
		305284 => x"FF",
		305285 => x"FF",
		305286 => x"FF",
		305287 => x"FF",
		305288 => x"FF",
		305289 => x"FF",
		305290 => x"FF",
		305291 => x"FF",
		305292 => x"FF",
		305293 => x"FF",
		305294 => x"FF",
		305295 => x"FF",
		305296 => x"FF",
		305297 => x"FF",
		305298 => x"FF",
		305299 => x"FF",
		305300 => x"FF",
		305301 => x"FF",
		305302 => x"FF",
		305303 => x"FF",
		305304 => x"FF",
		305305 => x"FF",
		305306 => x"FF",
		305307 => x"FF",
		305308 => x"FF",
		305309 => x"FF",
		305310 => x"FF",
		305311 => x"FF",
		305312 => x"FF",
		305313 => x"FF",
		305314 => x"FF",
		305315 => x"FF",
		305316 => x"FF",
		305317 => x"FF",
		305318 => x"FF",
		305319 => x"FF",
		305320 => x"FF",
		305321 => x"FF",
		305322 => x"FF",
		305323 => x"FF",
		305324 => x"FF",
		305325 => x"FF",
		305326 => x"FF",
		305327 => x"FF",
		305328 => x"FF",
		305329 => x"FF",
		305330 => x"FF",
		305331 => x"FF",
		305332 => x"FF",
		305333 => x"FF",
		305334 => x"FF",
		305335 => x"FF",
		305336 => x"FF",
		305337 => x"FF",
		305338 => x"FF",
		305339 => x"FF",
		305340 => x"FF",
		305341 => x"FF",
		305342 => x"FF",
		305343 => x"FF",
		305344 => x"FF",
		305345 => x"FF",
		305346 => x"FF",
		305347 => x"FF",
		305348 => x"FF",
		305349 => x"FF",
		305350 => x"FF",
		305351 => x"FF",
		305352 => x"FF",
		305353 => x"FF",
		305354 => x"FF",
		305355 => x"FF",
		305356 => x"FF",
		305357 => x"FF",
		305358 => x"FF",
		305359 => x"FF",
		305360 => x"FF",
		305361 => x"FF",
		305362 => x"FF",
		305363 => x"FF",
		305364 => x"FF",
		305365 => x"FF",
		305366 => x"FF",
		305367 => x"FF",
		305368 => x"FF",
		305369 => x"FF",
		305370 => x"FF",
		305371 => x"FF",
		305372 => x"FF",
		305373 => x"FF",
		305374 => x"FF",
		305375 => x"FF",
		305376 => x"FF",
		305377 => x"FF",
		305378 => x"FF",
		305379 => x"FF",
		305380 => x"FF",
		305381 => x"FF",
		305382 => x"FF",
		305383 => x"FF",
		305384 => x"FF",
		305385 => x"FF",
		305386 => x"FF",
		305387 => x"FF",
		305388 => x"FF",
		305389 => x"FF",
		305390 => x"FF",
		305391 => x"FF",
		305392 => x"FF",
		305393 => x"FF",
		305394 => x"FF",
		305395 => x"FF",
		305396 => x"FF",
		305397 => x"FF",
		305398 => x"FF",
		305399 => x"FF",
		305400 => x"FF",
		305401 => x"FF",
		305402 => x"FF",
		305403 => x"FF",
		305404 => x"FF",
		305405 => x"FF",
		305406 => x"FF",
		305407 => x"FF",
		305408 => x"FF",
		305409 => x"FF",
		305410 => x"FF",
		305411 => x"FF",
		305412 => x"FF",
		305413 => x"FF",
		305414 => x"FF",
		305415 => x"FF",
		305416 => x"FF",
		305417 => x"FF",
		305418 => x"FF",
		305419 => x"FF",
		305420 => x"FF",
		305421 => x"FF",
		305422 => x"FF",
		305423 => x"FF",
		305424 => x"FF",
		305425 => x"FF",
		305426 => x"FF",
		305427 => x"FF",
		305428 => x"FF",
		305429 => x"FF",
		305430 => x"FF",
		305431 => x"FF",
		305432 => x"FF",
		305433 => x"FF",
		305434 => x"FF",
		305435 => x"FF",
		305436 => x"FF",
		305437 => x"FF",
		305438 => x"FF",
		305439 => x"FF",
		305440 => x"FF",
		305441 => x"FF",
		305442 => x"FF",
		305443 => x"FF",
		305444 => x"FF",
		305445 => x"FF",
		305446 => x"FF",
		305447 => x"FF",
		305448 => x"FF",
		305449 => x"FF",
		305450 => x"FF",
		305451 => x"FF",
		305452 => x"FF",
		305453 => x"FF",
		305454 => x"FF",
		305455 => x"FF",
		305456 => x"FF",
		305457 => x"FF",
		305458 => x"FF",
		305459 => x"FF",
		305460 => x"FF",
		305461 => x"FF",
		305462 => x"FF",
		305463 => x"FF",
		305464 => x"FF",
		305465 => x"FF",
		305466 => x"FF",
		305467 => x"FF",
		305468 => x"FF",
		305469 => x"FF",
		305470 => x"FF",
		305471 => x"FF",
		305472 => x"FF",
		305473 => x"FF",
		305474 => x"FF",
		305475 => x"FF",
		305476 => x"FF",
		305477 => x"FF",
		305478 => x"FF",
		305479 => x"FF",
		305480 => x"FF",
		305481 => x"FF",
		305482 => x"FF",
		305483 => x"FF",
		305484 => x"FF",
		305485 => x"FF",
		305486 => x"FF",
		305487 => x"FF",
		305488 => x"FF",
		305489 => x"FF",
		305490 => x"FF",
		305491 => x"FF",
		305492 => x"FF",
		305493 => x"FF",
		305494 => x"FF",
		305495 => x"FF",
		305496 => x"FF",
		305497 => x"FF",
		305498 => x"FF",
		305499 => x"FF",
		305500 => x"FF",
		305501 => x"FF",
		305502 => x"FF",
		305503 => x"FF",
		305504 => x"FF",
		305505 => x"FF",
		305506 => x"FF",
		305507 => x"FF",
		305508 => x"FF",
		305509 => x"FF",
		305510 => x"FF",
		305511 => x"FF",
		305512 => x"FF",
		305513 => x"FF",
		305514 => x"FF",
		305515 => x"FF",
		305516 => x"FF",
		305517 => x"FF",
		305518 => x"FF",
		305519 => x"FF",
		305520 => x"FF",
		305521 => x"FF",
		305522 => x"FF",
		305523 => x"FF",
		305524 => x"FF",
		305525 => x"FF",
		305526 => x"FF",
		305527 => x"FF",
		305528 => x"FF",
		305529 => x"FF",
		305530 => x"FF",
		305531 => x"FF",
		305532 => x"FF",
		305533 => x"FF",
		305534 => x"FF",
		305535 => x"FF",
		305536 => x"FF",
		305537 => x"FF",
		305538 => x"FF",
		305539 => x"FF",
		305540 => x"FF",
		305541 => x"FF",
		305542 => x"FF",
		305543 => x"FF",
		305544 => x"FF",
		305545 => x"FF",
		305546 => x"FF",
		305547 => x"FF",
		305548 => x"FF",
		305549 => x"FF",
		305550 => x"FF",
		305551 => x"FF",
		305552 => x"FF",
		305553 => x"FF",
		305554 => x"FF",
		305555 => x"FF",
		305556 => x"FF",
		305557 => x"FF",
		305558 => x"FF",
		305559 => x"FF",
		305560 => x"FF",
		305561 => x"FF",
		305562 => x"FF",
		305563 => x"FF",
		305564 => x"FF",
		305565 => x"FF",
		305566 => x"FF",
		305567 => x"FF",
		305568 => x"FF",
		305569 => x"FF",
		305570 => x"FF",
		305571 => x"FF",
		305572 => x"FF",
		305573 => x"FF",
		305574 => x"FF",
		305575 => x"FF",
		305576 => x"FF",
		305577 => x"FF",
		305578 => x"FF",
		305579 => x"FF",
		305580 => x"FF",
		305581 => x"FF",
		305582 => x"FF",
		305583 => x"FF",
		305584 => x"FF",
		305585 => x"FF",
		305586 => x"FF",
		305587 => x"FF",
		305588 => x"FF",
		305589 => x"FF",
		305590 => x"FF",
		305591 => x"FF",
		305592 => x"FF",
		305593 => x"FF",
		305594 => x"FF",
		305595 => x"FF",
		305596 => x"FF",
		305597 => x"FF",
		305598 => x"FF",
		305599 => x"FF",
		305600 => x"FF",
		305601 => x"FF",
		305602 => x"FF",
		305603 => x"FF",
		305604 => x"FF",
		305605 => x"FF",
		305606 => x"FF",
		305607 => x"FF",
		305608 => x"FF",
		305609 => x"FF",
		305610 => x"FF",
		305611 => x"FF",
		305612 => x"FF",
		305613 => x"FF",
		305614 => x"FF",
		305615 => x"FF",
		305616 => x"FF",
		305617 => x"FF",
		305618 => x"FF",
		305619 => x"FF",
		305620 => x"FF",
		305621 => x"FF",
		305622 => x"FF",
		305623 => x"FF",
		305624 => x"FF",
		305625 => x"FF",
		305626 => x"FF",
		305627 => x"FF",
		305628 => x"FF",
		305629 => x"FF",
		305630 => x"FF",
		305631 => x"FF",
		305632 => x"FF",
		305633 => x"FF",
		305634 => x"FF",
		305635 => x"FF",
		305636 => x"FF",
		305637 => x"FF",
		305638 => x"FF",
		305639 => x"FF",
		305640 => x"FF",
		305641 => x"FF",
		305642 => x"FF",
		305643 => x"FF",
		305644 => x"FF",
		305645 => x"FF",
		305646 => x"FF",
		305647 => x"FF",
		305648 => x"FF",
		305649 => x"FF",
		306294 => x"FF",
		306295 => x"FF",
		306296 => x"FF",
		306297 => x"FF",
		306298 => x"FF",
		306299 => x"FF",
		306300 => x"FF",
		306301 => x"FF",
		306302 => x"FF",
		306303 => x"FF",
		306304 => x"FF",
		306305 => x"FF",
		306306 => x"FF",
		306307 => x"FF",
		306308 => x"FF",
		306309 => x"FF",
		306310 => x"FF",
		306311 => x"FF",
		306312 => x"FF",
		306313 => x"FF",
		306314 => x"FF",
		306315 => x"FF",
		306316 => x"FF",
		306317 => x"FF",
		306318 => x"FF",
		306319 => x"FF",
		306320 => x"FF",
		306321 => x"FF",
		306322 => x"FF",
		306323 => x"FF",
		306324 => x"FF",
		306325 => x"FF",
		306326 => x"FF",
		306327 => x"FF",
		306328 => x"FF",
		306329 => x"FF",
		306330 => x"FF",
		306331 => x"FF",
		306332 => x"FF",
		306333 => x"FF",
		306334 => x"FF",
		306335 => x"FF",
		306336 => x"FF",
		306337 => x"FF",
		306338 => x"FF",
		306339 => x"FF",
		306340 => x"FF",
		306341 => x"FF",
		306342 => x"FF",
		306343 => x"FF",
		306344 => x"FF",
		306345 => x"FF",
		306346 => x"FF",
		306347 => x"FF",
		306348 => x"FF",
		306349 => x"FF",
		306350 => x"FF",
		306351 => x"FF",
		306352 => x"FF",
		306353 => x"FF",
		306354 => x"FF",
		306355 => x"FF",
		306356 => x"FF",
		306357 => x"FF",
		306358 => x"FF",
		306359 => x"FF",
		306360 => x"FF",
		306361 => x"FF",
		306362 => x"FF",
		306363 => x"FF",
		306364 => x"FF",
		306365 => x"FF",
		306366 => x"FF",
		306367 => x"FF",
		306368 => x"FF",
		306369 => x"FF",
		306370 => x"FF",
		306371 => x"FF",
		306372 => x"FF",
		306373 => x"FF",
		306374 => x"FF",
		306375 => x"FF",
		306376 => x"FF",
		306377 => x"FF",
		306378 => x"FF",
		306379 => x"FF",
		306380 => x"FF",
		306381 => x"FF",
		306382 => x"FF",
		306383 => x"FF",
		306384 => x"FF",
		306385 => x"FF",
		306386 => x"FF",
		306387 => x"FF",
		306388 => x"FF",
		306389 => x"FF",
		306390 => x"FF",
		306391 => x"FF",
		306392 => x"FF",
		306393 => x"FF",
		306394 => x"FF",
		306395 => x"FF",
		306396 => x"FF",
		306397 => x"FF",
		306398 => x"FF",
		306399 => x"FF",
		306400 => x"FF",
		306401 => x"FF",
		306402 => x"FF",
		306403 => x"FF",
		306404 => x"FF",
		306405 => x"FF",
		306406 => x"FF",
		306407 => x"FF",
		306408 => x"FF",
		306409 => x"FF",
		306410 => x"FF",
		306411 => x"FF",
		306412 => x"FF",
		306413 => x"FF",
		306414 => x"FF",
		306415 => x"FF",
		306416 => x"FF",
		306417 => x"FF",
		306418 => x"FF",
		306419 => x"FF",
		306420 => x"FF",
		306421 => x"FF",
		306422 => x"FF",
		306423 => x"FF",
		306424 => x"FF",
		306425 => x"FF",
		306426 => x"FF",
		306427 => x"FF",
		306428 => x"FF",
		306429 => x"FF",
		306430 => x"FF",
		306431 => x"FF",
		306432 => x"FF",
		306433 => x"FF",
		306434 => x"FF",
		306435 => x"FF",
		306436 => x"FF",
		306437 => x"FF",
		306438 => x"FF",
		306439 => x"FF",
		306440 => x"FF",
		306441 => x"FF",
		306442 => x"FF",
		306443 => x"FF",
		306444 => x"FF",
		306445 => x"FF",
		306446 => x"FF",
		306447 => x"FF",
		306448 => x"FF",
		306449 => x"FF",
		306450 => x"FF",
		306451 => x"FF",
		306452 => x"FF",
		306453 => x"FF",
		306454 => x"FF",
		306455 => x"FF",
		306456 => x"FF",
		306457 => x"FF",
		306458 => x"FF",
		306459 => x"FF",
		306460 => x"FF",
		306461 => x"FF",
		306462 => x"FF",
		306463 => x"FF",
		306464 => x"FF",
		306465 => x"FF",
		306466 => x"FF",
		306467 => x"FF",
		306468 => x"FF",
		306469 => x"FF",
		306470 => x"FF",
		306471 => x"FF",
		306472 => x"FF",
		306473 => x"FF",
		306474 => x"FF",
		306475 => x"FF",
		306476 => x"FF",
		306477 => x"FF",
		306478 => x"FF",
		306479 => x"FF",
		306480 => x"FF",
		306481 => x"FF",
		306482 => x"FF",
		306483 => x"FF",
		306484 => x"FF",
		306485 => x"FF",
		306486 => x"FF",
		306487 => x"FF",
		306488 => x"FF",
		306489 => x"FF",
		306490 => x"FF",
		306491 => x"FF",
		306492 => x"FF",
		306493 => x"FF",
		306494 => x"FF",
		306495 => x"FF",
		306496 => x"FF",
		306497 => x"FF",
		306498 => x"FF",
		306499 => x"FF",
		306500 => x"FF",
		306501 => x"FF",
		306502 => x"FF",
		306503 => x"FF",
		306504 => x"FF",
		306505 => x"FF",
		306506 => x"FF",
		306507 => x"FF",
		306508 => x"FF",
		306509 => x"FF",
		306510 => x"FF",
		306511 => x"FF",
		306512 => x"FF",
		306513 => x"FF",
		306514 => x"FF",
		306515 => x"FF",
		306516 => x"FF",
		306517 => x"FF",
		306518 => x"FF",
		306519 => x"FF",
		306520 => x"FF",
		306521 => x"FF",
		306522 => x"FF",
		306523 => x"FF",
		306524 => x"FF",
		306525 => x"FF",
		306526 => x"FF",
		306527 => x"FF",
		306528 => x"FF",
		306529 => x"FF",
		306530 => x"FF",
		306531 => x"FF",
		306532 => x"FF",
		306533 => x"FF",
		306534 => x"FF",
		306535 => x"FF",
		306536 => x"FF",
		306537 => x"FF",
		306538 => x"FF",
		306539 => x"FF",
		306540 => x"FF",
		306541 => x"FF",
		306542 => x"FF",
		306543 => x"FF",
		306544 => x"FF",
		306545 => x"FF",
		306546 => x"FF",
		306547 => x"FF",
		306548 => x"FF",
		306549 => x"FF",
		306550 => x"FF",
		306551 => x"FF",
		306552 => x"FF",
		306553 => x"FF",
		306554 => x"FF",
		306555 => x"FF",
		306556 => x"FF",
		306557 => x"FF",
		306558 => x"FF",
		306559 => x"FF",
		306560 => x"FF",
		306561 => x"FF",
		306562 => x"FF",
		306563 => x"FF",
		306564 => x"FF",
		306565 => x"FF",
		306566 => x"FF",
		306567 => x"FF",
		306568 => x"FF",
		306569 => x"FF",
		306570 => x"FF",
		306571 => x"FF",
		306572 => x"FF",
		306573 => x"FF",
		306574 => x"FF",
		306575 => x"FF",
		306576 => x"FF",
		306577 => x"FF",
		306578 => x"FF",
		306579 => x"FF",
		306580 => x"FF",
		306581 => x"FF",
		306582 => x"FF",
		306583 => x"FF",
		306584 => x"FF",
		306585 => x"FF",
		306586 => x"FF",
		306587 => x"FF",
		306588 => x"FF",
		306589 => x"FF",
		306590 => x"FF",
		306591 => x"FF",
		306592 => x"FF",
		306593 => x"FF",
		306594 => x"FF",
		306595 => x"FF",
		306596 => x"FF",
		306597 => x"FF",
		306598 => x"FF",
		306599 => x"FF",
		306600 => x"FF",
		306601 => x"FF",
		306602 => x"FF",
		306603 => x"FF",
		306604 => x"FF",
		306605 => x"FF",
		306606 => x"FF",
		306607 => x"FF",
		306608 => x"FF",
		306609 => x"FF",
		306610 => x"FF",
		306611 => x"FF",
		306612 => x"FF",
		306613 => x"FF",
		306614 => x"FF",
		306615 => x"FF",
		306616 => x"FF",
		306617 => x"FF",
		306618 => x"FF",
		306619 => x"FF",
		306620 => x"FF",
		306621 => x"FF",
		306622 => x"FF",
		306623 => x"FF",
		306624 => x"FF",
		306625 => x"FF",
		306626 => x"FF",
		306627 => x"FF",
		306628 => x"FF",
		306629 => x"FF",
		306630 => x"FF",
		306631 => x"FF",
		306632 => x"FF",
		306633 => x"FF",
		306634 => x"FF",
		306635 => x"FF",
		306636 => x"FF",
		306637 => x"FF",
		306638 => x"FF",
		306639 => x"FF",
		306640 => x"FF",
		306641 => x"FF",
		306642 => x"FF",
		306643 => x"FF",
		306644 => x"FF",
		306645 => x"FF",
		306646 => x"FF",
		306647 => x"FF",
		306648 => x"FF",
		306649 => x"FF",
		306650 => x"FF",
		306651 => x"FF",
		306652 => x"FF",
		306653 => x"FF",
		306654 => x"FF",
		306655 => x"FF",
		306656 => x"FF",
		306657 => x"FF",
		306658 => x"FF",
		306659 => x"FF",
		306660 => x"FF",
		306661 => x"FF",
		306662 => x"FF",
		306663 => x"FF",
		306664 => x"FF",
		306665 => x"FF",
		306666 => x"FF",
		306667 => x"FF",
		306668 => x"FF",
		306669 => x"FF",
		306670 => x"FF",
		306671 => x"FF",
		306672 => x"FF",
		306673 => x"FF",
		307318 => x"FF",
		307319 => x"FF",
		307320 => x"FF",
		307321 => x"FF",
		307322 => x"FF",
		307323 => x"FF",
		307324 => x"FF",
		307325 => x"FF",
		307326 => x"FF",
		307327 => x"FF",
		307328 => x"FF",
		307329 => x"FF",
		307330 => x"FF",
		307331 => x"FF",
		307332 => x"FF",
		307333 => x"FF",
		307334 => x"FF",
		307335 => x"FF",
		307336 => x"FF",
		307337 => x"FF",
		307338 => x"FF",
		307339 => x"FF",
		307340 => x"FF",
		307341 => x"FF",
		307342 => x"FF",
		307343 => x"FF",
		307344 => x"FF",
		307345 => x"FF",
		307346 => x"FF",
		307347 => x"FF",
		307348 => x"FF",
		307349 => x"FF",
		307350 => x"FF",
		307351 => x"FF",
		307352 => x"FF",
		307353 => x"FF",
		307354 => x"FF",
		307355 => x"FF",
		307356 => x"FF",
		307357 => x"FF",
		307358 => x"FF",
		307359 => x"FF",
		307360 => x"FF",
		307361 => x"FF",
		307362 => x"FF",
		307363 => x"FF",
		307364 => x"FF",
		307365 => x"FF",
		307366 => x"FF",
		307367 => x"FF",
		307368 => x"FF",
		307369 => x"FF",
		307370 => x"FF",
		307371 => x"FF",
		307372 => x"FF",
		307373 => x"FF",
		307374 => x"FF",
		307375 => x"FF",
		307376 => x"FF",
		307377 => x"FF",
		307378 => x"FF",
		307379 => x"FF",
		307380 => x"FF",
		307381 => x"FF",
		307382 => x"FF",
		307383 => x"FF",
		307384 => x"FF",
		307385 => x"FF",
		307386 => x"FF",
		307387 => x"FF",
		307388 => x"FF",
		307389 => x"FF",
		307390 => x"FF",
		307391 => x"FF",
		307392 => x"FF",
		307393 => x"FF",
		307394 => x"FF",
		307395 => x"FF",
		307396 => x"FF",
		307397 => x"FF",
		307398 => x"FF",
		307399 => x"FF",
		307400 => x"FF",
		307401 => x"FF",
		307402 => x"FF",
		307403 => x"FF",
		307404 => x"FF",
		307405 => x"FF",
		307406 => x"FF",
		307407 => x"FF",
		307408 => x"FF",
		307409 => x"FF",
		307410 => x"FF",
		307411 => x"FF",
		307412 => x"FF",
		307413 => x"FF",
		307414 => x"FF",
		307415 => x"FF",
		307416 => x"FF",
		307417 => x"FF",
		307418 => x"FF",
		307419 => x"FF",
		307420 => x"FF",
		307421 => x"FF",
		307422 => x"FF",
		307423 => x"FF",
		307424 => x"FF",
		307425 => x"FF",
		307426 => x"FF",
		307427 => x"FF",
		307428 => x"FF",
		307429 => x"FF",
		307430 => x"FF",
		307431 => x"FF",
		307432 => x"FF",
		307433 => x"FF",
		307434 => x"FF",
		307435 => x"FF",
		307436 => x"FF",
		307437 => x"FF",
		307438 => x"FF",
		307439 => x"FF",
		307440 => x"FF",
		307441 => x"FF",
		307442 => x"FF",
		307443 => x"FF",
		307444 => x"FF",
		307445 => x"FF",
		307446 => x"FF",
		307447 => x"FF",
		307448 => x"FF",
		307449 => x"FF",
		307450 => x"FF",
		307451 => x"FF",
		307452 => x"FF",
		307453 => x"FF",
		307454 => x"FF",
		307455 => x"FF",
		307456 => x"FF",
		307457 => x"FF",
		307458 => x"FF",
		307459 => x"FF",
		307460 => x"FF",
		307461 => x"FF",
		307462 => x"FF",
		307463 => x"FF",
		307464 => x"FF",
		307465 => x"FF",
		307466 => x"FF",
		307467 => x"FF",
		307468 => x"FF",
		307469 => x"FF",
		307470 => x"FF",
		307471 => x"FF",
		307472 => x"FF",
		307473 => x"FF",
		307474 => x"FF",
		307475 => x"FF",
		307476 => x"FF",
		307477 => x"FF",
		307478 => x"FF",
		307479 => x"FF",
		307480 => x"FF",
		307481 => x"FF",
		307482 => x"FF",
		307483 => x"FF",
		307484 => x"FF",
		307485 => x"FF",
		307486 => x"FF",
		307487 => x"FF",
		307488 => x"FF",
		307489 => x"FF",
		307490 => x"FF",
		307491 => x"FF",
		307492 => x"FF",
		307493 => x"FF",
		307494 => x"FF",
		307495 => x"FF",
		307496 => x"FF",
		307497 => x"FF",
		307498 => x"FF",
		307499 => x"FF",
		307500 => x"FF",
		307501 => x"FF",
		307502 => x"FF",
		307503 => x"FF",
		307504 => x"FF",
		307505 => x"FF",
		307506 => x"FF",
		307507 => x"FF",
		307508 => x"FF",
		307509 => x"FF",
		307510 => x"FF",
		307511 => x"FF",
		307512 => x"FF",
		307513 => x"FF",
		307514 => x"FF",
		307515 => x"FF",
		307516 => x"FF",
		307517 => x"FF",
		307518 => x"FF",
		307519 => x"FF",
		307520 => x"FF",
		307521 => x"FF",
		307522 => x"FF",
		307523 => x"FF",
		307524 => x"FF",
		307525 => x"FF",
		307526 => x"FF",
		307527 => x"FF",
		307528 => x"FF",
		307529 => x"FF",
		307530 => x"FF",
		307531 => x"FF",
		307532 => x"FF",
		307533 => x"FF",
		307534 => x"FF",
		307535 => x"FF",
		307536 => x"FF",
		307537 => x"FF",
		307538 => x"FF",
		307539 => x"FF",
		307540 => x"FF",
		307541 => x"FF",
		307542 => x"FF",
		307543 => x"FF",
		307544 => x"FF",
		307545 => x"FF",
		307546 => x"FF",
		307547 => x"FF",
		307548 => x"FF",
		307549 => x"FF",
		307550 => x"FF",
		307551 => x"FF",
		307552 => x"FF",
		307553 => x"FF",
		307554 => x"FF",
		307555 => x"FF",
		307556 => x"FF",
		307557 => x"FF",
		307558 => x"FF",
		307559 => x"FF",
		307560 => x"FF",
		307561 => x"FF",
		307562 => x"FF",
		307563 => x"FF",
		307564 => x"FF",
		307565 => x"FF",
		307566 => x"FF",
		307567 => x"FF",
		307568 => x"FF",
		307569 => x"FF",
		307570 => x"FF",
		307571 => x"FF",
		307572 => x"FF",
		307573 => x"FF",
		307574 => x"FF",
		307575 => x"FF",
		307576 => x"FF",
		307577 => x"FF",
		307578 => x"FF",
		307579 => x"FF",
		307580 => x"FF",
		307581 => x"FF",
		307582 => x"FF",
		307583 => x"FF",
		307584 => x"FF",
		307585 => x"FF",
		307586 => x"FF",
		307587 => x"FF",
		307588 => x"FF",
		307589 => x"FF",
		307590 => x"FF",
		307591 => x"FF",
		307592 => x"FF",
		307593 => x"FF",
		307594 => x"FF",
		307595 => x"FF",
		307596 => x"FF",
		307597 => x"FF",
		307598 => x"FF",
		307599 => x"FF",
		307600 => x"FF",
		307601 => x"FF",
		307602 => x"FF",
		307603 => x"FF",
		307604 => x"FF",
		307605 => x"FF",
		307606 => x"FF",
		307607 => x"FF",
		307608 => x"FF",
		307609 => x"FF",
		307610 => x"FF",
		307611 => x"FF",
		307612 => x"FF",
		307613 => x"FF",
		307614 => x"FF",
		307615 => x"FF",
		307616 => x"FF",
		307617 => x"FF",
		307618 => x"FF",
		307619 => x"FF",
		307620 => x"FF",
		307621 => x"FF",
		307622 => x"FF",
		307623 => x"FF",
		307624 => x"FF",
		307625 => x"FF",
		307626 => x"FF",
		307627 => x"FF",
		307628 => x"FF",
		307629 => x"FF",
		307630 => x"FF",
		307631 => x"FF",
		307632 => x"FF",
		307633 => x"FF",
		307634 => x"FF",
		307635 => x"FF",
		307636 => x"FF",
		307637 => x"FF",
		307638 => x"FF",
		307639 => x"FF",
		307640 => x"FF",
		307641 => x"FF",
		307642 => x"FF",
		307643 => x"FF",
		307644 => x"FF",
		307645 => x"FF",
		307646 => x"FF",
		307647 => x"FF",
		307648 => x"FF",
		307649 => x"FF",
		307650 => x"FF",
		307651 => x"FF",
		307652 => x"FF",
		307653 => x"FF",
		307654 => x"FF",
		307655 => x"FF",
		307656 => x"FF",
		307657 => x"FF",
		307658 => x"FF",
		307659 => x"FF",
		307660 => x"FF",
		307661 => x"FF",
		307662 => x"FF",
		307663 => x"FF",
		307664 => x"FF",
		307665 => x"FF",
		307666 => x"FF",
		307667 => x"FF",
		307668 => x"FF",
		307669 => x"FF",
		307670 => x"FF",
		307671 => x"FF",
		307672 => x"FF",
		307673 => x"FF",
		307674 => x"FF",
		307675 => x"FF",
		307676 => x"FF",
		307677 => x"FF",
		307678 => x"FF",
		307679 => x"FF",
		307680 => x"FF",
		307681 => x"FF",
		307682 => x"FF",
		307683 => x"FF",
		307684 => x"FF",
		307685 => x"FF",
		307686 => x"FF",
		307687 => x"FF",
		307688 => x"FF",
		307689 => x"FF",
		307690 => x"FF",
		307691 => x"FF",
		307692 => x"FF",
		307693 => x"FF",
		307694 => x"FF",
		307695 => x"FF",
		307696 => x"FF",
		307697 => x"FF",
		308342 => x"FF",
		308343 => x"FF",
		308344 => x"FF",
		308345 => x"FF",
		308346 => x"FF",
		308347 => x"FF",
		308348 => x"FF",
		308349 => x"FF",
		308350 => x"FF",
		308351 => x"FF",
		308352 => x"FF",
		308353 => x"FF",
		308354 => x"FF",
		308355 => x"FF",
		308356 => x"FF",
		308357 => x"FF",
		308358 => x"FF",
		308359 => x"FF",
		308360 => x"FF",
		308361 => x"FF",
		308362 => x"FF",
		308363 => x"FF",
		308364 => x"FF",
		308365 => x"FF",
		308366 => x"FF",
		308367 => x"FF",
		308368 => x"FF",
		308369 => x"FF",
		308370 => x"FF",
		308371 => x"FF",
		308372 => x"FF",
		308373 => x"FF",
		308374 => x"FF",
		308375 => x"FF",
		308376 => x"FF",
		308377 => x"FF",
		308378 => x"FF",
		308379 => x"FF",
		308380 => x"FF",
		308381 => x"FF",
		308382 => x"FF",
		308383 => x"FF",
		308384 => x"FF",
		308385 => x"FF",
		308386 => x"FF",
		308387 => x"FF",
		308388 => x"FF",
		308389 => x"FF",
		308390 => x"FF",
		308391 => x"FF",
		308392 => x"FF",
		308393 => x"FF",
		308394 => x"FF",
		308395 => x"FF",
		308396 => x"FF",
		308397 => x"FF",
		308398 => x"FF",
		308399 => x"FF",
		308400 => x"FF",
		308401 => x"FF",
		308402 => x"FF",
		308403 => x"FF",
		308404 => x"FF",
		308405 => x"FF",
		308406 => x"FF",
		308407 => x"FF",
		308408 => x"FF",
		308409 => x"FF",
		308410 => x"FF",
		308411 => x"FF",
		308412 => x"FF",
		308413 => x"FF",
		308414 => x"FF",
		308415 => x"FF",
		308416 => x"FF",
		308417 => x"FF",
		308418 => x"FF",
		308419 => x"FF",
		308420 => x"FF",
		308421 => x"FF",
		308422 => x"FF",
		308423 => x"FF",
		308424 => x"FF",
		308425 => x"FF",
		308426 => x"FF",
		308427 => x"FF",
		308428 => x"FF",
		308429 => x"FF",
		308430 => x"FF",
		308431 => x"FF",
		308432 => x"FF",
		308433 => x"FF",
		308434 => x"FF",
		308435 => x"FF",
		308436 => x"FF",
		308437 => x"FF",
		308438 => x"FF",
		308439 => x"FF",
		308440 => x"FF",
		308441 => x"FF",
		308442 => x"FF",
		308443 => x"FF",
		308444 => x"FF",
		308445 => x"FF",
		308446 => x"FF",
		308447 => x"FF",
		308448 => x"FF",
		308449 => x"FF",
		308450 => x"FF",
		308451 => x"FF",
		308452 => x"FF",
		308453 => x"FF",
		308454 => x"FF",
		308455 => x"FF",
		308456 => x"FF",
		308457 => x"FF",
		308458 => x"FF",
		308459 => x"FF",
		308460 => x"FF",
		308461 => x"FF",
		308462 => x"FF",
		308463 => x"FF",
		308464 => x"FF",
		308465 => x"FF",
		308466 => x"FF",
		308467 => x"FF",
		308468 => x"FF",
		308469 => x"FF",
		308470 => x"FF",
		308471 => x"FF",
		308472 => x"FF",
		308473 => x"FF",
		308474 => x"FF",
		308475 => x"FF",
		308476 => x"FF",
		308477 => x"FF",
		308478 => x"FF",
		308479 => x"FF",
		308480 => x"FF",
		308481 => x"FF",
		308482 => x"FF",
		308483 => x"FF",
		308484 => x"FF",
		308485 => x"FF",
		308486 => x"FF",
		308487 => x"FF",
		308488 => x"FF",
		308489 => x"FF",
		308490 => x"FF",
		308491 => x"FF",
		308492 => x"FF",
		308493 => x"FF",
		308494 => x"FF",
		308495 => x"FF",
		308496 => x"FF",
		308497 => x"FF",
		308498 => x"FF",
		308499 => x"FF",
		308500 => x"FF",
		308501 => x"FF",
		308502 => x"FF",
		308503 => x"FF",
		308504 => x"FF",
		308505 => x"FF",
		308506 => x"FF",
		308507 => x"FF",
		308508 => x"FF",
		308509 => x"FF",
		308510 => x"FF",
		308511 => x"FF",
		308512 => x"FF",
		308513 => x"FF",
		308514 => x"FF",
		308515 => x"FF",
		308516 => x"FF",
		308517 => x"FF",
		308518 => x"FF",
		308519 => x"FF",
		308520 => x"FF",
		308521 => x"FF",
		308522 => x"FF",
		308523 => x"FF",
		308524 => x"FF",
		308525 => x"FF",
		308526 => x"FF",
		308527 => x"FF",
		308528 => x"FF",
		308529 => x"FF",
		308530 => x"FF",
		308531 => x"FF",
		308532 => x"FF",
		308533 => x"FF",
		308534 => x"FF",
		308535 => x"FF",
		308536 => x"FF",
		308537 => x"FF",
		308538 => x"FF",
		308539 => x"FF",
		308540 => x"FF",
		308541 => x"FF",
		308542 => x"FF",
		308543 => x"FF",
		308544 => x"FF",
		308545 => x"FF",
		308546 => x"FF",
		308547 => x"FF",
		308548 => x"FF",
		308549 => x"FF",
		308550 => x"FF",
		308551 => x"FF",
		308552 => x"FF",
		308553 => x"FF",
		308554 => x"FF",
		308555 => x"FF",
		308556 => x"FF",
		308557 => x"FF",
		308558 => x"FF",
		308559 => x"FF",
		308560 => x"FF",
		308561 => x"FF",
		308562 => x"FF",
		308563 => x"FF",
		308564 => x"FF",
		308565 => x"FF",
		308566 => x"FF",
		308567 => x"FF",
		308568 => x"FF",
		308569 => x"FF",
		308570 => x"FF",
		308571 => x"FF",
		308572 => x"FF",
		308573 => x"FF",
		308574 => x"FF",
		308575 => x"FF",
		308576 => x"FF",
		308577 => x"FF",
		308578 => x"FF",
		308579 => x"FF",
		308580 => x"FF",
		308581 => x"FF",
		308582 => x"FF",
		308583 => x"FF",
		308584 => x"FF",
		308585 => x"FF",
		308586 => x"FF",
		308587 => x"FF",
		308588 => x"FF",
		308589 => x"FF",
		308590 => x"FF",
		308591 => x"FF",
		308592 => x"FF",
		308593 => x"FF",
		308594 => x"FF",
		308595 => x"FF",
		308596 => x"FF",
		308597 => x"FF",
		308598 => x"FF",
		308599 => x"FF",
		308600 => x"FF",
		308601 => x"FF",
		308602 => x"FF",
		308603 => x"FF",
		308604 => x"FF",
		308605 => x"FF",
		308606 => x"FF",
		308607 => x"FF",
		308608 => x"FF",
		308609 => x"FF",
		308610 => x"FF",
		308611 => x"FF",
		308612 => x"FF",
		308613 => x"FF",
		308614 => x"FF",
		308615 => x"FF",
		308616 => x"FF",
		308617 => x"FF",
		308618 => x"FF",
		308619 => x"FF",
		308620 => x"FF",
		308621 => x"FF",
		308622 => x"FF",
		308623 => x"FF",
		308624 => x"FF",
		308625 => x"FF",
		308626 => x"FF",
		308627 => x"FF",
		308628 => x"FF",
		308629 => x"FF",
		308630 => x"FF",
		308631 => x"FF",
		308632 => x"FF",
		308633 => x"FF",
		308634 => x"FF",
		308635 => x"FF",
		308636 => x"FF",
		308637 => x"FF",
		308638 => x"FF",
		308639 => x"FF",
		308640 => x"FF",
		308641 => x"FF",
		308642 => x"FF",
		308643 => x"FF",
		308644 => x"FF",
		308645 => x"FF",
		308646 => x"FF",
		308647 => x"FF",
		308648 => x"FF",
		308649 => x"FF",
		308650 => x"FF",
		308651 => x"FF",
		308652 => x"FF",
		308653 => x"FF",
		308654 => x"FF",
		308655 => x"FF",
		308656 => x"FF",
		308657 => x"FF",
		308658 => x"FF",
		308659 => x"FF",
		308660 => x"FF",
		308661 => x"FF",
		308662 => x"FF",
		308663 => x"FF",
		308664 => x"FF",
		308665 => x"FF",
		308666 => x"FF",
		308667 => x"FF",
		308668 => x"FF",
		308669 => x"FF",
		308670 => x"FF",
		308671 => x"FF",
		308672 => x"FF",
		308673 => x"FF",
		308674 => x"FF",
		308675 => x"FF",
		308676 => x"FF",
		308677 => x"FF",
		308678 => x"FF",
		308679 => x"FF",
		308680 => x"FF",
		308681 => x"FF",
		308682 => x"FF",
		308683 => x"FF",
		308684 => x"FF",
		308685 => x"FF",
		308686 => x"FF",
		308687 => x"FF",
		308688 => x"FF",
		308689 => x"FF",
		308690 => x"FF",
		308691 => x"FF",
		308692 => x"FF",
		308693 => x"FF",
		308694 => x"FF",
		308695 => x"FF",
		308696 => x"FF",
		308697 => x"FF",
		308698 => x"FF",
		308699 => x"FF",
		308700 => x"FF",
		308701 => x"FF",
		308702 => x"FF",
		308703 => x"FF",
		308704 => x"FF",
		308705 => x"FF",
		308706 => x"FF",
		308707 => x"FF",
		308708 => x"FF",
		308709 => x"FF",
		308710 => x"FF",
		308711 => x"FF",
		308712 => x"FF",
		308713 => x"FF",
		308714 => x"FF",
		308715 => x"FF",
		308716 => x"FF",
		308717 => x"FF",
		308718 => x"FF",
		308719 => x"FF",
		308720 => x"FF",
		308721 => x"FF",
		309366 => x"FF",
		309367 => x"FF",
		309368 => x"FF",
		309369 => x"FF",
		309370 => x"FF",
		309371 => x"FF",
		309372 => x"FF",
		309373 => x"FF",
		309374 => x"FF",
		309375 => x"FF",
		309376 => x"FF",
		309377 => x"FF",
		309378 => x"FF",
		309379 => x"FF",
		309380 => x"FF",
		309381 => x"FF",
		309382 => x"FF",
		309383 => x"FF",
		309384 => x"FF",
		309385 => x"FF",
		309386 => x"FF",
		309387 => x"FF",
		309388 => x"FF",
		309389 => x"FF",
		309390 => x"FF",
		309391 => x"FF",
		309392 => x"FF",
		309393 => x"FF",
		309394 => x"FF",
		309395 => x"FF",
		309396 => x"FF",
		309397 => x"FF",
		309398 => x"FF",
		309399 => x"FF",
		309400 => x"FF",
		309401 => x"FF",
		309402 => x"FF",
		309403 => x"FF",
		309404 => x"FF",
		309405 => x"FF",
		309406 => x"FF",
		309407 => x"FF",
		309408 => x"FF",
		309409 => x"FF",
		309410 => x"FF",
		309411 => x"FF",
		309412 => x"FF",
		309413 => x"FF",
		309414 => x"FF",
		309415 => x"FF",
		309416 => x"FF",
		309417 => x"FF",
		309418 => x"FF",
		309419 => x"FF",
		309420 => x"FF",
		309421 => x"FF",
		309422 => x"FF",
		309423 => x"FF",
		309424 => x"FF",
		309425 => x"FF",
		309426 => x"FF",
		309427 => x"FF",
		309428 => x"FF",
		309429 => x"FF",
		309430 => x"FF",
		309431 => x"FF",
		309432 => x"FF",
		309433 => x"FF",
		309434 => x"FF",
		309435 => x"FF",
		309436 => x"FF",
		309437 => x"FF",
		309438 => x"FF",
		309439 => x"FF",
		309440 => x"FF",
		309441 => x"FF",
		309442 => x"FF",
		309443 => x"FF",
		309444 => x"FF",
		309445 => x"FF",
		309446 => x"FF",
		309447 => x"FF",
		309448 => x"FF",
		309449 => x"FF",
		309450 => x"FF",
		309451 => x"FF",
		309452 => x"FF",
		309453 => x"FF",
		309454 => x"FF",
		309455 => x"FF",
		309456 => x"FF",
		309457 => x"FF",
		309458 => x"FF",
		309459 => x"FF",
		309460 => x"FF",
		309461 => x"FF",
		309462 => x"FF",
		309463 => x"FF",
		309464 => x"FF",
		309465 => x"FF",
		309466 => x"FF",
		309467 => x"FF",
		309468 => x"FF",
		309469 => x"FF",
		309470 => x"FF",
		309471 => x"FF",
		309472 => x"FF",
		309473 => x"FF",
		309474 => x"FF",
		309475 => x"FF",
		309476 => x"FF",
		309477 => x"FF",
		309478 => x"FF",
		309479 => x"FF",
		309480 => x"FF",
		309481 => x"FF",
		309482 => x"FF",
		309483 => x"FF",
		309484 => x"FF",
		309485 => x"FF",
		309486 => x"FF",
		309487 => x"FF",
		309488 => x"FF",
		309489 => x"FF",
		309490 => x"FF",
		309491 => x"FF",
		309492 => x"FF",
		309493 => x"FF",
		309494 => x"FF",
		309495 => x"FF",
		309496 => x"FF",
		309497 => x"FF",
		309498 => x"FF",
		309499 => x"FF",
		309500 => x"FF",
		309501 => x"FF",
		309502 => x"FF",
		309503 => x"FF",
		309504 => x"FF",
		309505 => x"FF",
		309506 => x"FF",
		309507 => x"FF",
		309508 => x"FF",
		309509 => x"FF",
		309510 => x"FF",
		309511 => x"FF",
		309512 => x"FF",
		309513 => x"FF",
		309514 => x"FF",
		309515 => x"FF",
		309516 => x"FF",
		309517 => x"FF",
		309518 => x"FF",
		309519 => x"FF",
		309520 => x"FF",
		309521 => x"FF",
		309522 => x"FF",
		309523 => x"FF",
		309524 => x"FF",
		309525 => x"FF",
		309526 => x"FF",
		309527 => x"FF",
		309528 => x"FF",
		309529 => x"FF",
		309530 => x"FF",
		309531 => x"FF",
		309532 => x"FF",
		309533 => x"FF",
		309534 => x"FF",
		309535 => x"FF",
		309536 => x"FF",
		309537 => x"FF",
		309538 => x"FF",
		309539 => x"FF",
		309540 => x"FF",
		309541 => x"FF",
		309542 => x"FF",
		309543 => x"FF",
		309544 => x"FF",
		309545 => x"FF",
		309546 => x"FF",
		309547 => x"FF",
		309548 => x"FF",
		309549 => x"FF",
		309550 => x"FF",
		309551 => x"FF",
		309552 => x"FF",
		309553 => x"FF",
		309554 => x"FF",
		309555 => x"FF",
		309556 => x"FF",
		309557 => x"FF",
		309558 => x"FF",
		309559 => x"FF",
		309560 => x"FF",
		309561 => x"FF",
		309562 => x"FF",
		309563 => x"FF",
		309564 => x"FF",
		309565 => x"FF",
		309566 => x"FF",
		309567 => x"FF",
		309568 => x"FF",
		309569 => x"FF",
		309570 => x"FF",
		309571 => x"FF",
		309572 => x"FF",
		309573 => x"FF",
		309574 => x"FF",
		309575 => x"FF",
		309576 => x"FF",
		309577 => x"FF",
		309578 => x"FF",
		309579 => x"FF",
		309580 => x"FF",
		309581 => x"FF",
		309582 => x"FF",
		309583 => x"FF",
		309584 => x"FF",
		309585 => x"FF",
		309586 => x"FF",
		309587 => x"FF",
		309588 => x"FF",
		309589 => x"FF",
		309590 => x"FF",
		309591 => x"FF",
		309592 => x"FF",
		309593 => x"FF",
		309594 => x"FF",
		309595 => x"FF",
		309596 => x"FF",
		309597 => x"FF",
		309598 => x"FF",
		309599 => x"FF",
		309600 => x"FF",
		309601 => x"FF",
		309602 => x"FF",
		309603 => x"FF",
		309604 => x"FF",
		309605 => x"FF",
		309606 => x"FF",
		309607 => x"FF",
		309608 => x"FF",
		309609 => x"FF",
		309610 => x"FF",
		309611 => x"FF",
		309612 => x"FF",
		309613 => x"FF",
		309614 => x"FF",
		309615 => x"FF",
		309616 => x"FF",
		309617 => x"FF",
		309618 => x"FF",
		309619 => x"FF",
		309620 => x"FF",
		309621 => x"FF",
		309622 => x"FF",
		309623 => x"FF",
		309624 => x"FF",
		309625 => x"FF",
		309626 => x"FF",
		309627 => x"FF",
		309628 => x"FF",
		309629 => x"FF",
		309630 => x"FF",
		309631 => x"FF",
		309632 => x"FF",
		309633 => x"FF",
		309634 => x"FF",
		309635 => x"FF",
		309636 => x"FF",
		309637 => x"FF",
		309638 => x"FF",
		309639 => x"FF",
		309640 => x"FF",
		309641 => x"FF",
		309642 => x"FF",
		309643 => x"FF",
		309644 => x"FF",
		309645 => x"FF",
		309646 => x"FF",
		309647 => x"FF",
		309648 => x"FF",
		309649 => x"FF",
		309650 => x"FF",
		309651 => x"FF",
		309652 => x"FF",
		309653 => x"FF",
		309654 => x"FF",
		309655 => x"FF",
		309656 => x"FF",
		309657 => x"FF",
		309658 => x"FF",
		309659 => x"FF",
		309660 => x"FF",
		309661 => x"FF",
		309662 => x"FF",
		309663 => x"FF",
		309664 => x"FF",
		309665 => x"FF",
		309666 => x"FF",
		309667 => x"FF",
		309668 => x"FF",
		309669 => x"FF",
		309670 => x"FF",
		309671 => x"FF",
		309672 => x"FF",
		309673 => x"FF",
		309674 => x"FF",
		309675 => x"FF",
		309676 => x"FF",
		309677 => x"FF",
		309678 => x"FF",
		309679 => x"FF",
		309680 => x"FF",
		309681 => x"FF",
		309682 => x"FF",
		309683 => x"FF",
		309684 => x"FF",
		309685 => x"FF",
		309686 => x"FF",
		309687 => x"FF",
		309688 => x"FF",
		309689 => x"FF",
		309690 => x"FF",
		309691 => x"FF",
		309692 => x"FF",
		309693 => x"FF",
		309694 => x"FF",
		309695 => x"FF",
		309696 => x"FF",
		309697 => x"FF",
		309698 => x"FF",
		309699 => x"FF",
		309700 => x"FF",
		309701 => x"FF",
		309702 => x"FF",
		309703 => x"FF",
		309704 => x"FF",
		309705 => x"FF",
		309706 => x"FF",
		309707 => x"FF",
		309708 => x"FF",
		309709 => x"FF",
		309710 => x"FF",
		309711 => x"FF",
		309712 => x"FF",
		309713 => x"FF",
		309714 => x"FF",
		309715 => x"FF",
		309716 => x"FF",
		309717 => x"FF",
		309718 => x"FF",
		309719 => x"FF",
		309720 => x"FF",
		309721 => x"FF",
		309722 => x"FF",
		309723 => x"FF",
		309724 => x"FF",
		309725 => x"FF",
		309726 => x"FF",
		309727 => x"FF",
		309728 => x"FF",
		309729 => x"FF",
		309730 => x"FF",
		309731 => x"FF",
		309732 => x"FF",
		309733 => x"FF",
		309734 => x"FF",
		309735 => x"FF",
		309736 => x"FF",
		309737 => x"FF",
		309738 => x"FF",
		309739 => x"FF",
		309740 => x"FF",
		309741 => x"FF",
		309742 => x"FF",
		309743 => x"FF",
		309744 => x"FF",
		309745 => x"FF",
		310390 => x"FF",
		310391 => x"FF",
		310392 => x"FF",
		310393 => x"FF",
		310394 => x"FF",
		310515 => x"FF",
		310516 => x"FF",
		310517 => x"FF",
		310518 => x"FF",
		310519 => x"FF",
		310640 => x"FF",
		310641 => x"FF",
		310642 => x"FF",
		310643 => x"FF",
		310644 => x"FF",
		310765 => x"FF",
		310766 => x"FF",
		310767 => x"FF",
		310768 => x"FF",
		310769 => x"FF",
		311414 => x"FF",
		311415 => x"FF",
		311416 => x"FF",
		311417 => x"FF",
		311418 => x"FF",
		311539 => x"FF",
		311540 => x"FF",
		311541 => x"FF",
		311542 => x"FF",
		311543 => x"FF",
		311664 => x"FF",
		311665 => x"FF",
		311666 => x"FF",
		311667 => x"FF",
		311668 => x"FF",
		311789 => x"FF",
		311790 => x"FF",
		311791 => x"FF",
		311792 => x"FF",
		311793 => x"FF",
		312438 => x"FF",
		312439 => x"FF",
		312440 => x"FF",
		312441 => x"FF",
		312442 => x"FF",
		312563 => x"FF",
		312564 => x"FF",
		312565 => x"FF",
		312566 => x"FF",
		312567 => x"FF",
		312688 => x"FF",
		312689 => x"FF",
		312690 => x"FF",
		312691 => x"FF",
		312692 => x"FF",
		312813 => x"FF",
		312814 => x"FF",
		312815 => x"FF",
		312816 => x"FF",
		312817 => x"FF",
		313462 => x"FF",
		313463 => x"FF",
		313464 => x"FF",
		313465 => x"FF",
		313466 => x"FF",
		313587 => x"FF",
		313588 => x"FF",
		313589 => x"FF",
		313590 => x"FF",
		313591 => x"FF",
		313712 => x"FF",
		313713 => x"FF",
		313714 => x"FF",
		313715 => x"FF",
		313716 => x"FF",
		313837 => x"FF",
		313838 => x"FF",
		313839 => x"FF",
		313840 => x"FF",
		313841 => x"FF",
		314486 => x"FF",
		314487 => x"FF",
		314488 => x"FF",
		314489 => x"FF",
		314490 => x"FF",
		314611 => x"FF",
		314612 => x"FF",
		314613 => x"FF",
		314614 => x"FF",
		314615 => x"FF",
		314736 => x"FF",
		314737 => x"FF",
		314738 => x"FF",
		314739 => x"FF",
		314740 => x"FF",
		314861 => x"FF",
		314862 => x"FF",
		314863 => x"FF",
		314864 => x"FF",
		314865 => x"FF",
		315510 => x"FF",
		315511 => x"FF",
		315512 => x"FF",
		315513 => x"FF",
		315514 => x"FF",
		315635 => x"FF",
		315636 => x"FF",
		315637 => x"FF",
		315638 => x"FF",
		315639 => x"FF",
		315760 => x"FF",
		315761 => x"FF",
		315762 => x"FF",
		315763 => x"FF",
		315764 => x"FF",
		315885 => x"FF",
		315886 => x"FF",
		315887 => x"FF",
		315888 => x"FF",
		315889 => x"FF",
		316534 => x"FF",
		316535 => x"FF",
		316536 => x"FF",
		316537 => x"FF",
		316538 => x"FF",
		316659 => x"FF",
		316660 => x"FF",
		316661 => x"FF",
		316662 => x"FF",
		316663 => x"FF",
		316784 => x"FF",
		316785 => x"FF",
		316786 => x"FF",
		316787 => x"FF",
		316788 => x"FF",
		316909 => x"FF",
		316910 => x"FF",
		316911 => x"FF",
		316912 => x"FF",
		316913 => x"FF",
		317558 => x"FF",
		317559 => x"FF",
		317560 => x"FF",
		317561 => x"FF",
		317562 => x"FF",
		317683 => x"FF",
		317684 => x"FF",
		317685 => x"FF",
		317686 => x"FF",
		317687 => x"FF",
		317808 => x"FF",
		317809 => x"FF",
		317810 => x"FF",
		317811 => x"FF",
		317812 => x"FF",
		317933 => x"FF",
		317934 => x"FF",
		317935 => x"FF",
		317936 => x"FF",
		317937 => x"FF",
		318582 => x"FF",
		318583 => x"FF",
		318584 => x"FF",
		318585 => x"FF",
		318586 => x"FF",
		318707 => x"FF",
		318708 => x"FF",
		318709 => x"FF",
		318710 => x"FF",
		318711 => x"FF",
		318832 => x"FF",
		318833 => x"FF",
		318834 => x"FF",
		318835 => x"FF",
		318836 => x"FF",
		318957 => x"FF",
		318958 => x"FF",
		318959 => x"FF",
		318960 => x"FF",
		318961 => x"FF",
		319606 => x"FF",
		319607 => x"FF",
		319608 => x"FF",
		319609 => x"FF",
		319610 => x"FF",
		319731 => x"FF",
		319732 => x"FF",
		319733 => x"FF",
		319734 => x"FF",
		319735 => x"FF",
		319856 => x"FF",
		319857 => x"FF",
		319858 => x"FF",
		319859 => x"FF",
		319860 => x"FF",
		319981 => x"FF",
		319982 => x"FF",
		319983 => x"FF",
		319984 => x"FF",
		319985 => x"FF",
		320630 => x"FF",
		320631 => x"FF",
		320632 => x"FF",
		320633 => x"FF",
		320634 => x"FF",
		320755 => x"FF",
		320756 => x"FF",
		320757 => x"FF",
		320758 => x"FF",
		320759 => x"FF",
		320880 => x"FF",
		320881 => x"FF",
		320882 => x"FF",
		320883 => x"FF",
		320884 => x"FF",
		321005 => x"FF",
		321006 => x"FF",
		321007 => x"FF",
		321008 => x"FF",
		321009 => x"FF",
		321654 => x"FF",
		321655 => x"FF",
		321656 => x"FF",
		321657 => x"FF",
		321658 => x"FF",
		321779 => x"FF",
		321780 => x"FF",
		321781 => x"FF",
		321782 => x"FF",
		321783 => x"FF",
		321904 => x"FF",
		321905 => x"FF",
		321906 => x"FF",
		321907 => x"FF",
		321908 => x"FF",
		322029 => x"FF",
		322030 => x"FF",
		322031 => x"FF",
		322032 => x"FF",
		322033 => x"FF",
		322678 => x"FF",
		322679 => x"FF",
		322680 => x"FF",
		322681 => x"FF",
		322682 => x"FF",
		322803 => x"FF",
		322804 => x"FF",
		322805 => x"FF",
		322806 => x"FF",
		322807 => x"FF",
		322928 => x"FF",
		322929 => x"FF",
		322930 => x"FF",
		322931 => x"FF",
		322932 => x"FF",
		323053 => x"FF",
		323054 => x"FF",
		323055 => x"FF",
		323056 => x"FF",
		323057 => x"FF",
		323702 => x"FF",
		323703 => x"FF",
		323704 => x"FF",
		323705 => x"FF",
		323706 => x"FF",
		323827 => x"FF",
		323828 => x"FF",
		323829 => x"FF",
		323830 => x"FF",
		323831 => x"FF",
		323952 => x"FF",
		323953 => x"FF",
		323954 => x"FF",
		323955 => x"FF",
		323956 => x"FF",
		324077 => x"FF",
		324078 => x"FF",
		324079 => x"FF",
		324080 => x"FF",
		324081 => x"FF",
		324726 => x"FF",
		324727 => x"FF",
		324728 => x"FF",
		324729 => x"FF",
		324730 => x"FF",
		324851 => x"FF",
		324852 => x"FF",
		324853 => x"FF",
		324854 => x"FF",
		324855 => x"FF",
		324976 => x"FF",
		324977 => x"FF",
		324978 => x"FF",
		324979 => x"FF",
		324980 => x"FF",
		325101 => x"FF",
		325102 => x"FF",
		325103 => x"FF",
		325104 => x"FF",
		325105 => x"FF",
		325750 => x"FF",
		325751 => x"FF",
		325752 => x"FF",
		325753 => x"FF",
		325754 => x"FF",
		325875 => x"FF",
		325876 => x"FF",
		325877 => x"FF",
		325878 => x"FF",
		325879 => x"FF",
		326000 => x"FF",
		326001 => x"FF",
		326002 => x"FF",
		326003 => x"FF",
		326004 => x"FF",
		326125 => x"FF",
		326126 => x"FF",
		326127 => x"FF",
		326128 => x"FF",
		326129 => x"FF",
		326774 => x"FF",
		326775 => x"FF",
		326776 => x"FF",
		326777 => x"FF",
		326778 => x"FF",
		326899 => x"FF",
		326900 => x"FF",
		326901 => x"FF",
		326902 => x"FF",
		326903 => x"FF",
		327024 => x"FF",
		327025 => x"FF",
		327026 => x"FF",
		327027 => x"FF",
		327028 => x"FF",
		327149 => x"FF",
		327150 => x"FF",
		327151 => x"FF",
		327152 => x"FF",
		327153 => x"FF",
		327798 => x"FF",
		327799 => x"FF",
		327800 => x"FF",
		327801 => x"FF",
		327802 => x"FF",
		327923 => x"FF",
		327924 => x"FF",
		327925 => x"FF",
		327926 => x"FF",
		327927 => x"FF",
		328048 => x"FF",
		328049 => x"FF",
		328050 => x"FF",
		328051 => x"FF",
		328052 => x"FF",
		328173 => x"FF",
		328174 => x"FF",
		328175 => x"FF",
		328176 => x"FF",
		328177 => x"FF",
		328822 => x"FF",
		328823 => x"FF",
		328824 => x"FF",
		328825 => x"FF",
		328826 => x"FF",
		328947 => x"FF",
		328948 => x"FF",
		328949 => x"FF",
		328950 => x"FF",
		328951 => x"FF",
		329072 => x"FF",
		329073 => x"FF",
		329074 => x"FF",
		329075 => x"FF",
		329076 => x"FF",
		329197 => x"FF",
		329198 => x"FF",
		329199 => x"FF",
		329200 => x"FF",
		329201 => x"FF",
		329846 => x"FF",
		329847 => x"FF",
		329848 => x"FF",
		329849 => x"FF",
		329850 => x"FF",
		329971 => x"FF",
		329972 => x"FF",
		329973 => x"FF",
		329974 => x"FF",
		329975 => x"FF",
		330096 => x"FF",
		330097 => x"FF",
		330098 => x"FF",
		330099 => x"FF",
		330100 => x"FF",
		330221 => x"FF",
		330222 => x"FF",
		330223 => x"FF",
		330224 => x"FF",
		330225 => x"FF",
		330870 => x"FF",
		330871 => x"FF",
		330872 => x"FF",
		330873 => x"FF",
		330874 => x"FF",
		330995 => x"FF",
		330996 => x"FF",
		330997 => x"FF",
		330998 => x"FF",
		330999 => x"FF",
		331120 => x"FF",
		331121 => x"FF",
		331122 => x"FF",
		331123 => x"FF",
		331124 => x"FF",
		331245 => x"FF",
		331246 => x"FF",
		331247 => x"FF",
		331248 => x"FF",
		331249 => x"FF",
		331894 => x"FF",
		331895 => x"FF",
		331896 => x"FF",
		331897 => x"FF",
		331898 => x"FF",
		332019 => x"FF",
		332020 => x"FF",
		332021 => x"FF",
		332022 => x"FF",
		332023 => x"FF",
		332144 => x"FF",
		332145 => x"FF",
		332146 => x"FF",
		332147 => x"FF",
		332148 => x"FF",
		332269 => x"FF",
		332270 => x"FF",
		332271 => x"FF",
		332272 => x"FF",
		332273 => x"FF",
		332918 => x"FF",
		332919 => x"FF",
		332920 => x"FF",
		332921 => x"FF",
		332922 => x"FF",
		333043 => x"FF",
		333044 => x"FF",
		333045 => x"FF",
		333046 => x"FF",
		333047 => x"FF",
		333168 => x"FF",
		333169 => x"FF",
		333170 => x"FF",
		333171 => x"FF",
		333172 => x"FF",
		333293 => x"FF",
		333294 => x"FF",
		333295 => x"FF",
		333296 => x"FF",
		333297 => x"FF",
		333942 => x"FF",
		333943 => x"FF",
		333944 => x"FF",
		333945 => x"FF",
		333946 => x"FF",
		334067 => x"FF",
		334068 => x"FF",
		334069 => x"FF",
		334070 => x"FF",
		334071 => x"FF",
		334192 => x"FF",
		334193 => x"FF",
		334194 => x"FF",
		334195 => x"FF",
		334196 => x"FF",
		334317 => x"FF",
		334318 => x"FF",
		334319 => x"FF",
		334320 => x"FF",
		334321 => x"FF",
		334966 => x"FF",
		334967 => x"FF",
		334968 => x"FF",
		334969 => x"FF",
		334970 => x"FF",
		335091 => x"FF",
		335092 => x"FF",
		335093 => x"FF",
		335094 => x"FF",
		335095 => x"FF",
		335216 => x"FF",
		335217 => x"FF",
		335218 => x"FF",
		335219 => x"FF",
		335220 => x"FF",
		335341 => x"FF",
		335342 => x"FF",
		335343 => x"FF",
		335344 => x"FF",
		335345 => x"FF",
		335990 => x"FF",
		335991 => x"FF",
		335992 => x"FF",
		335993 => x"FF",
		335994 => x"FF",
		336115 => x"FF",
		336116 => x"FF",
		336117 => x"FF",
		336118 => x"FF",
		336119 => x"FF",
		336240 => x"FF",
		336241 => x"FF",
		336242 => x"FF",
		336243 => x"FF",
		336244 => x"FF",
		336365 => x"FF",
		336366 => x"FF",
		336367 => x"FF",
		336368 => x"FF",
		336369 => x"FF",
		337014 => x"FF",
		337015 => x"FF",
		337016 => x"FF",
		337017 => x"FF",
		337018 => x"FF",
		337139 => x"FF",
		337140 => x"FF",
		337141 => x"FF",
		337142 => x"FF",
		337143 => x"FF",
		337264 => x"FF",
		337265 => x"FF",
		337266 => x"FF",
		337267 => x"FF",
		337268 => x"FF",
		337389 => x"FF",
		337390 => x"FF",
		337391 => x"FF",
		337392 => x"FF",
		337393 => x"FF",
		338038 => x"FF",
		338039 => x"FF",
		338040 => x"FF",
		338041 => x"FF",
		338042 => x"FF",
		338163 => x"FF",
		338164 => x"FF",
		338165 => x"FF",
		338166 => x"FF",
		338167 => x"FF",
		338288 => x"FF",
		338289 => x"FF",
		338290 => x"FF",
		338291 => x"FF",
		338292 => x"FF",
		338413 => x"FF",
		338414 => x"FF",
		338415 => x"FF",
		338416 => x"FF",
		338417 => x"FF",
		339062 => x"FF",
		339063 => x"FF",
		339064 => x"FF",
		339065 => x"FF",
		339066 => x"FF",
		339187 => x"FF",
		339188 => x"FF",
		339189 => x"FF",
		339190 => x"FF",
		339191 => x"FF",
		339312 => x"FF",
		339313 => x"FF",
		339314 => x"FF",
		339315 => x"FF",
		339316 => x"FF",
		339437 => x"FF",
		339438 => x"FF",
		339439 => x"FF",
		339440 => x"FF",
		339441 => x"FF",
		340086 => x"FF",
		340087 => x"FF",
		340088 => x"FF",
		340089 => x"FF",
		340090 => x"FF",
		340211 => x"FF",
		340212 => x"FF",
		340213 => x"FF",
		340214 => x"FF",
		340215 => x"FF",
		340336 => x"FF",
		340337 => x"FF",
		340338 => x"FF",
		340339 => x"FF",
		340340 => x"FF",
		340461 => x"FF",
		340462 => x"FF",
		340463 => x"FF",
		340464 => x"FF",
		340465 => x"FF",
		341110 => x"FF",
		341111 => x"FF",
		341112 => x"FF",
		341113 => x"FF",
		341114 => x"FF",
		341235 => x"FF",
		341236 => x"FF",
		341237 => x"FF",
		341238 => x"FF",
		341239 => x"FF",
		341360 => x"FF",
		341361 => x"FF",
		341362 => x"FF",
		341363 => x"FF",
		341364 => x"FF",
		341485 => x"FF",
		341486 => x"FF",
		341487 => x"FF",
		341488 => x"FF",
		341489 => x"FF",
		342134 => x"FF",
		342135 => x"FF",
		342136 => x"FF",
		342137 => x"FF",
		342138 => x"FF",
		342259 => x"FF",
		342260 => x"FF",
		342261 => x"FF",
		342262 => x"FF",
		342263 => x"FF",
		342384 => x"FF",
		342385 => x"FF",
		342386 => x"FF",
		342387 => x"FF",
		342388 => x"FF",
		342509 => x"FF",
		342510 => x"FF",
		342511 => x"FF",
		342512 => x"FF",
		342513 => x"FF",
		343158 => x"FF",
		343159 => x"FF",
		343160 => x"FF",
		343161 => x"FF",
		343162 => x"FF",
		343283 => x"FF",
		343284 => x"FF",
		343285 => x"FF",
		343286 => x"FF",
		343287 => x"FF",
		343408 => x"FF",
		343409 => x"FF",
		343410 => x"FF",
		343411 => x"FF",
		343412 => x"FF",
		343533 => x"FF",
		343534 => x"FF",
		343535 => x"FF",
		343536 => x"FF",
		343537 => x"FF",
		344182 => x"FF",
		344183 => x"FF",
		344184 => x"FF",
		344185 => x"FF",
		344186 => x"FF",
		344307 => x"FF",
		344308 => x"FF",
		344309 => x"FF",
		344310 => x"FF",
		344311 => x"FF",
		344432 => x"FF",
		344433 => x"FF",
		344434 => x"FF",
		344435 => x"FF",
		344436 => x"FF",
		344557 => x"FF",
		344558 => x"FF",
		344559 => x"FF",
		344560 => x"FF",
		344561 => x"FF",
		345206 => x"FF",
		345207 => x"FF",
		345208 => x"FF",
		345209 => x"FF",
		345210 => x"FF",
		345331 => x"FF",
		345332 => x"FF",
		345333 => x"FF",
		345334 => x"FF",
		345335 => x"FF",
		345456 => x"FF",
		345457 => x"FF",
		345458 => x"FF",
		345459 => x"FF",
		345460 => x"FF",
		345581 => x"FF",
		345582 => x"FF",
		345583 => x"FF",
		345584 => x"FF",
		345585 => x"FF",
		346230 => x"FF",
		346231 => x"FF",
		346232 => x"FF",
		346233 => x"FF",
		346234 => x"FF",
		346355 => x"FF",
		346356 => x"FF",
		346357 => x"FF",
		346358 => x"FF",
		346359 => x"FF",
		346480 => x"FF",
		346481 => x"FF",
		346482 => x"FF",
		346483 => x"FF",
		346484 => x"FF",
		346605 => x"FF",
		346606 => x"FF",
		346607 => x"FF",
		346608 => x"FF",
		346609 => x"FF",
		347254 => x"FF",
		347255 => x"FF",
		347256 => x"FF",
		347257 => x"FF",
		347258 => x"FF",
		347379 => x"FF",
		347380 => x"FF",
		347381 => x"FF",
		347382 => x"FF",
		347383 => x"FF",
		347504 => x"FF",
		347505 => x"FF",
		347506 => x"FF",
		347507 => x"FF",
		347508 => x"FF",
		347629 => x"FF",
		347630 => x"FF",
		347631 => x"FF",
		347632 => x"FF",
		347633 => x"FF",
		348278 => x"FF",
		348279 => x"FF",
		348280 => x"FF",
		348281 => x"FF",
		348282 => x"FF",
		348403 => x"FF",
		348404 => x"FF",
		348405 => x"FF",
		348406 => x"FF",
		348407 => x"FF",
		348528 => x"FF",
		348529 => x"FF",
		348530 => x"FF",
		348531 => x"FF",
		348532 => x"FF",
		348653 => x"FF",
		348654 => x"FF",
		348655 => x"FF",
		348656 => x"FF",
		348657 => x"FF",
		349302 => x"FF",
		349303 => x"FF",
		349304 => x"FF",
		349305 => x"FF",
		349306 => x"FF",
		349427 => x"FF",
		349428 => x"FF",
		349429 => x"FF",
		349430 => x"FF",
		349431 => x"FF",
		349552 => x"FF",
		349553 => x"FF",
		349554 => x"FF",
		349555 => x"FF",
		349556 => x"FF",
		349677 => x"FF",
		349678 => x"FF",
		349679 => x"FF",
		349680 => x"FF",
		349681 => x"FF",
		350326 => x"FF",
		350327 => x"FF",
		350328 => x"FF",
		350329 => x"FF",
		350330 => x"FF",
		350451 => x"FF",
		350452 => x"FF",
		350453 => x"FF",
		350454 => x"FF",
		350455 => x"FF",
		350576 => x"FF",
		350577 => x"FF",
		350578 => x"FF",
		350579 => x"FF",
		350580 => x"FF",
		350701 => x"FF",
		350702 => x"FF",
		350703 => x"FF",
		350704 => x"FF",
		350705 => x"FF",
		351350 => x"FF",
		351351 => x"FF",
		351352 => x"FF",
		351353 => x"FF",
		351354 => x"FF",
		351475 => x"FF",
		351476 => x"FF",
		351477 => x"FF",
		351478 => x"FF",
		351479 => x"FF",
		351600 => x"FF",
		351601 => x"FF",
		351602 => x"FF",
		351603 => x"FF",
		351604 => x"FF",
		351725 => x"FF",
		351726 => x"FF",
		351727 => x"FF",
		351728 => x"FF",
		351729 => x"FF",
		352374 => x"FF",
		352375 => x"FF",
		352376 => x"FF",
		352377 => x"FF",
		352378 => x"FF",
		352499 => x"FF",
		352500 => x"FF",
		352501 => x"FF",
		352502 => x"FF",
		352503 => x"FF",
		352624 => x"FF",
		352625 => x"FF",
		352626 => x"FF",
		352627 => x"FF",
		352628 => x"FF",
		352749 => x"FF",
		352750 => x"FF",
		352751 => x"FF",
		352752 => x"FF",
		352753 => x"FF",
		353398 => x"FF",
		353399 => x"FF",
		353400 => x"FF",
		353401 => x"FF",
		353402 => x"FF",
		353523 => x"FF",
		353524 => x"FF",
		353525 => x"FF",
		353526 => x"FF",
		353527 => x"FF",
		353648 => x"FF",
		353649 => x"FF",
		353650 => x"FF",
		353651 => x"FF",
		353652 => x"FF",
		353773 => x"FF",
		353774 => x"FF",
		353775 => x"FF",
		353776 => x"FF",
		353777 => x"FF",
		354422 => x"FF",
		354423 => x"FF",
		354424 => x"FF",
		354425 => x"FF",
		354426 => x"FF",
		354547 => x"FF",
		354548 => x"FF",
		354549 => x"FF",
		354550 => x"FF",
		354551 => x"FF",
		354672 => x"FF",
		354673 => x"FF",
		354674 => x"FF",
		354675 => x"FF",
		354676 => x"FF",
		354797 => x"FF",
		354798 => x"FF",
		354799 => x"FF",
		354800 => x"FF",
		354801 => x"FF",
		355446 => x"FF",
		355447 => x"FF",
		355448 => x"FF",
		355449 => x"FF",
		355450 => x"FF",
		355571 => x"FF",
		355572 => x"FF",
		355573 => x"FF",
		355574 => x"FF",
		355575 => x"FF",
		355696 => x"FF",
		355697 => x"FF",
		355698 => x"FF",
		355699 => x"FF",
		355700 => x"FF",
		355821 => x"FF",
		355822 => x"FF",
		355823 => x"FF",
		355824 => x"FF",
		355825 => x"FF",
		356470 => x"FF",
		356471 => x"FF",
		356472 => x"FF",
		356473 => x"FF",
		356474 => x"FF",
		356595 => x"FF",
		356596 => x"FF",
		356597 => x"FF",
		356598 => x"FF",
		356599 => x"FF",
		356720 => x"FF",
		356721 => x"FF",
		356722 => x"FF",
		356723 => x"FF",
		356724 => x"FF",
		356845 => x"FF",
		356846 => x"FF",
		356847 => x"FF",
		356848 => x"FF",
		356849 => x"FF",
		357494 => x"FF",
		357495 => x"FF",
		357496 => x"FF",
		357497 => x"FF",
		357498 => x"FF",
		357619 => x"FF",
		357620 => x"FF",
		357621 => x"FF",
		357622 => x"FF",
		357623 => x"FF",
		357744 => x"FF",
		357745 => x"FF",
		357746 => x"FF",
		357747 => x"FF",
		357748 => x"FF",
		357869 => x"FF",
		357870 => x"FF",
		357871 => x"FF",
		357872 => x"FF",
		357873 => x"FF",
		358518 => x"FF",
		358519 => x"FF",
		358520 => x"FF",
		358521 => x"FF",
		358522 => x"FF",
		358643 => x"FF",
		358644 => x"FF",
		358645 => x"FF",
		358646 => x"FF",
		358647 => x"FF",
		358768 => x"FF",
		358769 => x"FF",
		358770 => x"FF",
		358771 => x"FF",
		358772 => x"FF",
		358893 => x"FF",
		358894 => x"FF",
		358895 => x"FF",
		358896 => x"FF",
		358897 => x"FF",
		359542 => x"FF",
		359543 => x"FF",
		359544 => x"FF",
		359545 => x"FF",
		359546 => x"FF",
		359667 => x"FF",
		359668 => x"FF",
		359669 => x"FF",
		359670 => x"FF",
		359671 => x"FF",
		359792 => x"FF",
		359793 => x"FF",
		359794 => x"FF",
		359795 => x"FF",
		359796 => x"FF",
		359917 => x"FF",
		359918 => x"FF",
		359919 => x"FF",
		359920 => x"FF",
		359921 => x"FF",
		360566 => x"FF",
		360567 => x"FF",
		360568 => x"FF",
		360569 => x"FF",
		360570 => x"FF",
		360691 => x"FF",
		360692 => x"FF",
		360693 => x"FF",
		360694 => x"FF",
		360695 => x"FF",
		360816 => x"FF",
		360817 => x"FF",
		360818 => x"FF",
		360819 => x"FF",
		360820 => x"FF",
		360941 => x"FF",
		360942 => x"FF",
		360943 => x"FF",
		360944 => x"FF",
		360945 => x"FF",
		361590 => x"FF",
		361591 => x"FF",
		361592 => x"FF",
		361593 => x"FF",
		361594 => x"FF",
		361715 => x"FF",
		361716 => x"FF",
		361717 => x"FF",
		361718 => x"FF",
		361719 => x"FF",
		361840 => x"FF",
		361841 => x"FF",
		361842 => x"FF",
		361843 => x"FF",
		361844 => x"FF",
		361965 => x"FF",
		361966 => x"FF",
		361967 => x"FF",
		361968 => x"FF",
		361969 => x"FF",
		362614 => x"FF",
		362615 => x"FF",
		362616 => x"FF",
		362617 => x"FF",
		362618 => x"FF",
		362739 => x"FF",
		362740 => x"FF",
		362741 => x"FF",
		362742 => x"FF",
		362743 => x"FF",
		362864 => x"FF",
		362865 => x"FF",
		362866 => x"FF",
		362867 => x"FF",
		362868 => x"FF",
		362989 => x"FF",
		362990 => x"FF",
		362991 => x"FF",
		362992 => x"FF",
		362993 => x"FF",
		363638 => x"FF",
		363639 => x"FF",
		363640 => x"FF",
		363641 => x"FF",
		363642 => x"FF",
		363763 => x"FF",
		363764 => x"FF",
		363765 => x"FF",
		363766 => x"FF",
		363767 => x"FF",
		363888 => x"FF",
		363889 => x"FF",
		363890 => x"FF",
		363891 => x"FF",
		363892 => x"FF",
		364013 => x"FF",
		364014 => x"FF",
		364015 => x"FF",
		364016 => x"FF",
		364017 => x"FF",
		364662 => x"FF",
		364663 => x"FF",
		364664 => x"FF",
		364665 => x"FF",
		364666 => x"FF",
		364787 => x"FF",
		364788 => x"FF",
		364789 => x"FF",
		364790 => x"FF",
		364791 => x"FF",
		364912 => x"FF",
		364913 => x"FF",
		364914 => x"FF",
		364915 => x"FF",
		364916 => x"FF",
		365037 => x"FF",
		365038 => x"FF",
		365039 => x"FF",
		365040 => x"FF",
		365041 => x"FF",
		365686 => x"FF",
		365687 => x"FF",
		365688 => x"FF",
		365689 => x"FF",
		365690 => x"FF",
		365811 => x"FF",
		365812 => x"FF",
		365813 => x"FF",
		365814 => x"FF",
		365815 => x"FF",
		365936 => x"FF",
		365937 => x"FF",
		365938 => x"FF",
		365939 => x"FF",
		365940 => x"FF",
		366061 => x"FF",
		366062 => x"FF",
		366063 => x"FF",
		366064 => x"FF",
		366065 => x"FF",
		366710 => x"FF",
		366711 => x"FF",
		366712 => x"FF",
		366713 => x"FF",
		366714 => x"FF",
		366835 => x"FF",
		366836 => x"FF",
		366837 => x"FF",
		366838 => x"FF",
		366839 => x"FF",
		366960 => x"FF",
		366961 => x"FF",
		366962 => x"FF",
		366963 => x"FF",
		366964 => x"FF",
		367085 => x"FF",
		367086 => x"FF",
		367087 => x"FF",
		367088 => x"FF",
		367089 => x"FF",
		367734 => x"FF",
		367735 => x"FF",
		367736 => x"FF",
		367737 => x"FF",
		367738 => x"FF",
		367859 => x"FF",
		367860 => x"FF",
		367861 => x"FF",
		367862 => x"FF",
		367863 => x"FF",
		367984 => x"FF",
		367985 => x"FF",
		367986 => x"FF",
		367987 => x"FF",
		367988 => x"FF",
		368109 => x"FF",
		368110 => x"FF",
		368111 => x"FF",
		368112 => x"FF",
		368113 => x"FF",
		368758 => x"FF",
		368759 => x"FF",
		368760 => x"FF",
		368761 => x"FF",
		368762 => x"FF",
		368883 => x"FF",
		368884 => x"FF",
		368885 => x"FF",
		368886 => x"FF",
		368887 => x"FF",
		369008 => x"FF",
		369009 => x"FF",
		369010 => x"FF",
		369011 => x"FF",
		369012 => x"FF",
		369133 => x"FF",
		369134 => x"FF",
		369135 => x"FF",
		369136 => x"FF",
		369137 => x"FF",
		369782 => x"FF",
		369783 => x"FF",
		369784 => x"FF",
		369785 => x"FF",
		369786 => x"FF",
		369907 => x"FF",
		369908 => x"FF",
		369909 => x"FF",
		369910 => x"FF",
		369911 => x"FF",
		370032 => x"FF",
		370033 => x"FF",
		370034 => x"FF",
		370035 => x"FF",
		370036 => x"FF",
		370157 => x"FF",
		370158 => x"FF",
		370159 => x"FF",
		370160 => x"FF",
		370161 => x"FF",
		370806 => x"FF",
		370807 => x"FF",
		370808 => x"FF",
		370809 => x"FF",
		370810 => x"FF",
		370931 => x"FF",
		370932 => x"FF",
		370933 => x"FF",
		370934 => x"FF",
		370935 => x"FF",
		371056 => x"FF",
		371057 => x"FF",
		371058 => x"FF",
		371059 => x"FF",
		371060 => x"FF",
		371181 => x"FF",
		371182 => x"FF",
		371183 => x"FF",
		371184 => x"FF",
		371185 => x"FF",
		371830 => x"FF",
		371831 => x"FF",
		371832 => x"FF",
		371833 => x"FF",
		371834 => x"FF",
		371955 => x"FF",
		371956 => x"FF",
		371957 => x"FF",
		371958 => x"FF",
		371959 => x"FF",
		372080 => x"FF",
		372081 => x"FF",
		372082 => x"FF",
		372083 => x"FF",
		372084 => x"FF",
		372205 => x"FF",
		372206 => x"FF",
		372207 => x"FF",
		372208 => x"FF",
		372209 => x"FF",
		372854 => x"FF",
		372855 => x"FF",
		372856 => x"FF",
		372857 => x"FF",
		372858 => x"FF",
		372979 => x"FF",
		372980 => x"FF",
		372981 => x"FF",
		372982 => x"FF",
		372983 => x"FF",
		373104 => x"FF",
		373105 => x"FF",
		373106 => x"FF",
		373107 => x"FF",
		373108 => x"FF",
		373229 => x"FF",
		373230 => x"FF",
		373231 => x"FF",
		373232 => x"FF",
		373233 => x"FF",
		373878 => x"FF",
		373879 => x"FF",
		373880 => x"FF",
		373881 => x"FF",
		373882 => x"FF",
		374003 => x"FF",
		374004 => x"FF",
		374005 => x"FF",
		374006 => x"FF",
		374007 => x"FF",
		374128 => x"FF",
		374129 => x"FF",
		374130 => x"FF",
		374131 => x"FF",
		374132 => x"FF",
		374253 => x"FF",
		374254 => x"FF",
		374255 => x"FF",
		374256 => x"FF",
		374257 => x"FF",
		374902 => x"FF",
		374903 => x"FF",
		374904 => x"FF",
		374905 => x"FF",
		374906 => x"FF",
		375027 => x"FF",
		375028 => x"FF",
		375029 => x"FF",
		375030 => x"FF",
		375031 => x"FF",
		375152 => x"FF",
		375153 => x"FF",
		375154 => x"FF",
		375155 => x"FF",
		375156 => x"FF",
		375277 => x"FF",
		375278 => x"FF",
		375279 => x"FF",
		375280 => x"FF",
		375281 => x"FF",
		375926 => x"FF",
		375927 => x"FF",
		375928 => x"FF",
		375929 => x"FF",
		375930 => x"FF",
		376051 => x"FF",
		376052 => x"FF",
		376053 => x"FF",
		376054 => x"FF",
		376055 => x"FF",
		376176 => x"FF",
		376177 => x"FF",
		376178 => x"FF",
		376179 => x"FF",
		376180 => x"FF",
		376301 => x"FF",
		376302 => x"FF",
		376303 => x"FF",
		376304 => x"FF",
		376305 => x"FF",
		376950 => x"FF",
		376951 => x"FF",
		376952 => x"FF",
		376953 => x"FF",
		376954 => x"FF",
		377075 => x"FF",
		377076 => x"FF",
		377077 => x"FF",
		377078 => x"FF",
		377079 => x"FF",
		377200 => x"FF",
		377201 => x"FF",
		377202 => x"FF",
		377203 => x"FF",
		377204 => x"FF",
		377325 => x"FF",
		377326 => x"FF",
		377327 => x"FF",
		377328 => x"FF",
		377329 => x"FF",
		377974 => x"FF",
		377975 => x"FF",
		377976 => x"FF",
		377977 => x"FF",
		377978 => x"FF",
		378099 => x"FF",
		378100 => x"FF",
		378101 => x"FF",
		378102 => x"FF",
		378103 => x"FF",
		378224 => x"FF",
		378225 => x"FF",
		378226 => x"FF",
		378227 => x"FF",
		378228 => x"FF",
		378349 => x"FF",
		378350 => x"FF",
		378351 => x"FF",
		378352 => x"FF",
		378353 => x"FF",
		378998 => x"FF",
		378999 => x"FF",
		379000 => x"FF",
		379001 => x"FF",
		379002 => x"FF",
		379123 => x"FF",
		379124 => x"FF",
		379125 => x"FF",
		379126 => x"FF",
		379127 => x"FF",
		379248 => x"FF",
		379249 => x"FF",
		379250 => x"FF",
		379251 => x"FF",
		379252 => x"FF",
		379373 => x"FF",
		379374 => x"FF",
		379375 => x"FF",
		379376 => x"FF",
		379377 => x"FF",
		380022 => x"FF",
		380023 => x"FF",
		380024 => x"FF",
		380025 => x"FF",
		380026 => x"FF",
		380147 => x"FF",
		380148 => x"FF",
		380149 => x"FF",
		380150 => x"FF",
		380151 => x"FF",
		380272 => x"FF",
		380273 => x"FF",
		380274 => x"FF",
		380275 => x"FF",
		380276 => x"FF",
		380397 => x"FF",
		380398 => x"FF",
		380399 => x"FF",
		380400 => x"FF",
		380401 => x"FF",
		381046 => x"FF",
		381047 => x"FF",
		381048 => x"FF",
		381049 => x"FF",
		381050 => x"FF",
		381171 => x"FF",
		381172 => x"FF",
		381173 => x"FF",
		381174 => x"FF",
		381175 => x"FF",
		381296 => x"FF",
		381297 => x"FF",
		381298 => x"FF",
		381299 => x"FF",
		381300 => x"FF",
		381421 => x"FF",
		381422 => x"FF",
		381423 => x"FF",
		381424 => x"FF",
		381425 => x"FF",
		382070 => x"FF",
		382071 => x"FF",
		382072 => x"FF",
		382073 => x"FF",
		382074 => x"FF",
		382195 => x"FF",
		382196 => x"FF",
		382197 => x"FF",
		382198 => x"FF",
		382199 => x"FF",
		382320 => x"FF",
		382321 => x"FF",
		382322 => x"FF",
		382323 => x"FF",
		382324 => x"FF",
		382445 => x"FF",
		382446 => x"FF",
		382447 => x"FF",
		382448 => x"FF",
		382449 => x"FF",
		383094 => x"FF",
		383095 => x"FF",
		383096 => x"FF",
		383097 => x"FF",
		383098 => x"FF",
		383219 => x"FF",
		383220 => x"FF",
		383221 => x"FF",
		383222 => x"FF",
		383223 => x"FF",
		383344 => x"FF",
		383345 => x"FF",
		383346 => x"FF",
		383347 => x"FF",
		383348 => x"FF",
		383469 => x"FF",
		383470 => x"FF",
		383471 => x"FF",
		383472 => x"FF",
		383473 => x"FF",
		384118 => x"FF",
		384119 => x"FF",
		384120 => x"FF",
		384121 => x"FF",
		384122 => x"FF",
		384243 => x"FF",
		384244 => x"FF",
		384245 => x"FF",
		384246 => x"FF",
		384247 => x"FF",
		384368 => x"FF",
		384369 => x"FF",
		384370 => x"FF",
		384371 => x"FF",
		384372 => x"FF",
		384493 => x"FF",
		384494 => x"FF",
		384495 => x"FF",
		384496 => x"FF",
		384497 => x"FF",
		385142 => x"FF",
		385143 => x"FF",
		385144 => x"FF",
		385145 => x"FF",
		385146 => x"FF",
		385267 => x"FF",
		385268 => x"FF",
		385269 => x"FF",
		385270 => x"FF",
		385271 => x"FF",
		385392 => x"FF",
		385393 => x"FF",
		385394 => x"FF",
		385395 => x"FF",
		385396 => x"FF",
		385517 => x"FF",
		385518 => x"FF",
		385519 => x"FF",
		385520 => x"FF",
		385521 => x"FF",
		386166 => x"FF",
		386167 => x"FF",
		386168 => x"FF",
		386169 => x"FF",
		386170 => x"FF",
		386291 => x"FF",
		386292 => x"FF",
		386293 => x"FF",
		386294 => x"FF",
		386295 => x"FF",
		386416 => x"FF",
		386417 => x"FF",
		386418 => x"FF",
		386419 => x"FF",
		386420 => x"FF",
		386541 => x"FF",
		386542 => x"FF",
		386543 => x"FF",
		386544 => x"FF",
		386545 => x"FF",
		387190 => x"FF",
		387191 => x"FF",
		387192 => x"FF",
		387193 => x"FF",
		387194 => x"FF",
		387315 => x"FF",
		387316 => x"FF",
		387317 => x"FF",
		387318 => x"FF",
		387319 => x"FF",
		387440 => x"FF",
		387441 => x"FF",
		387442 => x"FF",
		387443 => x"FF",
		387444 => x"FF",
		387565 => x"FF",
		387566 => x"FF",
		387567 => x"FF",
		387568 => x"FF",
		387569 => x"FF",
		388214 => x"FF",
		388215 => x"FF",
		388216 => x"FF",
		388217 => x"FF",
		388218 => x"FF",
		388339 => x"FF",
		388340 => x"FF",
		388341 => x"FF",
		388342 => x"FF",
		388343 => x"FF",
		388464 => x"FF",
		388465 => x"FF",
		388466 => x"FF",
		388467 => x"FF",
		388468 => x"FF",
		388589 => x"FF",
		388590 => x"FF",
		388591 => x"FF",
		388592 => x"FF",
		388593 => x"FF",
		389238 => x"FF",
		389239 => x"FF",
		389240 => x"FF",
		389241 => x"FF",
		389242 => x"FF",
		389363 => x"FF",
		389364 => x"FF",
		389365 => x"FF",
		389366 => x"FF",
		389367 => x"FF",
		389488 => x"FF",
		389489 => x"FF",
		389490 => x"FF",
		389491 => x"FF",
		389492 => x"FF",
		389613 => x"FF",
		389614 => x"FF",
		389615 => x"FF",
		389616 => x"FF",
		389617 => x"FF",
		390262 => x"FF",
		390263 => x"FF",
		390264 => x"FF",
		390265 => x"FF",
		390266 => x"FF",
		390387 => x"FF",
		390388 => x"FF",
		390389 => x"FF",
		390390 => x"FF",
		390391 => x"FF",
		390512 => x"FF",
		390513 => x"FF",
		390514 => x"FF",
		390515 => x"FF",
		390516 => x"FF",
		390637 => x"FF",
		390638 => x"FF",
		390639 => x"FF",
		390640 => x"FF",
		390641 => x"FF",
		391286 => x"FF",
		391287 => x"FF",
		391288 => x"FF",
		391289 => x"FF",
		391290 => x"FF",
		391411 => x"FF",
		391412 => x"FF",
		391413 => x"FF",
		391414 => x"FF",
		391415 => x"FF",
		391536 => x"FF",
		391537 => x"FF",
		391538 => x"FF",
		391539 => x"FF",
		391540 => x"FF",
		391661 => x"FF",
		391662 => x"FF",
		391663 => x"FF",
		391664 => x"FF",
		391665 => x"FF",
		392310 => x"FF",
		392311 => x"FF",
		392312 => x"FF",
		392313 => x"FF",
		392314 => x"FF",
		392435 => x"FF",
		392436 => x"FF",
		392437 => x"FF",
		392438 => x"FF",
		392439 => x"FF",
		392560 => x"FF",
		392561 => x"FF",
		392562 => x"FF",
		392563 => x"FF",
		392564 => x"FF",
		392685 => x"FF",
		392686 => x"FF",
		392687 => x"FF",
		392688 => x"FF",
		392689 => x"FF",
		393334 => x"FF",
		393335 => x"FF",
		393336 => x"FF",
		393337 => x"FF",
		393338 => x"FF",
		393459 => x"FF",
		393460 => x"FF",
		393461 => x"FF",
		393462 => x"FF",
		393463 => x"FF",
		393584 => x"FF",
		393585 => x"FF",
		393586 => x"FF",
		393587 => x"FF",
		393588 => x"FF",
		393709 => x"FF",
		393710 => x"FF",
		393711 => x"FF",
		393712 => x"FF",
		393713 => x"FF",
		394358 => x"FF",
		394359 => x"FF",
		394360 => x"FF",
		394361 => x"FF",
		394362 => x"FF",
		394483 => x"FF",
		394484 => x"FF",
		394485 => x"FF",
		394486 => x"FF",
		394487 => x"FF",
		394608 => x"FF",
		394609 => x"FF",
		394610 => x"FF",
		394611 => x"FF",
		394612 => x"FF",
		394733 => x"FF",
		394734 => x"FF",
		394735 => x"FF",
		394736 => x"FF",
		394737 => x"FF",
		395382 => x"FF",
		395383 => x"FF",
		395384 => x"FF",
		395385 => x"FF",
		395386 => x"FF",
		395507 => x"FF",
		395508 => x"FF",
		395509 => x"FF",
		395510 => x"FF",
		395511 => x"FF",
		395632 => x"FF",
		395633 => x"FF",
		395634 => x"FF",
		395635 => x"FF",
		395636 => x"FF",
		395757 => x"FF",
		395758 => x"FF",
		395759 => x"FF",
		395760 => x"FF",
		395761 => x"FF",
		396406 => x"FF",
		396407 => x"FF",
		396408 => x"FF",
		396409 => x"FF",
		396410 => x"FF",
		396531 => x"FF",
		396532 => x"FF",
		396533 => x"FF",
		396534 => x"FF",
		396535 => x"FF",
		396656 => x"FF",
		396657 => x"FF",
		396658 => x"FF",
		396659 => x"FF",
		396660 => x"FF",
		396781 => x"FF",
		396782 => x"FF",
		396783 => x"FF",
		396784 => x"FF",
		396785 => x"FF",
		397430 => x"FF",
		397431 => x"FF",
		397432 => x"FF",
		397433 => x"FF",
		397434 => x"FF",
		397555 => x"FF",
		397556 => x"FF",
		397557 => x"FF",
		397558 => x"FF",
		397559 => x"FF",
		397680 => x"FF",
		397681 => x"FF",
		397682 => x"FF",
		397683 => x"FF",
		397684 => x"FF",
		397805 => x"FF",
		397806 => x"FF",
		397807 => x"FF",
		397808 => x"FF",
		397809 => x"FF",
		398454 => x"FF",
		398455 => x"FF",
		398456 => x"FF",
		398457 => x"FF",
		398458 => x"FF",
		398579 => x"FF",
		398580 => x"FF",
		398581 => x"FF",
		398582 => x"FF",
		398583 => x"FF",
		398704 => x"FF",
		398705 => x"FF",
		398706 => x"FF",
		398707 => x"FF",
		398708 => x"FF",
		398829 => x"FF",
		398830 => x"FF",
		398831 => x"FF",
		398832 => x"FF",
		398833 => x"FF",
		399478 => x"FF",
		399479 => x"FF",
		399480 => x"FF",
		399481 => x"FF",
		399482 => x"FF",
		399603 => x"FF",
		399604 => x"FF",
		399605 => x"FF",
		399606 => x"FF",
		399607 => x"FF",
		399728 => x"FF",
		399729 => x"FF",
		399730 => x"FF",
		399731 => x"FF",
		399732 => x"FF",
		399853 => x"FF",
		399854 => x"FF",
		399855 => x"FF",
		399856 => x"FF",
		399857 => x"FF",
		400502 => x"FF",
		400503 => x"FF",
		400504 => x"FF",
		400505 => x"FF",
		400506 => x"FF",
		400627 => x"FF",
		400628 => x"FF",
		400629 => x"FF",
		400630 => x"FF",
		400631 => x"FF",
		400752 => x"FF",
		400753 => x"FF",
		400754 => x"FF",
		400755 => x"FF",
		400756 => x"FF",
		400877 => x"FF",
		400878 => x"FF",
		400879 => x"FF",
		400880 => x"FF",
		400881 => x"FF",
		401526 => x"FF",
		401527 => x"FF",
		401528 => x"FF",
		401529 => x"FF",
		401530 => x"FF",
		401651 => x"FF",
		401652 => x"FF",
		401653 => x"FF",
		401654 => x"FF",
		401655 => x"FF",
		401776 => x"FF",
		401777 => x"FF",
		401778 => x"FF",
		401779 => x"FF",
		401780 => x"FF",
		401901 => x"FF",
		401902 => x"FF",
		401903 => x"FF",
		401904 => x"FF",
		401905 => x"FF",
		402550 => x"FF",
		402551 => x"FF",
		402552 => x"FF",
		402553 => x"FF",
		402554 => x"FF",
		402675 => x"FF",
		402676 => x"FF",
		402677 => x"FF",
		402678 => x"FF",
		402679 => x"FF",
		402800 => x"FF",
		402801 => x"FF",
		402802 => x"FF",
		402803 => x"FF",
		402804 => x"FF",
		402925 => x"FF",
		402926 => x"FF",
		402927 => x"FF",
		402928 => x"FF",
		402929 => x"FF",
		403574 => x"FF",
		403575 => x"FF",
		403576 => x"FF",
		403577 => x"FF",
		403578 => x"FF",
		403699 => x"FF",
		403700 => x"FF",
		403701 => x"FF",
		403702 => x"FF",
		403703 => x"FF",
		403824 => x"FF",
		403825 => x"FF",
		403826 => x"FF",
		403827 => x"FF",
		403828 => x"FF",
		403949 => x"FF",
		403950 => x"FF",
		403951 => x"FF",
		403952 => x"FF",
		403953 => x"FF",
		404598 => x"FF",
		404599 => x"FF",
		404600 => x"FF",
		404601 => x"FF",
		404602 => x"FF",
		404723 => x"FF",
		404724 => x"FF",
		404725 => x"FF",
		404726 => x"FF",
		404727 => x"FF",
		404848 => x"FF",
		404849 => x"FF",
		404850 => x"FF",
		404851 => x"FF",
		404852 => x"FF",
		404973 => x"FF",
		404974 => x"FF",
		404975 => x"FF",
		404976 => x"FF",
		404977 => x"FF",
		405622 => x"FF",
		405623 => x"FF",
		405624 => x"FF",
		405625 => x"FF",
		405626 => x"FF",
		405747 => x"FF",
		405748 => x"FF",
		405749 => x"FF",
		405750 => x"FF",
		405751 => x"FF",
		405872 => x"FF",
		405873 => x"FF",
		405874 => x"FF",
		405875 => x"FF",
		405876 => x"FF",
		405997 => x"FF",
		405998 => x"FF",
		405999 => x"FF",
		406000 => x"FF",
		406001 => x"FF",
		406646 => x"FF",
		406647 => x"FF",
		406648 => x"FF",
		406649 => x"FF",
		406650 => x"FF",
		406771 => x"FF",
		406772 => x"FF",
		406773 => x"FF",
		406774 => x"FF",
		406775 => x"FF",
		406896 => x"FF",
		406897 => x"FF",
		406898 => x"FF",
		406899 => x"FF",
		406900 => x"FF",
		407021 => x"FF",
		407022 => x"FF",
		407023 => x"FF",
		407024 => x"FF",
		407025 => x"FF",
		407670 => x"FF",
		407671 => x"FF",
		407672 => x"FF",
		407673 => x"FF",
		407674 => x"FF",
		407795 => x"FF",
		407796 => x"FF",
		407797 => x"FF",
		407798 => x"FF",
		407799 => x"FF",
		407920 => x"FF",
		407921 => x"FF",
		407922 => x"FF",
		407923 => x"FF",
		407924 => x"FF",
		408045 => x"FF",
		408046 => x"FF",
		408047 => x"FF",
		408048 => x"FF",
		408049 => x"FF",
		408694 => x"FF",
		408695 => x"FF",
		408696 => x"FF",
		408697 => x"FF",
		408698 => x"FF",
		408819 => x"FF",
		408820 => x"FF",
		408821 => x"FF",
		408822 => x"FF",
		408823 => x"FF",
		408944 => x"FF",
		408945 => x"FF",
		408946 => x"FF",
		408947 => x"FF",
		408948 => x"FF",
		409069 => x"FF",
		409070 => x"FF",
		409071 => x"FF",
		409072 => x"FF",
		409073 => x"FF",
		409718 => x"FF",
		409719 => x"FF",
		409720 => x"FF",
		409721 => x"FF",
		409722 => x"FF",
		409843 => x"FF",
		409844 => x"FF",
		409845 => x"FF",
		409846 => x"FF",
		409847 => x"FF",
		409968 => x"FF",
		409969 => x"FF",
		409970 => x"FF",
		409971 => x"FF",
		409972 => x"FF",
		410093 => x"FF",
		410094 => x"FF",
		410095 => x"FF",
		410096 => x"FF",
		410097 => x"FF",
		410742 => x"FF",
		410743 => x"FF",
		410744 => x"FF",
		410745 => x"FF",
		410746 => x"FF",
		410867 => x"FF",
		410868 => x"FF",
		410869 => x"FF",
		410870 => x"FF",
		410871 => x"FF",
		410992 => x"FF",
		410993 => x"FF",
		410994 => x"FF",
		410995 => x"FF",
		410996 => x"FF",
		411117 => x"FF",
		411118 => x"FF",
		411119 => x"FF",
		411120 => x"FF",
		411121 => x"FF",
		411766 => x"FF",
		411767 => x"FF",
		411768 => x"FF",
		411769 => x"FF",
		411770 => x"FF",
		411891 => x"FF",
		411892 => x"FF",
		411893 => x"FF",
		411894 => x"FF",
		411895 => x"FF",
		412016 => x"FF",
		412017 => x"FF",
		412018 => x"FF",
		412019 => x"FF",
		412020 => x"FF",
		412141 => x"FF",
		412142 => x"FF",
		412143 => x"FF",
		412144 => x"FF",
		412145 => x"FF",
		412790 => x"FF",
		412791 => x"FF",
		412792 => x"FF",
		412793 => x"FF",
		412794 => x"FF",
		412915 => x"FF",
		412916 => x"FF",
		412917 => x"FF",
		412918 => x"FF",
		412919 => x"FF",
		413040 => x"FF",
		413041 => x"FF",
		413042 => x"FF",
		413043 => x"FF",
		413044 => x"FF",
		413165 => x"FF",
		413166 => x"FF",
		413167 => x"FF",
		413168 => x"FF",
		413169 => x"FF",
		413814 => x"FF",
		413815 => x"FF",
		413816 => x"FF",
		413817 => x"FF",
		413818 => x"FF",
		413939 => x"FF",
		413940 => x"FF",
		413941 => x"FF",
		413942 => x"FF",
		413943 => x"FF",
		414064 => x"FF",
		414065 => x"FF",
		414066 => x"FF",
		414067 => x"FF",
		414068 => x"FF",
		414189 => x"FF",
		414190 => x"FF",
		414191 => x"FF",
		414192 => x"FF",
		414193 => x"FF",
		414838 => x"FF",
		414839 => x"FF",
		414840 => x"FF",
		414841 => x"FF",
		414842 => x"FF",
		414963 => x"FF",
		414964 => x"FF",
		414965 => x"FF",
		414966 => x"FF",
		414967 => x"FF",
		415088 => x"FF",
		415089 => x"FF",
		415090 => x"FF",
		415091 => x"FF",
		415092 => x"FF",
		415213 => x"FF",
		415214 => x"FF",
		415215 => x"FF",
		415216 => x"FF",
		415217 => x"FF",
		415862 => x"FF",
		415863 => x"FF",
		415864 => x"FF",
		415865 => x"FF",
		415866 => x"FF",
		415987 => x"FF",
		415988 => x"FF",
		415989 => x"FF",
		415990 => x"FF",
		415991 => x"FF",
		416112 => x"FF",
		416113 => x"FF",
		416114 => x"FF",
		416115 => x"FF",
		416116 => x"FF",
		416237 => x"FF",
		416238 => x"FF",
		416239 => x"FF",
		416240 => x"FF",
		416241 => x"FF",
		416886 => x"FF",
		416887 => x"FF",
		416888 => x"FF",
		416889 => x"FF",
		416890 => x"FF",
		417011 => x"FF",
		417012 => x"FF",
		417013 => x"FF",
		417014 => x"FF",
		417015 => x"FF",
		417136 => x"FF",
		417137 => x"FF",
		417138 => x"FF",
		417139 => x"FF",
		417140 => x"FF",
		417261 => x"FF",
		417262 => x"FF",
		417263 => x"FF",
		417264 => x"FF",
		417265 => x"FF",
		417910 => x"FF",
		417911 => x"FF",
		417912 => x"FF",
		417913 => x"FF",
		417914 => x"FF",
		418035 => x"FF",
		418036 => x"FF",
		418037 => x"FF",
		418038 => x"FF",
		418039 => x"FF",
		418160 => x"FF",
		418161 => x"FF",
		418162 => x"FF",
		418163 => x"FF",
		418164 => x"FF",
		418285 => x"FF",
		418286 => x"FF",
		418287 => x"FF",
		418288 => x"FF",
		418289 => x"FF",
		418934 => x"FF",
		418935 => x"FF",
		418936 => x"FF",
		418937 => x"FF",
		418938 => x"FF",
		419059 => x"FF",
		419060 => x"FF",
		419061 => x"FF",
		419062 => x"FF",
		419063 => x"FF",
		419184 => x"FF",
		419185 => x"FF",
		419186 => x"FF",
		419187 => x"FF",
		419188 => x"FF",
		419309 => x"FF",
		419310 => x"FF",
		419311 => x"FF",
		419312 => x"FF",
		419313 => x"FF",
		419958 => x"FF",
		419959 => x"FF",
		419960 => x"FF",
		419961 => x"FF",
		419962 => x"FF",
		420083 => x"FF",
		420084 => x"FF",
		420085 => x"FF",
		420086 => x"FF",
		420087 => x"FF",
		420208 => x"FF",
		420209 => x"FF",
		420210 => x"FF",
		420211 => x"FF",
		420212 => x"FF",
		420333 => x"FF",
		420334 => x"FF",
		420335 => x"FF",
		420336 => x"FF",
		420337 => x"FF",
		420982 => x"FF",
		420983 => x"FF",
		420984 => x"FF",
		420985 => x"FF",
		420986 => x"FF",
		421107 => x"FF",
		421108 => x"FF",
		421109 => x"FF",
		421110 => x"FF",
		421111 => x"FF",
		421232 => x"FF",
		421233 => x"FF",
		421234 => x"FF",
		421235 => x"FF",
		421236 => x"FF",
		421357 => x"FF",
		421358 => x"FF",
		421359 => x"FF",
		421360 => x"FF",
		421361 => x"FF",
		422006 => x"FF",
		422007 => x"FF",
		422008 => x"FF",
		422009 => x"FF",
		422010 => x"FF",
		422131 => x"FF",
		422132 => x"FF",
		422133 => x"FF",
		422134 => x"FF",
		422135 => x"FF",
		422256 => x"FF",
		422257 => x"FF",
		422258 => x"FF",
		422259 => x"FF",
		422260 => x"FF",
		422381 => x"FF",
		422382 => x"FF",
		422383 => x"FF",
		422384 => x"FF",
		422385 => x"FF",
		423030 => x"FF",
		423031 => x"FF",
		423032 => x"FF",
		423033 => x"FF",
		423034 => x"FF",
		423155 => x"FF",
		423156 => x"FF",
		423157 => x"FF",
		423158 => x"FF",
		423159 => x"FF",
		423280 => x"FF",
		423281 => x"FF",
		423282 => x"FF",
		423283 => x"FF",
		423284 => x"FF",
		423405 => x"FF",
		423406 => x"FF",
		423407 => x"FF",
		423408 => x"FF",
		423409 => x"FF",
		424054 => x"FF",
		424055 => x"FF",
		424056 => x"FF",
		424057 => x"FF",
		424058 => x"FF",
		424179 => x"FF",
		424180 => x"FF",
		424181 => x"FF",
		424182 => x"FF",
		424183 => x"FF",
		424304 => x"FF",
		424305 => x"FF",
		424306 => x"FF",
		424307 => x"FF",
		424308 => x"FF",
		424429 => x"FF",
		424430 => x"FF",
		424431 => x"FF",
		424432 => x"FF",
		424433 => x"FF",
		425078 => x"FF",
		425079 => x"FF",
		425080 => x"FF",
		425081 => x"FF",
		425082 => x"FF",
		425203 => x"FF",
		425204 => x"FF",
		425205 => x"FF",
		425206 => x"FF",
		425207 => x"FF",
		425328 => x"FF",
		425329 => x"FF",
		425330 => x"FF",
		425331 => x"FF",
		425332 => x"FF",
		425453 => x"FF",
		425454 => x"FF",
		425455 => x"FF",
		425456 => x"FF",
		425457 => x"FF",
		426102 => x"FF",
		426103 => x"FF",
		426104 => x"FF",
		426105 => x"FF",
		426106 => x"FF",
		426227 => x"FF",
		426228 => x"FF",
		426229 => x"FF",
		426230 => x"FF",
		426231 => x"FF",
		426352 => x"FF",
		426353 => x"FF",
		426354 => x"FF",
		426355 => x"FF",
		426356 => x"FF",
		426477 => x"FF",
		426478 => x"FF",
		426479 => x"FF",
		426480 => x"FF",
		426481 => x"FF",
		427126 => x"FF",
		427127 => x"FF",
		427128 => x"FF",
		427129 => x"FF",
		427130 => x"FF",
		427251 => x"FF",
		427252 => x"FF",
		427253 => x"FF",
		427254 => x"FF",
		427255 => x"FF",
		427376 => x"FF",
		427377 => x"FF",
		427378 => x"FF",
		427379 => x"FF",
		427380 => x"FF",
		427501 => x"FF",
		427502 => x"FF",
		427503 => x"FF",
		427504 => x"FF",
		427505 => x"FF",
		428150 => x"FF",
		428151 => x"FF",
		428152 => x"FF",
		428153 => x"FF",
		428154 => x"FF",
		428275 => x"FF",
		428276 => x"FF",
		428277 => x"FF",
		428278 => x"FF",
		428279 => x"FF",
		428400 => x"FF",
		428401 => x"FF",
		428402 => x"FF",
		428403 => x"FF",
		428404 => x"FF",
		428525 => x"FF",
		428526 => x"FF",
		428527 => x"FF",
		428528 => x"FF",
		428529 => x"FF",
		429174 => x"FF",
		429175 => x"FF",
		429176 => x"FF",
		429177 => x"FF",
		429178 => x"FF",
		429299 => x"FF",
		429300 => x"FF",
		429301 => x"FF",
		429302 => x"FF",
		429303 => x"FF",
		429424 => x"FF",
		429425 => x"FF",
		429426 => x"FF",
		429427 => x"FF",
		429428 => x"FF",
		429549 => x"FF",
		429550 => x"FF",
		429551 => x"FF",
		429552 => x"FF",
		429553 => x"FF",
		430198 => x"FF",
		430199 => x"FF",
		430200 => x"FF",
		430201 => x"FF",
		430202 => x"FF",
		430323 => x"FF",
		430324 => x"FF",
		430325 => x"FF",
		430326 => x"FF",
		430327 => x"FF",
		430448 => x"FF",
		430449 => x"FF",
		430450 => x"FF",
		430451 => x"FF",
		430452 => x"FF",
		430573 => x"FF",
		430574 => x"FF",
		430575 => x"FF",
		430576 => x"FF",
		430577 => x"FF",
		431222 => x"FF",
		431223 => x"FF",
		431224 => x"FF",
		431225 => x"FF",
		431226 => x"FF",
		431347 => x"FF",
		431348 => x"FF",
		431349 => x"FF",
		431350 => x"FF",
		431351 => x"FF",
		431472 => x"FF",
		431473 => x"FF",
		431474 => x"FF",
		431475 => x"FF",
		431476 => x"FF",
		431597 => x"FF",
		431598 => x"FF",
		431599 => x"FF",
		431600 => x"FF",
		431601 => x"FF",
		432246 => x"FF",
		432247 => x"FF",
		432248 => x"FF",
		432249 => x"FF",
		432250 => x"FF",
		432371 => x"FF",
		432372 => x"FF",
		432373 => x"FF",
		432374 => x"FF",
		432375 => x"FF",
		432496 => x"FF",
		432497 => x"FF",
		432498 => x"FF",
		432499 => x"FF",
		432500 => x"FF",
		432621 => x"FF",
		432622 => x"FF",
		432623 => x"FF",
		432624 => x"FF",
		432625 => x"FF",
		433270 => x"FF",
		433271 => x"FF",
		433272 => x"FF",
		433273 => x"FF",
		433274 => x"FF",
		433275 => x"FF",
		433276 => x"FF",
		433277 => x"FF",
		433278 => x"FF",
		433279 => x"FF",
		433280 => x"FF",
		433281 => x"FF",
		433282 => x"FF",
		433283 => x"FF",
		433284 => x"FF",
		433285 => x"FF",
		433286 => x"FF",
		433287 => x"FF",
		433288 => x"FF",
		433289 => x"FF",
		433290 => x"FF",
		433291 => x"FF",
		433292 => x"FF",
		433293 => x"FF",
		433294 => x"FF",
		433295 => x"FF",
		433296 => x"FF",
		433297 => x"FF",
		433298 => x"FF",
		433299 => x"FF",
		433300 => x"FF",
		433301 => x"FF",
		433302 => x"FF",
		433303 => x"FF",
		433304 => x"FF",
		433305 => x"FF",
		433306 => x"FF",
		433307 => x"FF",
		433308 => x"FF",
		433309 => x"FF",
		433310 => x"FF",
		433311 => x"FF",
		433312 => x"FF",
		433313 => x"FF",
		433314 => x"FF",
		433315 => x"FF",
		433316 => x"FF",
		433317 => x"FF",
		433318 => x"FF",
		433319 => x"FF",
		433320 => x"FF",
		433321 => x"FF",
		433322 => x"FF",
		433323 => x"FF",
		433324 => x"FF",
		433325 => x"FF",
		433326 => x"FF",
		433327 => x"FF",
		433328 => x"FF",
		433329 => x"FF",
		433330 => x"FF",
		433331 => x"FF",
		433332 => x"FF",
		433333 => x"FF",
		433334 => x"FF",
		433335 => x"FF",
		433336 => x"FF",
		433337 => x"FF",
		433338 => x"FF",
		433339 => x"FF",
		433340 => x"FF",
		433341 => x"FF",
		433342 => x"FF",
		433343 => x"FF",
		433344 => x"FF",
		433345 => x"FF",
		433346 => x"FF",
		433347 => x"FF",
		433348 => x"FF",
		433349 => x"FF",
		433350 => x"FF",
		433351 => x"FF",
		433352 => x"FF",
		433353 => x"FF",
		433354 => x"FF",
		433355 => x"FF",
		433356 => x"FF",
		433357 => x"FF",
		433358 => x"FF",
		433359 => x"FF",
		433360 => x"FF",
		433361 => x"FF",
		433362 => x"FF",
		433363 => x"FF",
		433364 => x"FF",
		433365 => x"FF",
		433366 => x"FF",
		433367 => x"FF",
		433368 => x"FF",
		433369 => x"FF",
		433370 => x"FF",
		433371 => x"FF",
		433372 => x"FF",
		433373 => x"FF",
		433374 => x"FF",
		433375 => x"FF",
		433376 => x"FF",
		433377 => x"FF",
		433378 => x"FF",
		433379 => x"FF",
		433380 => x"FF",
		433381 => x"FF",
		433382 => x"FF",
		433383 => x"FF",
		433384 => x"FF",
		433385 => x"FF",
		433386 => x"FF",
		433387 => x"FF",
		433388 => x"FF",
		433389 => x"FF",
		433390 => x"FF",
		433391 => x"FF",
		433392 => x"FF",
		433393 => x"FF",
		433394 => x"FF",
		433395 => x"FF",
		433396 => x"FF",
		433397 => x"FF",
		433398 => x"FF",
		433399 => x"FF",
		433400 => x"FF",
		433401 => x"FF",
		433402 => x"FF",
		433403 => x"FF",
		433404 => x"FF",
		433405 => x"FF",
		433406 => x"FF",
		433407 => x"FF",
		433408 => x"FF",
		433409 => x"FF",
		433410 => x"FF",
		433411 => x"FF",
		433412 => x"FF",
		433413 => x"FF",
		433414 => x"FF",
		433415 => x"FF",
		433416 => x"FF",
		433417 => x"FF",
		433418 => x"FF",
		433419 => x"FF",
		433420 => x"FF",
		433421 => x"FF",
		433422 => x"FF",
		433423 => x"FF",
		433424 => x"FF",
		433425 => x"FF",
		433426 => x"FF",
		433427 => x"FF",
		433428 => x"FF",
		433429 => x"FF",
		433430 => x"FF",
		433431 => x"FF",
		433432 => x"FF",
		433433 => x"FF",
		433434 => x"FF",
		433435 => x"FF",
		433436 => x"FF",
		433437 => x"FF",
		433438 => x"FF",
		433439 => x"FF",
		433440 => x"FF",
		433441 => x"FF",
		433442 => x"FF",
		433443 => x"FF",
		433444 => x"FF",
		433445 => x"FF",
		433446 => x"FF",
		433447 => x"FF",
		433448 => x"FF",
		433449 => x"FF",
		433450 => x"FF",
		433451 => x"FF",
		433452 => x"FF",
		433453 => x"FF",
		433454 => x"FF",
		433455 => x"FF",
		433456 => x"FF",
		433457 => x"FF",
		433458 => x"FF",
		433459 => x"FF",
		433460 => x"FF",
		433461 => x"FF",
		433462 => x"FF",
		433463 => x"FF",
		433464 => x"FF",
		433465 => x"FF",
		433466 => x"FF",
		433467 => x"FF",
		433468 => x"FF",
		433469 => x"FF",
		433470 => x"FF",
		433471 => x"FF",
		433472 => x"FF",
		433473 => x"FF",
		433474 => x"FF",
		433475 => x"FF",
		433476 => x"FF",
		433477 => x"FF",
		433478 => x"FF",
		433479 => x"FF",
		433480 => x"FF",
		433481 => x"FF",
		433482 => x"FF",
		433483 => x"FF",
		433484 => x"FF",
		433485 => x"FF",
		433486 => x"FF",
		433487 => x"FF",
		433488 => x"FF",
		433489 => x"FF",
		433490 => x"FF",
		433491 => x"FF",
		433492 => x"FF",
		433493 => x"FF",
		433494 => x"FF",
		433495 => x"FF",
		433496 => x"FF",
		433497 => x"FF",
		433498 => x"FF",
		433499 => x"FF",
		433500 => x"FF",
		433501 => x"FF",
		433502 => x"FF",
		433503 => x"FF",
		433504 => x"FF",
		433505 => x"FF",
		433506 => x"FF",
		433507 => x"FF",
		433508 => x"FF",
		433509 => x"FF",
		433510 => x"FF",
		433511 => x"FF",
		433512 => x"FF",
		433513 => x"FF",
		433514 => x"FF",
		433515 => x"FF",
		433516 => x"FF",
		433517 => x"FF",
		433518 => x"FF",
		433519 => x"FF",
		433520 => x"FF",
		433521 => x"FF",
		433522 => x"FF",
		433523 => x"FF",
		433524 => x"FF",
		433525 => x"FF",
		433526 => x"FF",
		433527 => x"FF",
		433528 => x"FF",
		433529 => x"FF",
		433530 => x"FF",
		433531 => x"FF",
		433532 => x"FF",
		433533 => x"FF",
		433534 => x"FF",
		433535 => x"FF",
		433536 => x"FF",
		433537 => x"FF",
		433538 => x"FF",
		433539 => x"FF",
		433540 => x"FF",
		433541 => x"FF",
		433542 => x"FF",
		433543 => x"FF",
		433544 => x"FF",
		433545 => x"FF",
		433546 => x"FF",
		433547 => x"FF",
		433548 => x"FF",
		433549 => x"FF",
		433550 => x"FF",
		433551 => x"FF",
		433552 => x"FF",
		433553 => x"FF",
		433554 => x"FF",
		433555 => x"FF",
		433556 => x"FF",
		433557 => x"FF",
		433558 => x"FF",
		433559 => x"FF",
		433560 => x"FF",
		433561 => x"FF",
		433562 => x"FF",
		433563 => x"FF",
		433564 => x"FF",
		433565 => x"FF",
		433566 => x"FF",
		433567 => x"FF",
		433568 => x"FF",
		433569 => x"FF",
		433570 => x"FF",
		433571 => x"FF",
		433572 => x"FF",
		433573 => x"FF",
		433574 => x"FF",
		433575 => x"FF",
		433576 => x"FF",
		433577 => x"FF",
		433578 => x"FF",
		433579 => x"FF",
		433580 => x"FF",
		433581 => x"FF",
		433582 => x"FF",
		433583 => x"FF",
		433584 => x"FF",
		433585 => x"FF",
		433586 => x"FF",
		433587 => x"FF",
		433588 => x"FF",
		433589 => x"FF",
		433590 => x"FF",
		433591 => x"FF",
		433592 => x"FF",
		433593 => x"FF",
		433594 => x"FF",
		433595 => x"FF",
		433596 => x"FF",
		433597 => x"FF",
		433598 => x"FF",
		433599 => x"FF",
		433600 => x"FF",
		433601 => x"FF",
		433602 => x"FF",
		433603 => x"FF",
		433604 => x"FF",
		433605 => x"FF",
		433606 => x"FF",
		433607 => x"FF",
		433608 => x"FF",
		433609 => x"FF",
		433610 => x"FF",
		433611 => x"FF",
		433612 => x"FF",
		433613 => x"FF",
		433614 => x"FF",
		433615 => x"FF",
		433616 => x"FF",
		433617 => x"FF",
		433618 => x"FF",
		433619 => x"FF",
		433620 => x"FF",
		433621 => x"FF",
		433622 => x"FF",
		433623 => x"FF",
		433624 => x"FF",
		433625 => x"FF",
		433626 => x"FF",
		433627 => x"FF",
		433628 => x"FF",
		433629 => x"FF",
		433630 => x"FF",
		433631 => x"FF",
		433632 => x"FF",
		433633 => x"FF",
		433634 => x"FF",
		433635 => x"FF",
		433636 => x"FF",
		433637 => x"FF",
		433638 => x"FF",
		433639 => x"FF",
		433640 => x"FF",
		433641 => x"FF",
		433642 => x"FF",
		433643 => x"FF",
		433644 => x"FF",
		433645 => x"FF",
		433646 => x"FF",
		433647 => x"FF",
		433648 => x"FF",
		433649 => x"FF",
		434294 => x"FF",
		434295 => x"FF",
		434296 => x"FF",
		434297 => x"FF",
		434298 => x"FF",
		434299 => x"FF",
		434300 => x"FF",
		434301 => x"FF",
		434302 => x"FF",
		434303 => x"FF",
		434304 => x"FF",
		434305 => x"FF",
		434306 => x"FF",
		434307 => x"FF",
		434308 => x"FF",
		434309 => x"FF",
		434310 => x"FF",
		434311 => x"FF",
		434312 => x"FF",
		434313 => x"FF",
		434314 => x"FF",
		434315 => x"FF",
		434316 => x"FF",
		434317 => x"FF",
		434318 => x"FF",
		434319 => x"FF",
		434320 => x"FF",
		434321 => x"FF",
		434322 => x"FF",
		434323 => x"FF",
		434324 => x"FF",
		434325 => x"FF",
		434326 => x"FF",
		434327 => x"FF",
		434328 => x"FF",
		434329 => x"FF",
		434330 => x"FF",
		434331 => x"FF",
		434332 => x"FF",
		434333 => x"FF",
		434334 => x"FF",
		434335 => x"FF",
		434336 => x"FF",
		434337 => x"FF",
		434338 => x"FF",
		434339 => x"FF",
		434340 => x"FF",
		434341 => x"FF",
		434342 => x"FF",
		434343 => x"FF",
		434344 => x"FF",
		434345 => x"FF",
		434346 => x"FF",
		434347 => x"FF",
		434348 => x"FF",
		434349 => x"FF",
		434350 => x"FF",
		434351 => x"FF",
		434352 => x"FF",
		434353 => x"FF",
		434354 => x"FF",
		434355 => x"FF",
		434356 => x"FF",
		434357 => x"FF",
		434358 => x"FF",
		434359 => x"FF",
		434360 => x"FF",
		434361 => x"FF",
		434362 => x"FF",
		434363 => x"FF",
		434364 => x"FF",
		434365 => x"FF",
		434366 => x"FF",
		434367 => x"FF",
		434368 => x"FF",
		434369 => x"FF",
		434370 => x"FF",
		434371 => x"FF",
		434372 => x"FF",
		434373 => x"FF",
		434374 => x"FF",
		434375 => x"FF",
		434376 => x"FF",
		434377 => x"FF",
		434378 => x"FF",
		434379 => x"FF",
		434380 => x"FF",
		434381 => x"FF",
		434382 => x"FF",
		434383 => x"FF",
		434384 => x"FF",
		434385 => x"FF",
		434386 => x"FF",
		434387 => x"FF",
		434388 => x"FF",
		434389 => x"FF",
		434390 => x"FF",
		434391 => x"FF",
		434392 => x"FF",
		434393 => x"FF",
		434394 => x"FF",
		434395 => x"FF",
		434396 => x"FF",
		434397 => x"FF",
		434398 => x"FF",
		434399 => x"FF",
		434400 => x"FF",
		434401 => x"FF",
		434402 => x"FF",
		434403 => x"FF",
		434404 => x"FF",
		434405 => x"FF",
		434406 => x"FF",
		434407 => x"FF",
		434408 => x"FF",
		434409 => x"FF",
		434410 => x"FF",
		434411 => x"FF",
		434412 => x"FF",
		434413 => x"FF",
		434414 => x"FF",
		434415 => x"FF",
		434416 => x"FF",
		434417 => x"FF",
		434418 => x"FF",
		434419 => x"FF",
		434420 => x"FF",
		434421 => x"FF",
		434422 => x"FF",
		434423 => x"FF",
		434424 => x"FF",
		434425 => x"FF",
		434426 => x"FF",
		434427 => x"FF",
		434428 => x"FF",
		434429 => x"FF",
		434430 => x"FF",
		434431 => x"FF",
		434432 => x"FF",
		434433 => x"FF",
		434434 => x"FF",
		434435 => x"FF",
		434436 => x"FF",
		434437 => x"FF",
		434438 => x"FF",
		434439 => x"FF",
		434440 => x"FF",
		434441 => x"FF",
		434442 => x"FF",
		434443 => x"FF",
		434444 => x"FF",
		434445 => x"FF",
		434446 => x"FF",
		434447 => x"FF",
		434448 => x"FF",
		434449 => x"FF",
		434450 => x"FF",
		434451 => x"FF",
		434452 => x"FF",
		434453 => x"FF",
		434454 => x"FF",
		434455 => x"FF",
		434456 => x"FF",
		434457 => x"FF",
		434458 => x"FF",
		434459 => x"FF",
		434460 => x"FF",
		434461 => x"FF",
		434462 => x"FF",
		434463 => x"FF",
		434464 => x"FF",
		434465 => x"FF",
		434466 => x"FF",
		434467 => x"FF",
		434468 => x"FF",
		434469 => x"FF",
		434470 => x"FF",
		434471 => x"FF",
		434472 => x"FF",
		434473 => x"FF",
		434474 => x"FF",
		434475 => x"FF",
		434476 => x"FF",
		434477 => x"FF",
		434478 => x"FF",
		434479 => x"FF",
		434480 => x"FF",
		434481 => x"FF",
		434482 => x"FF",
		434483 => x"FF",
		434484 => x"FF",
		434485 => x"FF",
		434486 => x"FF",
		434487 => x"FF",
		434488 => x"FF",
		434489 => x"FF",
		434490 => x"FF",
		434491 => x"FF",
		434492 => x"FF",
		434493 => x"FF",
		434494 => x"FF",
		434495 => x"FF",
		434496 => x"FF",
		434497 => x"FF",
		434498 => x"FF",
		434499 => x"FF",
		434500 => x"FF",
		434501 => x"FF",
		434502 => x"FF",
		434503 => x"FF",
		434504 => x"FF",
		434505 => x"FF",
		434506 => x"FF",
		434507 => x"FF",
		434508 => x"FF",
		434509 => x"FF",
		434510 => x"FF",
		434511 => x"FF",
		434512 => x"FF",
		434513 => x"FF",
		434514 => x"FF",
		434515 => x"FF",
		434516 => x"FF",
		434517 => x"FF",
		434518 => x"FF",
		434519 => x"FF",
		434520 => x"FF",
		434521 => x"FF",
		434522 => x"FF",
		434523 => x"FF",
		434524 => x"FF",
		434525 => x"FF",
		434526 => x"FF",
		434527 => x"FF",
		434528 => x"FF",
		434529 => x"FF",
		434530 => x"FF",
		434531 => x"FF",
		434532 => x"FF",
		434533 => x"FF",
		434534 => x"FF",
		434535 => x"FF",
		434536 => x"FF",
		434537 => x"FF",
		434538 => x"FF",
		434539 => x"FF",
		434540 => x"FF",
		434541 => x"FF",
		434542 => x"FF",
		434543 => x"FF",
		434544 => x"FF",
		434545 => x"FF",
		434546 => x"FF",
		434547 => x"FF",
		434548 => x"FF",
		434549 => x"FF",
		434550 => x"FF",
		434551 => x"FF",
		434552 => x"FF",
		434553 => x"FF",
		434554 => x"FF",
		434555 => x"FF",
		434556 => x"FF",
		434557 => x"FF",
		434558 => x"FF",
		434559 => x"FF",
		434560 => x"FF",
		434561 => x"FF",
		434562 => x"FF",
		434563 => x"FF",
		434564 => x"FF",
		434565 => x"FF",
		434566 => x"FF",
		434567 => x"FF",
		434568 => x"FF",
		434569 => x"FF",
		434570 => x"FF",
		434571 => x"FF",
		434572 => x"FF",
		434573 => x"FF",
		434574 => x"FF",
		434575 => x"FF",
		434576 => x"FF",
		434577 => x"FF",
		434578 => x"FF",
		434579 => x"FF",
		434580 => x"FF",
		434581 => x"FF",
		434582 => x"FF",
		434583 => x"FF",
		434584 => x"FF",
		434585 => x"FF",
		434586 => x"FF",
		434587 => x"FF",
		434588 => x"FF",
		434589 => x"FF",
		434590 => x"FF",
		434591 => x"FF",
		434592 => x"FF",
		434593 => x"FF",
		434594 => x"FF",
		434595 => x"FF",
		434596 => x"FF",
		434597 => x"FF",
		434598 => x"FF",
		434599 => x"FF",
		434600 => x"FF",
		434601 => x"FF",
		434602 => x"FF",
		434603 => x"FF",
		434604 => x"FF",
		434605 => x"FF",
		434606 => x"FF",
		434607 => x"FF",
		434608 => x"FF",
		434609 => x"FF",
		434610 => x"FF",
		434611 => x"FF",
		434612 => x"FF",
		434613 => x"FF",
		434614 => x"FF",
		434615 => x"FF",
		434616 => x"FF",
		434617 => x"FF",
		434618 => x"FF",
		434619 => x"FF",
		434620 => x"FF",
		434621 => x"FF",
		434622 => x"FF",
		434623 => x"FF",
		434624 => x"FF",
		434625 => x"FF",
		434626 => x"FF",
		434627 => x"FF",
		434628 => x"FF",
		434629 => x"FF",
		434630 => x"FF",
		434631 => x"FF",
		434632 => x"FF",
		434633 => x"FF",
		434634 => x"FF",
		434635 => x"FF",
		434636 => x"FF",
		434637 => x"FF",
		434638 => x"FF",
		434639 => x"FF",
		434640 => x"FF",
		434641 => x"FF",
		434642 => x"FF",
		434643 => x"FF",
		434644 => x"FF",
		434645 => x"FF",
		434646 => x"FF",
		434647 => x"FF",
		434648 => x"FF",
		434649 => x"FF",
		434650 => x"FF",
		434651 => x"FF",
		434652 => x"FF",
		434653 => x"FF",
		434654 => x"FF",
		434655 => x"FF",
		434656 => x"FF",
		434657 => x"FF",
		434658 => x"FF",
		434659 => x"FF",
		434660 => x"FF",
		434661 => x"FF",
		434662 => x"FF",
		434663 => x"FF",
		434664 => x"FF",
		434665 => x"FF",
		434666 => x"FF",
		434667 => x"FF",
		434668 => x"FF",
		434669 => x"FF",
		434670 => x"FF",
		434671 => x"FF",
		434672 => x"FF",
		434673 => x"FF",
		435318 => x"FF",
		435319 => x"FF",
		435320 => x"FF",
		435321 => x"FF",
		435322 => x"FF",
		435323 => x"FF",
		435324 => x"FF",
		435325 => x"FF",
		435326 => x"FF",
		435327 => x"FF",
		435328 => x"FF",
		435329 => x"FF",
		435330 => x"FF",
		435331 => x"FF",
		435332 => x"FF",
		435333 => x"FF",
		435334 => x"FF",
		435335 => x"FF",
		435336 => x"FF",
		435337 => x"FF",
		435338 => x"FF",
		435339 => x"FF",
		435340 => x"FF",
		435341 => x"FF",
		435342 => x"FF",
		435343 => x"FF",
		435344 => x"FF",
		435345 => x"FF",
		435346 => x"FF",
		435347 => x"FF",
		435348 => x"FF",
		435349 => x"FF",
		435350 => x"FF",
		435351 => x"FF",
		435352 => x"FF",
		435353 => x"FF",
		435354 => x"FF",
		435355 => x"FF",
		435356 => x"FF",
		435357 => x"FF",
		435358 => x"FF",
		435359 => x"FF",
		435360 => x"FF",
		435361 => x"FF",
		435362 => x"FF",
		435363 => x"FF",
		435364 => x"FF",
		435365 => x"FF",
		435366 => x"FF",
		435367 => x"FF",
		435368 => x"FF",
		435369 => x"FF",
		435370 => x"FF",
		435371 => x"FF",
		435372 => x"FF",
		435373 => x"FF",
		435374 => x"FF",
		435375 => x"FF",
		435376 => x"FF",
		435377 => x"FF",
		435378 => x"FF",
		435379 => x"FF",
		435380 => x"FF",
		435381 => x"FF",
		435382 => x"FF",
		435383 => x"FF",
		435384 => x"FF",
		435385 => x"FF",
		435386 => x"FF",
		435387 => x"FF",
		435388 => x"FF",
		435389 => x"FF",
		435390 => x"FF",
		435391 => x"FF",
		435392 => x"FF",
		435393 => x"FF",
		435394 => x"FF",
		435395 => x"FF",
		435396 => x"FF",
		435397 => x"FF",
		435398 => x"FF",
		435399 => x"FF",
		435400 => x"FF",
		435401 => x"FF",
		435402 => x"FF",
		435403 => x"FF",
		435404 => x"FF",
		435405 => x"FF",
		435406 => x"FF",
		435407 => x"FF",
		435408 => x"FF",
		435409 => x"FF",
		435410 => x"FF",
		435411 => x"FF",
		435412 => x"FF",
		435413 => x"FF",
		435414 => x"FF",
		435415 => x"FF",
		435416 => x"FF",
		435417 => x"FF",
		435418 => x"FF",
		435419 => x"FF",
		435420 => x"FF",
		435421 => x"FF",
		435422 => x"FF",
		435423 => x"FF",
		435424 => x"FF",
		435425 => x"FF",
		435426 => x"FF",
		435427 => x"FF",
		435428 => x"FF",
		435429 => x"FF",
		435430 => x"FF",
		435431 => x"FF",
		435432 => x"FF",
		435433 => x"FF",
		435434 => x"FF",
		435435 => x"FF",
		435436 => x"FF",
		435437 => x"FF",
		435438 => x"FF",
		435439 => x"FF",
		435440 => x"FF",
		435441 => x"FF",
		435442 => x"FF",
		435443 => x"FF",
		435444 => x"FF",
		435445 => x"FF",
		435446 => x"FF",
		435447 => x"FF",
		435448 => x"FF",
		435449 => x"FF",
		435450 => x"FF",
		435451 => x"FF",
		435452 => x"FF",
		435453 => x"FF",
		435454 => x"FF",
		435455 => x"FF",
		435456 => x"FF",
		435457 => x"FF",
		435458 => x"FF",
		435459 => x"FF",
		435460 => x"FF",
		435461 => x"FF",
		435462 => x"FF",
		435463 => x"FF",
		435464 => x"FF",
		435465 => x"FF",
		435466 => x"FF",
		435467 => x"FF",
		435468 => x"FF",
		435469 => x"FF",
		435470 => x"FF",
		435471 => x"FF",
		435472 => x"FF",
		435473 => x"FF",
		435474 => x"FF",
		435475 => x"FF",
		435476 => x"FF",
		435477 => x"FF",
		435478 => x"FF",
		435479 => x"FF",
		435480 => x"FF",
		435481 => x"FF",
		435482 => x"FF",
		435483 => x"FF",
		435484 => x"FF",
		435485 => x"FF",
		435486 => x"FF",
		435487 => x"FF",
		435488 => x"FF",
		435489 => x"FF",
		435490 => x"FF",
		435491 => x"FF",
		435492 => x"FF",
		435493 => x"FF",
		435494 => x"FF",
		435495 => x"FF",
		435496 => x"FF",
		435497 => x"FF",
		435498 => x"FF",
		435499 => x"FF",
		435500 => x"FF",
		435501 => x"FF",
		435502 => x"FF",
		435503 => x"FF",
		435504 => x"FF",
		435505 => x"FF",
		435506 => x"FF",
		435507 => x"FF",
		435508 => x"FF",
		435509 => x"FF",
		435510 => x"FF",
		435511 => x"FF",
		435512 => x"FF",
		435513 => x"FF",
		435514 => x"FF",
		435515 => x"FF",
		435516 => x"FF",
		435517 => x"FF",
		435518 => x"FF",
		435519 => x"FF",
		435520 => x"FF",
		435521 => x"FF",
		435522 => x"FF",
		435523 => x"FF",
		435524 => x"FF",
		435525 => x"FF",
		435526 => x"FF",
		435527 => x"FF",
		435528 => x"FF",
		435529 => x"FF",
		435530 => x"FF",
		435531 => x"FF",
		435532 => x"FF",
		435533 => x"FF",
		435534 => x"FF",
		435535 => x"FF",
		435536 => x"FF",
		435537 => x"FF",
		435538 => x"FF",
		435539 => x"FF",
		435540 => x"FF",
		435541 => x"FF",
		435542 => x"FF",
		435543 => x"FF",
		435544 => x"FF",
		435545 => x"FF",
		435546 => x"FF",
		435547 => x"FF",
		435548 => x"FF",
		435549 => x"FF",
		435550 => x"FF",
		435551 => x"FF",
		435552 => x"FF",
		435553 => x"FF",
		435554 => x"FF",
		435555 => x"FF",
		435556 => x"FF",
		435557 => x"FF",
		435558 => x"FF",
		435559 => x"FF",
		435560 => x"FF",
		435561 => x"FF",
		435562 => x"FF",
		435563 => x"FF",
		435564 => x"FF",
		435565 => x"FF",
		435566 => x"FF",
		435567 => x"FF",
		435568 => x"FF",
		435569 => x"FF",
		435570 => x"FF",
		435571 => x"FF",
		435572 => x"FF",
		435573 => x"FF",
		435574 => x"FF",
		435575 => x"FF",
		435576 => x"FF",
		435577 => x"FF",
		435578 => x"FF",
		435579 => x"FF",
		435580 => x"FF",
		435581 => x"FF",
		435582 => x"FF",
		435583 => x"FF",
		435584 => x"FF",
		435585 => x"FF",
		435586 => x"FF",
		435587 => x"FF",
		435588 => x"FF",
		435589 => x"FF",
		435590 => x"FF",
		435591 => x"FF",
		435592 => x"FF",
		435593 => x"FF",
		435594 => x"FF",
		435595 => x"FF",
		435596 => x"FF",
		435597 => x"FF",
		435598 => x"FF",
		435599 => x"FF",
		435600 => x"FF",
		435601 => x"FF",
		435602 => x"FF",
		435603 => x"FF",
		435604 => x"FF",
		435605 => x"FF",
		435606 => x"FF",
		435607 => x"FF",
		435608 => x"FF",
		435609 => x"FF",
		435610 => x"FF",
		435611 => x"FF",
		435612 => x"FF",
		435613 => x"FF",
		435614 => x"FF",
		435615 => x"FF",
		435616 => x"FF",
		435617 => x"FF",
		435618 => x"FF",
		435619 => x"FF",
		435620 => x"FF",
		435621 => x"FF",
		435622 => x"FF",
		435623 => x"FF",
		435624 => x"FF",
		435625 => x"FF",
		435626 => x"FF",
		435627 => x"FF",
		435628 => x"FF",
		435629 => x"FF",
		435630 => x"FF",
		435631 => x"FF",
		435632 => x"FF",
		435633 => x"FF",
		435634 => x"FF",
		435635 => x"FF",
		435636 => x"FF",
		435637 => x"FF",
		435638 => x"FF",
		435639 => x"FF",
		435640 => x"FF",
		435641 => x"FF",
		435642 => x"FF",
		435643 => x"FF",
		435644 => x"FF",
		435645 => x"FF",
		435646 => x"FF",
		435647 => x"FF",
		435648 => x"FF",
		435649 => x"FF",
		435650 => x"FF",
		435651 => x"FF",
		435652 => x"FF",
		435653 => x"FF",
		435654 => x"FF",
		435655 => x"FF",
		435656 => x"FF",
		435657 => x"FF",
		435658 => x"FF",
		435659 => x"FF",
		435660 => x"FF",
		435661 => x"FF",
		435662 => x"FF",
		435663 => x"FF",
		435664 => x"FF",
		435665 => x"FF",
		435666 => x"FF",
		435667 => x"FF",
		435668 => x"FF",
		435669 => x"FF",
		435670 => x"FF",
		435671 => x"FF",
		435672 => x"FF",
		435673 => x"FF",
		435674 => x"FF",
		435675 => x"FF",
		435676 => x"FF",
		435677 => x"FF",
		435678 => x"FF",
		435679 => x"FF",
		435680 => x"FF",
		435681 => x"FF",
		435682 => x"FF",
		435683 => x"FF",
		435684 => x"FF",
		435685 => x"FF",
		435686 => x"FF",
		435687 => x"FF",
		435688 => x"FF",
		435689 => x"FF",
		435690 => x"FF",
		435691 => x"FF",
		435692 => x"FF",
		435693 => x"FF",
		435694 => x"FF",
		435695 => x"FF",
		435696 => x"FF",
		435697 => x"FF",
		436342 => x"FF",
		436343 => x"FF",
		436344 => x"FF",
		436345 => x"FF",
		436346 => x"FF",
		436347 => x"FF",
		436348 => x"FF",
		436349 => x"FF",
		436350 => x"FF",
		436351 => x"FF",
		436352 => x"FF",
		436353 => x"FF",
		436354 => x"FF",
		436355 => x"FF",
		436356 => x"FF",
		436357 => x"FF",
		436358 => x"FF",
		436359 => x"FF",
		436360 => x"FF",
		436361 => x"FF",
		436362 => x"FF",
		436363 => x"FF",
		436364 => x"FF",
		436365 => x"FF",
		436366 => x"FF",
		436367 => x"FF",
		436368 => x"FF",
		436369 => x"FF",
		436370 => x"FF",
		436371 => x"FF",
		436372 => x"FF",
		436373 => x"FF",
		436374 => x"FF",
		436375 => x"FF",
		436376 => x"FF",
		436377 => x"FF",
		436378 => x"FF",
		436379 => x"FF",
		436380 => x"FF",
		436381 => x"FF",
		436382 => x"FF",
		436383 => x"FF",
		436384 => x"FF",
		436385 => x"FF",
		436386 => x"FF",
		436387 => x"FF",
		436388 => x"FF",
		436389 => x"FF",
		436390 => x"FF",
		436391 => x"FF",
		436392 => x"FF",
		436393 => x"FF",
		436394 => x"FF",
		436395 => x"FF",
		436396 => x"FF",
		436397 => x"FF",
		436398 => x"FF",
		436399 => x"FF",
		436400 => x"FF",
		436401 => x"FF",
		436402 => x"FF",
		436403 => x"FF",
		436404 => x"FF",
		436405 => x"FF",
		436406 => x"FF",
		436407 => x"FF",
		436408 => x"FF",
		436409 => x"FF",
		436410 => x"FF",
		436411 => x"FF",
		436412 => x"FF",
		436413 => x"FF",
		436414 => x"FF",
		436415 => x"FF",
		436416 => x"FF",
		436417 => x"FF",
		436418 => x"FF",
		436419 => x"FF",
		436420 => x"FF",
		436421 => x"FF",
		436422 => x"FF",
		436423 => x"FF",
		436424 => x"FF",
		436425 => x"FF",
		436426 => x"FF",
		436427 => x"FF",
		436428 => x"FF",
		436429 => x"FF",
		436430 => x"FF",
		436431 => x"FF",
		436432 => x"FF",
		436433 => x"FF",
		436434 => x"FF",
		436435 => x"FF",
		436436 => x"FF",
		436437 => x"FF",
		436438 => x"FF",
		436439 => x"FF",
		436440 => x"FF",
		436441 => x"FF",
		436442 => x"FF",
		436443 => x"FF",
		436444 => x"FF",
		436445 => x"FF",
		436446 => x"FF",
		436447 => x"FF",
		436448 => x"FF",
		436449 => x"FF",
		436450 => x"FF",
		436451 => x"FF",
		436452 => x"FF",
		436453 => x"FF",
		436454 => x"FF",
		436455 => x"FF",
		436456 => x"FF",
		436457 => x"FF",
		436458 => x"FF",
		436459 => x"FF",
		436460 => x"FF",
		436461 => x"FF",
		436462 => x"FF",
		436463 => x"FF",
		436464 => x"FF",
		436465 => x"FF",
		436466 => x"FF",
		436467 => x"FF",
		436468 => x"FF",
		436469 => x"FF",
		436470 => x"FF",
		436471 => x"FF",
		436472 => x"FF",
		436473 => x"FF",
		436474 => x"FF",
		436475 => x"FF",
		436476 => x"FF",
		436477 => x"FF",
		436478 => x"FF",
		436479 => x"FF",
		436480 => x"FF",
		436481 => x"FF",
		436482 => x"FF",
		436483 => x"FF",
		436484 => x"FF",
		436485 => x"FF",
		436486 => x"FF",
		436487 => x"FF",
		436488 => x"FF",
		436489 => x"FF",
		436490 => x"FF",
		436491 => x"FF",
		436492 => x"FF",
		436493 => x"FF",
		436494 => x"FF",
		436495 => x"FF",
		436496 => x"FF",
		436497 => x"FF",
		436498 => x"FF",
		436499 => x"FF",
		436500 => x"FF",
		436501 => x"FF",
		436502 => x"FF",
		436503 => x"FF",
		436504 => x"FF",
		436505 => x"FF",
		436506 => x"FF",
		436507 => x"FF",
		436508 => x"FF",
		436509 => x"FF",
		436510 => x"FF",
		436511 => x"FF",
		436512 => x"FF",
		436513 => x"FF",
		436514 => x"FF",
		436515 => x"FF",
		436516 => x"FF",
		436517 => x"FF",
		436518 => x"FF",
		436519 => x"FF",
		436520 => x"FF",
		436521 => x"FF",
		436522 => x"FF",
		436523 => x"FF",
		436524 => x"FF",
		436525 => x"FF",
		436526 => x"FF",
		436527 => x"FF",
		436528 => x"FF",
		436529 => x"FF",
		436530 => x"FF",
		436531 => x"FF",
		436532 => x"FF",
		436533 => x"FF",
		436534 => x"FF",
		436535 => x"FF",
		436536 => x"FF",
		436537 => x"FF",
		436538 => x"FF",
		436539 => x"FF",
		436540 => x"FF",
		436541 => x"FF",
		436542 => x"FF",
		436543 => x"FF",
		436544 => x"FF",
		436545 => x"FF",
		436546 => x"FF",
		436547 => x"FF",
		436548 => x"FF",
		436549 => x"FF",
		436550 => x"FF",
		436551 => x"FF",
		436552 => x"FF",
		436553 => x"FF",
		436554 => x"FF",
		436555 => x"FF",
		436556 => x"FF",
		436557 => x"FF",
		436558 => x"FF",
		436559 => x"FF",
		436560 => x"FF",
		436561 => x"FF",
		436562 => x"FF",
		436563 => x"FF",
		436564 => x"FF",
		436565 => x"FF",
		436566 => x"FF",
		436567 => x"FF",
		436568 => x"FF",
		436569 => x"FF",
		436570 => x"FF",
		436571 => x"FF",
		436572 => x"FF",
		436573 => x"FF",
		436574 => x"FF",
		436575 => x"FF",
		436576 => x"FF",
		436577 => x"FF",
		436578 => x"FF",
		436579 => x"FF",
		436580 => x"FF",
		436581 => x"FF",
		436582 => x"FF",
		436583 => x"FF",
		436584 => x"FF",
		436585 => x"FF",
		436586 => x"FF",
		436587 => x"FF",
		436588 => x"FF",
		436589 => x"FF",
		436590 => x"FF",
		436591 => x"FF",
		436592 => x"FF",
		436593 => x"FF",
		436594 => x"FF",
		436595 => x"FF",
		436596 => x"FF",
		436597 => x"FF",
		436598 => x"FF",
		436599 => x"FF",
		436600 => x"FF",
		436601 => x"FF",
		436602 => x"FF",
		436603 => x"FF",
		436604 => x"FF",
		436605 => x"FF",
		436606 => x"FF",
		436607 => x"FF",
		436608 => x"FF",
		436609 => x"FF",
		436610 => x"FF",
		436611 => x"FF",
		436612 => x"FF",
		436613 => x"FF",
		436614 => x"FF",
		436615 => x"FF",
		436616 => x"FF",
		436617 => x"FF",
		436618 => x"FF",
		436619 => x"FF",
		436620 => x"FF",
		436621 => x"FF",
		436622 => x"FF",
		436623 => x"FF",
		436624 => x"FF",
		436625 => x"FF",
		436626 => x"FF",
		436627 => x"FF",
		436628 => x"FF",
		436629 => x"FF",
		436630 => x"FF",
		436631 => x"FF",
		436632 => x"FF",
		436633 => x"FF",
		436634 => x"FF",
		436635 => x"FF",
		436636 => x"FF",
		436637 => x"FF",
		436638 => x"FF",
		436639 => x"FF",
		436640 => x"FF",
		436641 => x"FF",
		436642 => x"FF",
		436643 => x"FF",
		436644 => x"FF",
		436645 => x"FF",
		436646 => x"FF",
		436647 => x"FF",
		436648 => x"FF",
		436649 => x"FF",
		436650 => x"FF",
		436651 => x"FF",
		436652 => x"FF",
		436653 => x"FF",
		436654 => x"FF",
		436655 => x"FF",
		436656 => x"FF",
		436657 => x"FF",
		436658 => x"FF",
		436659 => x"FF",
		436660 => x"FF",
		436661 => x"FF",
		436662 => x"FF",
		436663 => x"FF",
		436664 => x"FF",
		436665 => x"FF",
		436666 => x"FF",
		436667 => x"FF",
		436668 => x"FF",
		436669 => x"FF",
		436670 => x"FF",
		436671 => x"FF",
		436672 => x"FF",
		436673 => x"FF",
		436674 => x"FF",
		436675 => x"FF",
		436676 => x"FF",
		436677 => x"FF",
		436678 => x"FF",
		436679 => x"FF",
		436680 => x"FF",
		436681 => x"FF",
		436682 => x"FF",
		436683 => x"FF",
		436684 => x"FF",
		436685 => x"FF",
		436686 => x"FF",
		436687 => x"FF",
		436688 => x"FF",
		436689 => x"FF",
		436690 => x"FF",
		436691 => x"FF",
		436692 => x"FF",
		436693 => x"FF",
		436694 => x"FF",
		436695 => x"FF",
		436696 => x"FF",
		436697 => x"FF",
		436698 => x"FF",
		436699 => x"FF",
		436700 => x"FF",
		436701 => x"FF",
		436702 => x"FF",
		436703 => x"FF",
		436704 => x"FF",
		436705 => x"FF",
		436706 => x"FF",
		436707 => x"FF",
		436708 => x"FF",
		436709 => x"FF",
		436710 => x"FF",
		436711 => x"FF",
		436712 => x"FF",
		436713 => x"FF",
		436714 => x"FF",
		436715 => x"FF",
		436716 => x"FF",
		436717 => x"FF",
		436718 => x"FF",
		436719 => x"FF",
		436720 => x"FF",
		436721 => x"FF",
		437366 => x"FF",
		437367 => x"FF",
		437368 => x"FF",
		437369 => x"FF",
		437370 => x"FF",
		437371 => x"FF",
		437372 => x"FF",
		437373 => x"FF",
		437374 => x"FF",
		437375 => x"FF",
		437376 => x"FF",
		437377 => x"FF",
		437378 => x"FF",
		437379 => x"FF",
		437380 => x"FF",
		437381 => x"FF",
		437382 => x"FF",
		437383 => x"FF",
		437384 => x"FF",
		437385 => x"FF",
		437386 => x"FF",
		437387 => x"FF",
		437388 => x"FF",
		437389 => x"FF",
		437390 => x"FF",
		437391 => x"FF",
		437392 => x"FF",
		437393 => x"FF",
		437394 => x"FF",
		437395 => x"FF",
		437396 => x"FF",
		437397 => x"FF",
		437398 => x"FF",
		437399 => x"FF",
		437400 => x"FF",
		437401 => x"FF",
		437402 => x"FF",
		437403 => x"FF",
		437404 => x"FF",
		437405 => x"FF",
		437406 => x"FF",
		437407 => x"FF",
		437408 => x"FF",
		437409 => x"FF",
		437410 => x"FF",
		437411 => x"FF",
		437412 => x"FF",
		437413 => x"FF",
		437414 => x"FF",
		437415 => x"FF",
		437416 => x"FF",
		437417 => x"FF",
		437418 => x"FF",
		437419 => x"FF",
		437420 => x"FF",
		437421 => x"FF",
		437422 => x"FF",
		437423 => x"FF",
		437424 => x"FF",
		437425 => x"FF",
		437426 => x"FF",
		437427 => x"FF",
		437428 => x"FF",
		437429 => x"FF",
		437430 => x"FF",
		437431 => x"FF",
		437432 => x"FF",
		437433 => x"FF",
		437434 => x"FF",
		437435 => x"FF",
		437436 => x"FF",
		437437 => x"FF",
		437438 => x"FF",
		437439 => x"FF",
		437440 => x"FF",
		437441 => x"FF",
		437442 => x"FF",
		437443 => x"FF",
		437444 => x"FF",
		437445 => x"FF",
		437446 => x"FF",
		437447 => x"FF",
		437448 => x"FF",
		437449 => x"FF",
		437450 => x"FF",
		437451 => x"FF",
		437452 => x"FF",
		437453 => x"FF",
		437454 => x"FF",
		437455 => x"FF",
		437456 => x"FF",
		437457 => x"FF",
		437458 => x"FF",
		437459 => x"FF",
		437460 => x"FF",
		437461 => x"FF",
		437462 => x"FF",
		437463 => x"FF",
		437464 => x"FF",
		437465 => x"FF",
		437466 => x"FF",
		437467 => x"FF",
		437468 => x"FF",
		437469 => x"FF",
		437470 => x"FF",
		437471 => x"FF",
		437472 => x"FF",
		437473 => x"FF",
		437474 => x"FF",
		437475 => x"FF",
		437476 => x"FF",
		437477 => x"FF",
		437478 => x"FF",
		437479 => x"FF",
		437480 => x"FF",
		437481 => x"FF",
		437482 => x"FF",
		437483 => x"FF",
		437484 => x"FF",
		437485 => x"FF",
		437486 => x"FF",
		437487 => x"FF",
		437488 => x"FF",
		437489 => x"FF",
		437490 => x"FF",
		437491 => x"FF",
		437492 => x"FF",
		437493 => x"FF",
		437494 => x"FF",
		437495 => x"FF",
		437496 => x"FF",
		437497 => x"FF",
		437498 => x"FF",
		437499 => x"FF",
		437500 => x"FF",
		437501 => x"FF",
		437502 => x"FF",
		437503 => x"FF",
		437504 => x"FF",
		437505 => x"FF",
		437506 => x"FF",
		437507 => x"FF",
		437508 => x"FF",
		437509 => x"FF",
		437510 => x"FF",
		437511 => x"FF",
		437512 => x"FF",
		437513 => x"FF",
		437514 => x"FF",
		437515 => x"FF",
		437516 => x"FF",
		437517 => x"FF",
		437518 => x"FF",
		437519 => x"FF",
		437520 => x"FF",
		437521 => x"FF",
		437522 => x"FF",
		437523 => x"FF",
		437524 => x"FF",
		437525 => x"FF",
		437526 => x"FF",
		437527 => x"FF",
		437528 => x"FF",
		437529 => x"FF",
		437530 => x"FF",
		437531 => x"FF",
		437532 => x"FF",
		437533 => x"FF",
		437534 => x"FF",
		437535 => x"FF",
		437536 => x"FF",
		437537 => x"FF",
		437538 => x"FF",
		437539 => x"FF",
		437540 => x"FF",
		437541 => x"FF",
		437542 => x"FF",
		437543 => x"FF",
		437544 => x"FF",
		437545 => x"FF",
		437546 => x"FF",
		437547 => x"FF",
		437548 => x"FF",
		437549 => x"FF",
		437550 => x"FF",
		437551 => x"FF",
		437552 => x"FF",
		437553 => x"FF",
		437554 => x"FF",
		437555 => x"FF",
		437556 => x"FF",
		437557 => x"FF",
		437558 => x"FF",
		437559 => x"FF",
		437560 => x"FF",
		437561 => x"FF",
		437562 => x"FF",
		437563 => x"FF",
		437564 => x"FF",
		437565 => x"FF",
		437566 => x"FF",
		437567 => x"FF",
		437568 => x"FF",
		437569 => x"FF",
		437570 => x"FF",
		437571 => x"FF",
		437572 => x"FF",
		437573 => x"FF",
		437574 => x"FF",
		437575 => x"FF",
		437576 => x"FF",
		437577 => x"FF",
		437578 => x"FF",
		437579 => x"FF",
		437580 => x"FF",
		437581 => x"FF",
		437582 => x"FF",
		437583 => x"FF",
		437584 => x"FF",
		437585 => x"FF",
		437586 => x"FF",
		437587 => x"FF",
		437588 => x"FF",
		437589 => x"FF",
		437590 => x"FF",
		437591 => x"FF",
		437592 => x"FF",
		437593 => x"FF",
		437594 => x"FF",
		437595 => x"FF",
		437596 => x"FF",
		437597 => x"FF",
		437598 => x"FF",
		437599 => x"FF",
		437600 => x"FF",
		437601 => x"FF",
		437602 => x"FF",
		437603 => x"FF",
		437604 => x"FF",
		437605 => x"FF",
		437606 => x"FF",
		437607 => x"FF",
		437608 => x"FF",
		437609 => x"FF",
		437610 => x"FF",
		437611 => x"FF",
		437612 => x"FF",
		437613 => x"FF",
		437614 => x"FF",
		437615 => x"FF",
		437616 => x"FF",
		437617 => x"FF",
		437618 => x"FF",
		437619 => x"FF",
		437620 => x"FF",
		437621 => x"FF",
		437622 => x"FF",
		437623 => x"FF",
		437624 => x"FF",
		437625 => x"FF",
		437626 => x"FF",
		437627 => x"FF",
		437628 => x"FF",
		437629 => x"FF",
		437630 => x"FF",
		437631 => x"FF",
		437632 => x"FF",
		437633 => x"FF",
		437634 => x"FF",
		437635 => x"FF",
		437636 => x"FF",
		437637 => x"FF",
		437638 => x"FF",
		437639 => x"FF",
		437640 => x"FF",
		437641 => x"FF",
		437642 => x"FF",
		437643 => x"FF",
		437644 => x"FF",
		437645 => x"FF",
		437646 => x"FF",
		437647 => x"FF",
		437648 => x"FF",
		437649 => x"FF",
		437650 => x"FF",
		437651 => x"FF",
		437652 => x"FF",
		437653 => x"FF",
		437654 => x"FF",
		437655 => x"FF",
		437656 => x"FF",
		437657 => x"FF",
		437658 => x"FF",
		437659 => x"FF",
		437660 => x"FF",
		437661 => x"FF",
		437662 => x"FF",
		437663 => x"FF",
		437664 => x"FF",
		437665 => x"FF",
		437666 => x"FF",
		437667 => x"FF",
		437668 => x"FF",
		437669 => x"FF",
		437670 => x"FF",
		437671 => x"FF",
		437672 => x"FF",
		437673 => x"FF",
		437674 => x"FF",
		437675 => x"FF",
		437676 => x"FF",
		437677 => x"FF",
		437678 => x"FF",
		437679 => x"FF",
		437680 => x"FF",
		437681 => x"FF",
		437682 => x"FF",
		437683 => x"FF",
		437684 => x"FF",
		437685 => x"FF",
		437686 => x"FF",
		437687 => x"FF",
		437688 => x"FF",
		437689 => x"FF",
		437690 => x"FF",
		437691 => x"FF",
		437692 => x"FF",
		437693 => x"FF",
		437694 => x"FF",
		437695 => x"FF",
		437696 => x"FF",
		437697 => x"FF",
		437698 => x"FF",
		437699 => x"FF",
		437700 => x"FF",
		437701 => x"FF",
		437702 => x"FF",
		437703 => x"FF",
		437704 => x"FF",
		437705 => x"FF",
		437706 => x"FF",
		437707 => x"FF",
		437708 => x"FF",
		437709 => x"FF",
		437710 => x"FF",
		437711 => x"FF",
		437712 => x"FF",
		437713 => x"FF",
		437714 => x"FF",
		437715 => x"FF",
		437716 => x"FF",
		437717 => x"FF",
		437718 => x"FF",
		437719 => x"FF",
		437720 => x"FF",
		437721 => x"FF",
		437722 => x"FF",
		437723 => x"FF",
		437724 => x"FF",
		437725 => x"FF",
		437726 => x"FF",
		437727 => x"FF",
		437728 => x"FF",
		437729 => x"FF",
		437730 => x"FF",
		437731 => x"FF",
		437732 => x"FF",
		437733 => x"FF",
		437734 => x"FF",
		437735 => x"FF",
		437736 => x"FF",
		437737 => x"FF",
		437738 => x"FF",
		437739 => x"FF",
		437740 => x"FF",
		437741 => x"FF",
		437742 => x"FF",
		437743 => x"FF",
		437744 => x"FF",
		437745 => x"FF",
