		8200 => x"FF",
		8201 => x"FF",
		8202 => x"FF",
		8203 => x"FF",
		8204 => x"FF",
		8205 => x"FF",
		8206 => x"FF",
		8207 => x"FF",
		8208 => x"FF",
		8209 => x"FF",
		8210 => x"FF",
		8211 => x"FF",
		8212 => x"FF",
		8213 => x"FF",
		8214 => x"FF",
		8215 => x"FF",
		8216 => x"FF",
		8217 => x"FF",
		8218 => x"FF",
		8219 => x"FF",
		8220 => x"FF",
		8221 => x"FF",
		8222 => x"FF",
		8223 => x"FF",
		8224 => x"FF",
		8225 => x"FF",
		8226 => x"FF",
		8227 => x"FF",
		8228 => x"FF",
		8229 => x"FF",
		8230 => x"FF",
		8231 => x"FF",
		8232 => x"FF",
		8233 => x"FF",
		8234 => x"FF",
		8235 => x"FF",
		8236 => x"FF",
		8237 => x"FF",
		8238 => x"FF",
		8239 => x"FF",
		8240 => x"FF",
		8241 => x"FF",
		8242 => x"FF",
		8243 => x"FF",
		8244 => x"FF",
		8245 => x"FF",
		8246 => x"FF",
		8247 => x"FF",
		8248 => x"FF",
		8249 => x"FF",
		8250 => x"FF",
		8251 => x"FF",
		8252 => x"FF",
		8253 => x"FF",
		8254 => x"FF",
		8255 => x"FF",
		8256 => x"FF",
		8257 => x"FF",
		8258 => x"FF",
		8259 => x"FF",
		8260 => x"FF",
		8261 => x"FF",
		8262 => x"FF",
		8263 => x"FF",
		8264 => x"FF",
		8265 => x"FF",
		8266 => x"FF",
		8267 => x"FF",
		8268 => x"FF",
		8269 => x"FF",
		8270 => x"FF",
		8271 => x"FF",
		8272 => x"FF",
		8273 => x"FF",
		8274 => x"FF",
		8275 => x"FF",
		8276 => x"FF",
		8277 => x"FF",
		8278 => x"FF",
		8279 => x"FF",
		8280 => x"FF",
		8281 => x"FF",
		8282 => x"FF",
		8283 => x"FF",
		8284 => x"FF",
		8285 => x"FF",
		8286 => x"FF",
		8287 => x"FF",
		8288 => x"FF",
		8289 => x"FF",
		8290 => x"FF",
		8291 => x"FF",
		8292 => x"FF",
		8293 => x"FF",
		9224 => x"FF",
		9255 => x"FF",
		9286 => x"FF",
		9317 => x"FF",
		10248 => x"FF",
		10279 => x"FF",
		10310 => x"FF",
		10341 => x"FF",
		11272 => x"FF",
		11303 => x"FF",
		11334 => x"FF",
		11365 => x"FF",
		12296 => x"FF",
		12327 => x"FF",
		12358 => x"FF",
		12389 => x"FF",
		13320 => x"FF",
		13351 => x"FF",
		13382 => x"FF",
		13413 => x"FF",
		14344 => x"FF",
		14375 => x"FF",
		14406 => x"FF",
		14437 => x"FF",
		15368 => x"FF",
		15399 => x"FF",
		15430 => x"FF",
		15461 => x"FF",
		16392 => x"FF",
		16423 => x"FF",
		16454 => x"FF",
		16485 => x"FF",
		17416 => x"FF",
		17447 => x"FF",
		17478 => x"FF",
		17509 => x"FF",
		18440 => x"FF",
		18471 => x"FF",
		18502 => x"FF",
		18533 => x"FF",
		19464 => x"FF",
		19495 => x"FF",
		19526 => x"FF",
		19557 => x"FF",
		20488 => x"FF",
		20519 => x"FF",
		20550 => x"FF",
		20581 => x"FF",
		21512 => x"FF",
		21543 => x"FF",
		21574 => x"FF",
		21605 => x"FF",
		22536 => x"FF",
		22567 => x"FF",
		22598 => x"FF",
		22629 => x"FF",
		23560 => x"FF",
		23591 => x"FF",
		23622 => x"FF",
		23653 => x"FF",
		24584 => x"FF",
		24615 => x"FF",
		24646 => x"FF",
		24677 => x"FF",
		25608 => x"FF",
		25639 => x"FF",
		25670 => x"FF",
		25701 => x"FF",
		26632 => x"FF",
		26663 => x"FF",
		26694 => x"FF",
		26725 => x"FF",
		27656 => x"FF",
		27687 => x"FF",
		27718 => x"FF",
		27749 => x"FF",
		28680 => x"FF",
		28711 => x"FF",
		28742 => x"FF",
		28773 => x"FF",
		29704 => x"FF",
		29735 => x"FF",
		29766 => x"FF",
		29797 => x"FF",
		30728 => x"FF",
		30759 => x"FF",
		30790 => x"FF",
		30821 => x"FF",
		31752 => x"FF",
		31783 => x"FF",
		31814 => x"FF",
		31845 => x"FF",
		32776 => x"FF",
		32807 => x"FF",
		32838 => x"FF",
		32869 => x"FF",
		33800 => x"FF",
		33831 => x"FF",
		33862 => x"FF",
		33893 => x"FF",
		34824 => x"FF",
		34855 => x"FF",
		34886 => x"FF",
		34917 => x"FF",
		35848 => x"FF",
		35879 => x"FF",
		35910 => x"FF",
		35941 => x"FF",
		36872 => x"FF",
		36903 => x"FF",
		36934 => x"FF",
		36965 => x"FF",
		37896 => x"FF",
		37927 => x"FF",
		37958 => x"FF",
		37989 => x"FF",
		38920 => x"FF",
		38951 => x"FF",
		38982 => x"FF",
		39013 => x"FF",
		39944 => x"FF",
		39945 => x"FF",
		39946 => x"FF",
		39947 => x"FF",
		39948 => x"FF",
		39949 => x"FF",
		39950 => x"FF",
		39951 => x"FF",
		39952 => x"FF",
		39953 => x"FF",
		39954 => x"FF",
		39955 => x"FF",
		39956 => x"FF",
		39957 => x"FF",
		39958 => x"FF",
		39959 => x"FF",
		39960 => x"FF",
		39961 => x"FF",
		39962 => x"FF",
		39963 => x"FF",
		39964 => x"FF",
		39965 => x"FF",
		39966 => x"FF",
		39967 => x"FF",
		39968 => x"FF",
		39969 => x"FF",
		39970 => x"FF",
		39971 => x"FF",
		39972 => x"FF",
		39973 => x"FF",
		39974 => x"FF",
		39975 => x"FF",
		39976 => x"FF",
		39977 => x"FF",
		39978 => x"FF",
		39979 => x"FF",
		39980 => x"FF",
		39981 => x"FF",
		39982 => x"FF",
		39983 => x"FF",
		39984 => x"FF",
		39985 => x"FF",
		39986 => x"FF",
		39987 => x"FF",
		39988 => x"FF",
		39989 => x"FF",
		39990 => x"FF",
		39991 => x"FF",
		39992 => x"FF",
		39993 => x"FF",
		39994 => x"FF",
		39995 => x"FF",
		39996 => x"FF",
		39997 => x"FF",
		39998 => x"FF",
		39999 => x"FF",
		40000 => x"FF",
		40001 => x"FF",
		40002 => x"FF",
		40003 => x"FF",
		40004 => x"FF",
		40005 => x"FF",
		40006 => x"FF",
		40007 => x"FF",
		40008 => x"FF",
		40009 => x"FF",
		40010 => x"FF",
		40011 => x"FF",
		40012 => x"FF",
		40013 => x"FF",
		40014 => x"FF",
		40015 => x"FF",
		40016 => x"FF",
		40017 => x"FF",
		40018 => x"FF",
		40019 => x"FF",
		40020 => x"FF",
		40021 => x"FF",
		40022 => x"FF",
		40023 => x"FF",
		40024 => x"FF",
		40025 => x"FF",
		40026 => x"FF",
		40027 => x"FF",
		40028 => x"FF",
		40029 => x"FF",
		40030 => x"FF",
		40031 => x"FF",
		40032 => x"FF",
		40033 => x"FF",
		40034 => x"FF",
		40035 => x"FF",
		40036 => x"FF",
		40037 => x"FF",
		40968 => x"FF",
		40999 => x"FF",
		41030 => x"FF",
		41061 => x"FF",
		41992 => x"FF",
		42023 => x"FF",
		42054 => x"FF",
		42085 => x"FF",
		43016 => x"FF",
		43047 => x"FF",
		43078 => x"FF",
		43109 => x"FF",
		44040 => x"FF",
		44071 => x"FF",
		44102 => x"FF",
		44133 => x"FF",
		45064 => x"FF",
		45095 => x"FF",
		45126 => x"FF",
		45157 => x"FF",
		46088 => x"FF",
		46119 => x"FF",
		46150 => x"FF",
		46181 => x"FF",
		47112 => x"FF",
		47143 => x"FF",
		47174 => x"FF",
		47205 => x"FF",
		48136 => x"FF",
		48167 => x"FF",
		48198 => x"FF",
		48229 => x"FF",
		49160 => x"FF",
		49191 => x"FF",
		49222 => x"FF",
		49253 => x"FF",
		50184 => x"FF",
		50215 => x"FF",
		50246 => x"FF",
		50277 => x"FF",
		51208 => x"FF",
		51239 => x"FF",
		51270 => x"FF",
		51301 => x"FF",
		52232 => x"FF",
		52263 => x"FF",
		52294 => x"FF",
		52325 => x"FF",
		53256 => x"FF",
		53287 => x"FF",
		53318 => x"FF",
		53349 => x"FF",
		54280 => x"FF",
		54311 => x"FF",
		54342 => x"FF",
		54373 => x"FF",
		55304 => x"FF",
		55335 => x"FF",
		55366 => x"FF",
		55397 => x"FF",
		56328 => x"FF",
		56359 => x"FF",
		56390 => x"FF",
		56421 => x"FF",
		57352 => x"FF",
		57383 => x"FF",
		57414 => x"FF",
		57445 => x"FF",
		58376 => x"FF",
		58407 => x"FF",
		58438 => x"FF",
		58469 => x"FF",
		59400 => x"FF",
		59431 => x"FF",
		59462 => x"FF",
		59493 => x"FF",
		60424 => x"FF",
		60455 => x"FF",
		60486 => x"FF",
		60517 => x"FF",
		61448 => x"FF",
		61479 => x"FF",
		61510 => x"FF",
		61541 => x"FF",
		62472 => x"FF",
		62503 => x"FF",
		62534 => x"FF",
		62565 => x"FF",
		63496 => x"FF",
		63527 => x"FF",
		63558 => x"FF",
		63589 => x"FF",
		64520 => x"FF",
		64551 => x"FF",
		64582 => x"FF",
		64613 => x"FF",
		65544 => x"FF",
		65575 => x"FF",
		65606 => x"FF",
		65637 => x"FF",
		66568 => x"FF",
		66599 => x"FF",
		66630 => x"FF",
		66661 => x"FF",
		67592 => x"FF",
		67623 => x"FF",
		67654 => x"FF",
		67685 => x"FF",
		68616 => x"FF",
		68647 => x"FF",
		68678 => x"FF",
		68709 => x"FF",
		69640 => x"FF",
		69671 => x"FF",
		69702 => x"FF",
		69733 => x"FF",
		70664 => x"FF",
		70695 => x"FF",
		70726 => x"FF",
		70757 => x"FF",
		71688 => x"FF",
		71689 => x"FF",
		71690 => x"FF",
		71691 => x"FF",
		71692 => x"FF",
		71693 => x"FF",
		71694 => x"FF",
		71695 => x"FF",
		71696 => x"FF",
		71697 => x"FF",
		71698 => x"FF",
		71699 => x"FF",
		71700 => x"FF",
		71701 => x"FF",
		71702 => x"FF",
		71703 => x"FF",
		71704 => x"FF",
		71705 => x"FF",
		71706 => x"FF",
		71707 => x"FF",
		71708 => x"FF",
		71709 => x"FF",
		71710 => x"FF",
		71711 => x"FF",
		71712 => x"FF",
		71713 => x"FF",
		71714 => x"FF",
		71715 => x"FF",
		71716 => x"FF",
		71717 => x"FF",
		71718 => x"FF",
		71719 => x"FF",
		71720 => x"FF",
		71721 => x"FF",
		71722 => x"FF",
		71723 => x"FF",
		71724 => x"FF",
		71725 => x"FF",
		71726 => x"FF",
		71727 => x"FF",
		71728 => x"FF",
		71729 => x"FF",
		71730 => x"FF",
		71731 => x"FF",
		71732 => x"FF",
		71733 => x"FF",
		71734 => x"FF",
		71735 => x"FF",
		71736 => x"FF",
		71737 => x"FF",
		71738 => x"FF",
		71739 => x"FF",
		71740 => x"FF",
		71741 => x"FF",
		71742 => x"FF",
		71743 => x"FF",
		71744 => x"FF",
		71745 => x"FF",
		71746 => x"FF",
		71747 => x"FF",
		71748 => x"FF",
		71749 => x"FF",
		71750 => x"FF",
		71751 => x"FF",
		71752 => x"FF",
		71753 => x"FF",
		71754 => x"FF",
		71755 => x"FF",
		71756 => x"FF",
		71757 => x"FF",
		71758 => x"FF",
		71759 => x"FF",
		71760 => x"FF",
		71761 => x"FF",
		71762 => x"FF",
		71763 => x"FF",
		71764 => x"FF",
		71765 => x"FF",
		71766 => x"FF",
		71767 => x"FF",
		71768 => x"FF",
		71769 => x"FF",
		71770 => x"FF",
		71771 => x"FF",
		71772 => x"FF",
		71773 => x"FF",
		71774 => x"FF",
		71775 => x"FF",
		71776 => x"FF",
		71777 => x"FF",
		71778 => x"FF",
		71779 => x"FF",
		71780 => x"FF",
		71781 => x"FF",
		72712 => x"FF",
		72743 => x"FF",
		72774 => x"FF",
		72805 => x"FF",
		73736 => x"FF",
		73767 => x"FF",
		73798 => x"FF",
		73829 => x"FF",
		74760 => x"FF",
		74791 => x"FF",
		74822 => x"FF",
		74853 => x"FF",
		75784 => x"FF",
		75815 => x"FF",
		75846 => x"FF",
		75877 => x"FF",
		76808 => x"FF",
		76839 => x"FF",
		76870 => x"FF",
		76901 => x"FF",
		77832 => x"FF",
		77863 => x"FF",
		77894 => x"FF",
		77925 => x"FF",
		78856 => x"FF",
		78887 => x"FF",
		78918 => x"FF",
		78949 => x"FF",
		79880 => x"FF",
		79911 => x"FF",
		79942 => x"FF",
		79973 => x"FF",
		80904 => x"FF",
		80935 => x"FF",
		80966 => x"FF",
		80997 => x"FF",
		81928 => x"FF",
		81959 => x"FF",
		81990 => x"FF",
		82021 => x"FF",
		82952 => x"FF",
		82983 => x"FF",
		83014 => x"FF",
		83045 => x"FF",
		83976 => x"FF",
		84007 => x"FF",
		84038 => x"FF",
		84069 => x"FF",
		85000 => x"FF",
		85031 => x"FF",
		85062 => x"FF",
		85093 => x"FF",
		86024 => x"FF",
		86055 => x"FF",
		86086 => x"FF",
		86117 => x"FF",
		87048 => x"FF",
		87079 => x"FF",
		87110 => x"FF",
		87141 => x"FF",
		88072 => x"FF",
		88103 => x"FF",
		88134 => x"FF",
		88165 => x"FF",
		89096 => x"FF",
		89127 => x"FF",
		89158 => x"FF",
		89189 => x"FF",
		90120 => x"FF",
		90151 => x"FF",
		90182 => x"FF",
		90213 => x"FF",
		91144 => x"FF",
		91175 => x"FF",
		91206 => x"FF",
		91237 => x"FF",
		92168 => x"FF",
		92199 => x"FF",
		92230 => x"FF",
		92261 => x"FF",
		93192 => x"FF",
		93223 => x"FF",
		93254 => x"FF",
		93285 => x"FF",
		94216 => x"FF",
		94247 => x"FF",
		94278 => x"FF",
		94309 => x"FF",
		95240 => x"FF",
		95271 => x"FF",
		95302 => x"FF",
		95333 => x"FF",
		96264 => x"FF",
		96295 => x"FF",
		96326 => x"FF",
		96357 => x"FF",
		97288 => x"FF",
		97319 => x"FF",
		97350 => x"FF",
		97381 => x"FF",
		98312 => x"FF",
		98343 => x"FF",
		98374 => x"FF",
		98405 => x"FF",
		99336 => x"FF",
		99367 => x"FF",
		99398 => x"FF",
		99429 => x"FF",
		100360 => x"FF",
		100391 => x"FF",
		100422 => x"FF",
		100453 => x"FF",
		101384 => x"FF",
		101415 => x"FF",
		101446 => x"FF",
		101477 => x"FF",
		102408 => x"FF",
		102439 => x"FF",
		102470 => x"FF",
		102501 => x"FF",
		103432 => x"FF",
		103433 => x"FF",
		103434 => x"FF",
		103435 => x"FF",
		103436 => x"FF",
		103437 => x"FF",
		103438 => x"FF",
		103439 => x"FF",
		103440 => x"FF",
		103441 => x"FF",
		103442 => x"FF",
		103443 => x"FF",
		103444 => x"FF",
		103445 => x"FF",
		103446 => x"FF",
		103447 => x"FF",
		103448 => x"FF",
		103449 => x"FF",
		103450 => x"FF",
		103451 => x"FF",
		103452 => x"FF",
		103453 => x"FF",
		103454 => x"FF",
		103455 => x"FF",
		103456 => x"FF",
		103457 => x"FF",
		103458 => x"FF",
		103459 => x"FF",
		103460 => x"FF",
		103461 => x"FF",
		103462 => x"FF",
		103463 => x"FF",
		103464 => x"FF",
		103465 => x"FF",
		103466 => x"FF",
		103467 => x"FF",
		103468 => x"FF",
		103469 => x"FF",
		103470 => x"FF",
		103471 => x"FF",
		103472 => x"FF",
		103473 => x"FF",
		103474 => x"FF",
		103475 => x"FF",
		103476 => x"FF",
		103477 => x"FF",
		103478 => x"FF",
		103479 => x"FF",
		103480 => x"FF",
		103481 => x"FF",
		103482 => x"FF",
		103483 => x"FF",
		103484 => x"FF",
		103485 => x"FF",
		103486 => x"FF",
		103487 => x"FF",
		103488 => x"FF",
		103489 => x"FF",
		103490 => x"FF",
		103491 => x"FF",
		103492 => x"FF",
		103493 => x"FF",
		103494 => x"FF",
		103495 => x"FF",
		103496 => x"FF",
		103497 => x"FF",
		103498 => x"FF",
		103499 => x"FF",
		103500 => x"FF",
		103501 => x"FF",
		103502 => x"FF",
		103503 => x"FF",
		103504 => x"FF",
		103505 => x"FF",
		103506 => x"FF",
		103507 => x"FF",
		103508 => x"FF",
		103509 => x"FF",
		103510 => x"FF",
		103511 => x"FF",
		103512 => x"FF",
		103513 => x"FF",
		103514 => x"FF",
		103515 => x"FF",
		103516 => x"FF",
		103517 => x"FF",
		103518 => x"FF",
		103519 => x"FF",
		103520 => x"FF",
		103521 => x"FF",
		103522 => x"FF",
		103523 => x"FF",
		103524 => x"FF",
		103525 => x"FF",
