		49270 to 49649 => "11111111",
		50294 to 50673 => "11111111",
		51318 to 51697 => "11111111",
		52342 to 52721 => "11111111",
		53366 to 53745 => "11111111",
		54390 to 54394 => "11111111",
		54515 to 54519 => "11111111",
		54640 to 54644 => "11111111",
		54765 to 54769 => "11111111",
		55414 to 55418 => "11111111",
		55539 to 55543 => "11111111",
		55664 to 55668 => "11111111",
		55789 to 55793 => "11111111",
		56438 to 56442 => "11111111",
		56563 to 56567 => "11111111",
		56688 to 56692 => "11111111",
		56813 to 56817 => "11111111",
		57462 to 57466 => "11111111",
		57587 to 57591 => "11111111",
		57712 to 57716 => "11111111",
		57837 to 57841 => "11111111",
		58486 to 58490 => "11111111",
		58611 to 58615 => "11111111",
		58736 to 58740 => "11111111",
		58861 to 58865 => "11111111",
		59510 to 59514 => "11111111",
		59635 to 59639 => "11111111",
		59760 to 59764 => "11111111",
		59885 to 59889 => "11111111",
		60534 to 60538 => "11111111",
		60659 to 60663 => "11111111",
		60784 to 60788 => "11111111",
		60909 to 60913 => "11111111",
		61558 to 61562 => "11111111",
		61683 to 61687 => "11111111",
		61808 to 61812 => "11111111",
		61933 to 61937 => "11111111",
		62582 to 62586 => "11111111",
		62707 to 62711 => "11111111",
		62832 to 62836 => "11111111",
		62957 to 62961 => "11111111",
		63606 to 63610 => "11111111",
		63731 to 63735 => "11111111",
		63856 to 63860 => "11111111",
		63981 to 63985 => "11111111",
		64630 to 64634 => "11111111",
		64755 to 64759 => "11111111",
		64880 to 64884 => "11111111",
		65005 to 65009 => "11111111",
		65654 to 65658 => "11111111",
		65779 to 65783 => "11111111",
		65904 to 65908 => "11111111",
		66029 to 66033 => "11111111",
		66678 to 66682 => "11111111",
		66803 to 66807 => "11111111",
		66928 to 66932 => "11111111",
		67053 to 67057 => "11111111",
		67702 to 67706 => "11111111",
		67827 to 67831 => "11111111",
		67952 to 67956 => "11111111",
		68077 to 68081 => "11111111",
		68726 to 68730 => "11111111",
		68851 to 68855 => "11111111",
		68976 to 68980 => "11111111",
		69101 to 69105 => "11111111",
		69750 to 69754 => "11111111",
		69875 to 69879 => "11111111",
		70000 to 70004 => "11111111",
		70125 to 70129 => "11111111",
		70774 to 70778 => "11111111",
		70899 to 70903 => "11111111",
		71024 to 71028 => "11111111",
		71149 to 71153 => "11111111",
		71798 to 71802 => "11111111",
		71923 to 71927 => "11111111",
		72048 to 72052 => "11111111",
		72173 to 72177 => "11111111",
		72822 to 72826 => "11111111",
		72947 to 72951 => "11111111",
		73072 to 73076 => "11111111",
		73197 to 73201 => "11111111",
		73846 to 73850 => "11111111",
		73971 to 73975 => "11111111",
		74096 to 74100 => "11111111",
		74221 to 74225 => "11111111",
		74870 to 74874 => "11111111",
		74995 to 74999 => "11111111",
		75120 to 75124 => "11111111",
		75245 to 75249 => "11111111",
		75894 to 75898 => "11111111",
		76019 to 76023 => "11111111",
		76144 to 76148 => "11111111",
		76269 to 76273 => "11111111",
		76918 to 76922 => "11111111",
		77043 to 77047 => "11111111",
		77168 to 77172 => "11111111",
		77293 to 77297 => "11111111",
		77942 to 77946 => "11111111",
		78067 to 78071 => "11111111",
		78192 to 78196 => "11111111",
		78317 to 78321 => "11111111",
		78966 to 78970 => "11111111",
		79091 to 79095 => "11111111",
		79216 to 79220 => "11111111",
		79341 to 79345 => "11111111",
		79990 to 79994 => "11111111",
		80115 to 80119 => "11111111",
		80240 to 80244 => "11111111",
		80365 to 80369 => "11111111",
		81014 to 81018 => "11111111",
		81139 to 81143 => "11111111",
		81264 to 81268 => "11111111",
		81389 to 81393 => "11111111",
		82038 to 82042 => "11111111",
		82163 to 82167 => "11111111",
		82288 to 82292 => "11111111",
		82413 to 82417 => "11111111",
		83062 to 83066 => "11111111",
		83187 to 83191 => "11111111",
		83312 to 83316 => "11111111",
		83437 to 83441 => "11111111",
		84086 to 84090 => "11111111",
		84211 to 84215 => "11111111",
		84336 to 84340 => "11111111",
		84461 to 84465 => "11111111",
		85110 to 85114 => "11111111",
		85235 to 85239 => "11111111",
		85360 to 85364 => "11111111",
		85485 to 85489 => "11111111",
		86134 to 86138 => "11111111",
		86259 to 86263 => "11111111",
		86384 to 86388 => "11111111",
		86509 to 86513 => "11111111",
		87158 to 87162 => "11111111",
		87283 to 87287 => "11111111",
		87408 to 87412 => "11111111",
		87533 to 87537 => "11111111",
		88182 to 88186 => "11111111",
		88307 to 88311 => "11111111",
		88432 to 88436 => "11111111",
		88557 to 88561 => "11111111",
		89206 to 89210 => "11111111",
		89331 to 89335 => "11111111",
		89456 to 89460 => "11111111",
		89581 to 89585 => "11111111",
		90230 to 90234 => "11111111",
		90355 to 90359 => "11111111",
		90480 to 90484 => "11111111",
		90605 to 90609 => "11111111",
		91254 to 91258 => "11111111",
		91379 to 91383 => "11111111",
		91504 to 91508 => "11111111",
		91629 to 91633 => "11111111",
		92278 to 92282 => "11111111",
		92403 to 92407 => "11111111",
		92528 to 92532 => "11111111",
		92653 to 92657 => "11111111",
		93302 to 93306 => "11111111",
		93427 to 93431 => "11111111",
		93552 to 93556 => "11111111",
		93677 to 93681 => "11111111",
		94326 to 94330 => "11111111",
		94451 to 94455 => "11111111",
		94576 to 94580 => "11111111",
		94701 to 94705 => "11111111",
		95350 to 95354 => "11111111",
		95475 to 95479 => "11111111",
		95600 to 95604 => "11111111",
		95725 to 95729 => "11111111",
		96374 to 96378 => "11111111",
		96499 to 96503 => "11111111",
		96624 to 96628 => "11111111",
		96749 to 96753 => "11111111",
		97398 to 97402 => "11111111",
		97523 to 97527 => "11111111",
		97648 to 97652 => "11111111",
		97773 to 97777 => "11111111",
		98422 to 98426 => "11111111",
		98547 to 98551 => "11111111",
		98672 to 98676 => "11111111",
		98797 to 98801 => "11111111",
		99446 to 99450 => "11111111",
		99571 to 99575 => "11111111",
		99696 to 99700 => "11111111",
		99821 to 99825 => "11111111",
		100470 to 100474 => "11111111",
		100595 to 100599 => "11111111",
		100720 to 100724 => "11111111",
		100845 to 100849 => "11111111",
		101494 to 101498 => "11111111",
		101619 to 101623 => "11111111",
		101744 to 101748 => "11111111",
		101869 to 101873 => "11111111",
		102518 to 102522 => "11111111",
		102643 to 102647 => "11111111",
		102768 to 102772 => "11111111",
		102893 to 102897 => "11111111",
		103542 to 103546 => "11111111",
		103667 to 103671 => "11111111",
		103792 to 103796 => "11111111",
		103917 to 103921 => "11111111",
		104566 to 104570 => "11111111",
		104691 to 104695 => "11111111",
		104816 to 104820 => "11111111",
		104941 to 104945 => "11111111",
		105590 to 105594 => "11111111",
		105715 to 105719 => "11111111",
		105840 to 105844 => "11111111",
		105965 to 105969 => "11111111",
		106614 to 106618 => "11111111",
		106739 to 106743 => "11111111",
		106864 to 106868 => "11111111",
		106989 to 106993 => "11111111",
		107638 to 107642 => "11111111",
		107763 to 107767 => "11111111",
		107888 to 107892 => "11111111",
		108013 to 108017 => "11111111",
		108662 to 108666 => "11111111",
		108787 to 108791 => "11111111",
		108912 to 108916 => "11111111",
		109037 to 109041 => "11111111",
		109686 to 109690 => "11111111",
		109811 to 109815 => "11111111",
		109936 to 109940 => "11111111",
		110061 to 110065 => "11111111",
		110710 to 110714 => "11111111",
		110835 to 110839 => "11111111",
		110960 to 110964 => "11111111",
		111085 to 111089 => "11111111",
		111734 to 111738 => "11111111",
		111859 to 111863 => "11111111",
		111984 to 111988 => "11111111",
		112109 to 112113 => "11111111",
		112758 to 112762 => "11111111",
		112883 to 112887 => "11111111",
		113008 to 113012 => "11111111",
		113133 to 113137 => "11111111",
		113782 to 113786 => "11111111",
		113907 to 113911 => "11111111",
		114032 to 114036 => "11111111",
		114157 to 114161 => "11111111",
		114806 to 114810 => "11111111",
		114931 to 114935 => "11111111",
		115056 to 115060 => "11111111",
		115181 to 115185 => "11111111",
		115830 to 115834 => "11111111",
		115955 to 115959 => "11111111",
		116080 to 116084 => "11111111",
		116205 to 116209 => "11111111",
		116854 to 116858 => "11111111",
		116979 to 116983 => "11111111",
		117104 to 117108 => "11111111",
		117229 to 117233 => "11111111",
		117878 to 117882 => "11111111",
		118003 to 118007 => "11111111",
		118128 to 118132 => "11111111",
		118253 to 118257 => "11111111",
		118902 to 118906 => "11111111",
		119027 to 119031 => "11111111",
		119152 to 119156 => "11111111",
		119277 to 119281 => "11111111",
		119926 to 119930 => "11111111",
		120051 to 120055 => "11111111",
		120176 to 120180 => "11111111",
		120301 to 120305 => "11111111",
		120950 to 120954 => "11111111",
		121075 to 121079 => "11111111",
		121200 to 121204 => "11111111",
		121325 to 121329 => "11111111",
		121974 to 121978 => "11111111",
		122099 to 122103 => "11111111",
		122224 to 122228 => "11111111",
		122349 to 122353 => "11111111",
		122998 to 123002 => "11111111",
		123123 to 123127 => "11111111",
		123248 to 123252 => "11111111",
		123373 to 123377 => "11111111",
		124022 to 124026 => "11111111",
		124147 to 124151 => "11111111",
		124272 to 124276 => "11111111",
		124397 to 124401 => "11111111",
		125046 to 125050 => "11111111",
		125171 to 125175 => "11111111",
		125296 to 125300 => "11111111",
		125421 to 125425 => "11111111",
		126070 to 126074 => "11111111",
		126195 to 126199 => "11111111",
		126320 to 126324 => "11111111",
		126445 to 126449 => "11111111",
		127094 to 127098 => "11111111",
		127219 to 127223 => "11111111",
		127344 to 127348 => "11111111",
		127469 to 127473 => "11111111",
		128118 to 128122 => "11111111",
		128243 to 128247 => "11111111",
		128368 to 128372 => "11111111",
		128493 to 128497 => "11111111",
		129142 to 129146 => "11111111",
		129267 to 129271 => "11111111",
		129392 to 129396 => "11111111",
		129517 to 129521 => "11111111",
		130166 to 130170 => "11111111",
		130291 to 130295 => "11111111",
		130416 to 130420 => "11111111",
		130541 to 130545 => "11111111",
		131190 to 131194 => "11111111",
		131315 to 131319 => "11111111",
		131440 to 131444 => "11111111",
		131565 to 131569 => "11111111",
		132214 to 132218 => "11111111",
		132339 to 132343 => "11111111",
		132464 to 132468 => "11111111",
		132589 to 132593 => "11111111",
		133238 to 133242 => "11111111",
		133363 to 133367 => "11111111",
		133488 to 133492 => "11111111",
		133613 to 133617 => "11111111",
		134262 to 134266 => "11111111",
		134387 to 134391 => "11111111",
		134512 to 134516 => "11111111",
		134637 to 134641 => "11111111",
		135286 to 135290 => "11111111",
		135411 to 135415 => "11111111",
		135536 to 135540 => "11111111",
		135661 to 135665 => "11111111",
		136310 to 136314 => "11111111",
		136435 to 136439 => "11111111",
		136560 to 136564 => "11111111",
		136685 to 136689 => "11111111",
		137334 to 137338 => "11111111",
		137459 to 137463 => "11111111",
		137584 to 137588 => "11111111",
		137709 to 137713 => "11111111",
		138358 to 138362 => "11111111",
		138483 to 138487 => "11111111",
		138608 to 138612 => "11111111",
		138733 to 138737 => "11111111",
		139382 to 139386 => "11111111",
		139507 to 139511 => "11111111",
		139632 to 139636 => "11111111",
		139757 to 139761 => "11111111",
		140406 to 140410 => "11111111",
		140531 to 140535 => "11111111",
		140656 to 140660 => "11111111",
		140781 to 140785 => "11111111",
		141430 to 141434 => "11111111",
		141555 to 141559 => "11111111",
		141680 to 141684 => "11111111",
		141805 to 141809 => "11111111",
		142454 to 142458 => "11111111",
		142579 to 142583 => "11111111",
		142704 to 142708 => "11111111",
		142829 to 142833 => "11111111",
		143478 to 143482 => "11111111",
		143603 to 143607 => "11111111",
		143728 to 143732 => "11111111",
		143853 to 143857 => "11111111",
		144502 to 144506 => "11111111",
		144627 to 144631 => "11111111",
		144752 to 144756 => "11111111",
		144877 to 144881 => "11111111",
		145526 to 145530 => "11111111",
		145651 to 145655 => "11111111",
		145776 to 145780 => "11111111",
		145901 to 145905 => "11111111",
		146550 to 146554 => "11111111",
		146675 to 146679 => "11111111",
		146800 to 146804 => "11111111",
		146925 to 146929 => "11111111",
		147574 to 147578 => "11111111",
		147699 to 147703 => "11111111",
		147824 to 147828 => "11111111",
		147949 to 147953 => "11111111",
		148598 to 148602 => "11111111",
		148723 to 148727 => "11111111",
		148848 to 148852 => "11111111",
		148973 to 148977 => "11111111",
		149622 to 149626 => "11111111",
		149747 to 149751 => "11111111",
		149872 to 149876 => "11111111",
		149997 to 150001 => "11111111",
		150646 to 150650 => "11111111",
		150771 to 150775 => "11111111",
		150896 to 150900 => "11111111",
		151021 to 151025 => "11111111",
		151670 to 151674 => "11111111",
		151795 to 151799 => "11111111",
		151920 to 151924 => "11111111",
		152045 to 152049 => "11111111",
		152694 to 152698 => "11111111",
		152819 to 152823 => "11111111",
		152944 to 152948 => "11111111",
		153069 to 153073 => "11111111",
		153718 to 153722 => "11111111",
		153843 to 153847 => "11111111",
		153968 to 153972 => "11111111",
		154093 to 154097 => "11111111",
		154742 to 154746 => "11111111",
		154867 to 154871 => "11111111",
		154992 to 154996 => "11111111",
		155117 to 155121 => "11111111",
		155766 to 155770 => "11111111",
		155891 to 155895 => "11111111",
		156016 to 156020 => "11111111",
		156141 to 156145 => "11111111",
		156790 to 156794 => "11111111",
		156915 to 156919 => "11111111",
		157040 to 157044 => "11111111",
		157165 to 157169 => "11111111",
		157814 to 157818 => "11111111",
		157939 to 157943 => "11111111",
		158064 to 158068 => "11111111",
		158189 to 158193 => "11111111",
		158838 to 158842 => "11111111",
		158963 to 158967 => "11111111",
		159088 to 159092 => "11111111",
		159213 to 159217 => "11111111",
		159862 to 159866 => "11111111",
		159987 to 159991 => "11111111",
		160112 to 160116 => "11111111",
		160237 to 160241 => "11111111",
		160886 to 160890 => "11111111",
		161011 to 161015 => "11111111",
		161136 to 161140 => "11111111",
		161261 to 161265 => "11111111",
		161910 to 161914 => "11111111",
		162035 to 162039 => "11111111",
		162160 to 162164 => "11111111",
		162285 to 162289 => "11111111",
		162934 to 162938 => "11111111",
		163059 to 163063 => "11111111",
		163184 to 163188 => "11111111",
		163309 to 163313 => "11111111",
		163958 to 163962 => "11111111",
		164083 to 164087 => "11111111",
		164208 to 164212 => "11111111",
		164333 to 164337 => "11111111",
		164982 to 164986 => "11111111",
		165107 to 165111 => "11111111",
		165232 to 165236 => "11111111",
		165357 to 165361 => "11111111",
		166006 to 166010 => "11111111",
		166131 to 166135 => "11111111",
		166256 to 166260 => "11111111",
		166381 to 166385 => "11111111",
		167030 to 167034 => "11111111",
		167155 to 167159 => "11111111",
		167280 to 167284 => "11111111",
		167405 to 167409 => "11111111",
		168054 to 168058 => "11111111",
		168179 to 168183 => "11111111",
		168304 to 168308 => "11111111",
		168429 to 168433 => "11111111",
		169078 to 169082 => "11111111",
		169203 to 169207 => "11111111",
		169328 to 169332 => "11111111",
		169453 to 169457 => "11111111",
		170102 to 170106 => "11111111",
		170227 to 170231 => "11111111",
		170352 to 170356 => "11111111",
		170477 to 170481 => "11111111",
		171126 to 171130 => "11111111",
		171251 to 171255 => "11111111",
		171376 to 171380 => "11111111",
		171501 to 171505 => "11111111",
		172150 to 172154 => "11111111",
		172275 to 172279 => "11111111",
		172400 to 172404 => "11111111",
		172525 to 172529 => "11111111",
		173174 to 173178 => "11111111",
		173299 to 173303 => "11111111",
		173424 to 173428 => "11111111",
		173549 to 173553 => "11111111",
		174198 to 174202 => "11111111",
		174323 to 174327 => "11111111",
		174448 to 174452 => "11111111",
		174573 to 174577 => "11111111",
		175222 to 175226 => "11111111",
		175347 to 175351 => "11111111",
		175472 to 175476 => "11111111",
		175597 to 175601 => "11111111",
		176246 to 176250 => "11111111",
		176371 to 176375 => "11111111",
		176496 to 176500 => "11111111",
		176621 to 176625 => "11111111",
		177270 to 177649 => "11111111",
		178294 to 178673 => "11111111",
		179318 to 179697 => "11111111",
		180342 to 180721 => "11111111",
		181366 to 181745 => "11111111",
		182390 to 182394 => "11111111",
		182515 to 182519 => "11111111",
		182640 to 182644 => "11111111",
		182765 to 182769 => "11111111",
		183414 to 183418 => "11111111",
		183539 to 183543 => "11111111",
		183664 to 183668 => "11111111",
		183789 to 183793 => "11111111",
		184438 to 184442 => "11111111",
		184563 to 184567 => "11111111",
		184688 to 184692 => "11111111",
		184813 to 184817 => "11111111",
		185462 to 185466 => "11111111",
		185587 to 185591 => "11111111",
		185712 to 185716 => "11111111",
		185837 to 185841 => "11111111",
		186486 to 186490 => "11111111",
		186611 to 186615 => "11111111",
		186736 to 186740 => "11111111",
		186861 to 186865 => "11111111",
		187510 to 187514 => "11111111",
		187635 to 187639 => "11111111",
		187760 to 187764 => "11111111",
		187885 to 187889 => "11111111",
		188534 to 188538 => "11111111",
		188659 to 188663 => "11111111",
		188784 to 188788 => "11111111",
		188909 to 188913 => "11111111",
		189558 to 189562 => "11111111",
		189683 to 189687 => "11111111",
		189808 to 189812 => "11111111",
		189933 to 189937 => "11111111",
		190582 to 190586 => "11111111",
		190707 to 190711 => "11111111",
		190832 to 190836 => "11111111",
		190957 to 190961 => "11111111",
		191606 to 191610 => "11111111",
		191731 to 191735 => "11111111",
		191856 to 191860 => "11111111",
		191981 to 191985 => "11111111",
		192630 to 192634 => "11111111",
		192755 to 192759 => "11111111",
		192880 to 192884 => "11111111",
		193005 to 193009 => "11111111",
		193654 to 193658 => "11111111",
		193779 to 193783 => "11111111",
		193904 to 193908 => "11111111",
		194029 to 194033 => "11111111",
		194678 to 194682 => "11111111",
		194803 to 194807 => "11111111",
		194928 to 194932 => "11111111",
		195053 to 195057 => "11111111",
		195702 to 195706 => "11111111",
		195827 to 195831 => "11111111",
		195952 to 195956 => "11111111",
		196077 to 196081 => "11111111",
		196726 to 196730 => "11111111",
		196851 to 196855 => "11111111",
		196976 to 196980 => "11111111",
		197101 to 197105 => "11111111",
		197750 to 197754 => "11111111",
		197875 to 197879 => "11111111",
		198000 to 198004 => "11111111",
		198125 to 198129 => "11111111",
		198774 to 198778 => "11111111",
		198899 to 198903 => "11111111",
		199024 to 199028 => "11111111",
		199149 to 199153 => "11111111",
		199798 to 199802 => "11111111",
		199923 to 199927 => "11111111",
		200048 to 200052 => "11111111",
		200173 to 200177 => "11111111",
		200822 to 200826 => "11111111",
		200947 to 200951 => "11111111",
		201072 to 201076 => "11111111",
		201197 to 201201 => "11111111",
		201846 to 201850 => "11111111",
		201971 to 201975 => "11111111",
		202096 to 202100 => "11111111",
		202221 to 202225 => "11111111",
		202870 to 202874 => "11111111",
		202995 to 202999 => "11111111",
		203120 to 203124 => "11111111",
		203245 to 203249 => "11111111",
		203894 to 203898 => "11111111",
		204019 to 204023 => "11111111",
		204144 to 204148 => "11111111",
		204269 to 204273 => "11111111",
		204918 to 204922 => "11111111",
		205043 to 205047 => "11111111",
		205168 to 205172 => "11111111",
		205293 to 205297 => "11111111",
		205942 to 205946 => "11111111",
		206067 to 206071 => "11111111",
		206192 to 206196 => "11111111",
		206317 to 206321 => "11111111",
		206966 to 206970 => "11111111",
		207091 to 207095 => "11111111",
		207216 to 207220 => "11111111",
		207341 to 207345 => "11111111",
		207990 to 207994 => "11111111",
		208115 to 208119 => "11111111",
		208240 to 208244 => "11111111",
		208365 to 208369 => "11111111",
		209014 to 209018 => "11111111",
		209139 to 209143 => "11111111",
		209264 to 209268 => "11111111",
		209389 to 209393 => "11111111",
		210038 to 210042 => "11111111",
		210163 to 210167 => "11111111",
		210288 to 210292 => "11111111",
		210413 to 210417 => "11111111",
		211062 to 211066 => "11111111",
		211187 to 211191 => "11111111",
		211312 to 211316 => "11111111",
		211437 to 211441 => "11111111",
		212086 to 212090 => "11111111",
		212211 to 212215 => "11111111",
		212336 to 212340 => "11111111",
		212461 to 212465 => "11111111",
		213110 to 213114 => "11111111",
		213235 to 213239 => "11111111",
		213360 to 213364 => "11111111",
		213485 to 213489 => "11111111",
		214134 to 214138 => "11111111",
		214259 to 214263 => "11111111",
		214384 to 214388 => "11111111",
		214509 to 214513 => "11111111",
		215158 to 215162 => "11111111",
		215283 to 215287 => "11111111",
		215408 to 215412 => "11111111",
		215533 to 215537 => "11111111",
		216182 to 216186 => "11111111",
		216307 to 216311 => "11111111",
		216432 to 216436 => "11111111",
		216557 to 216561 => "11111111",
		217206 to 217210 => "11111111",
		217331 to 217335 => "11111111",
		217456 to 217460 => "11111111",
		217581 to 217585 => "11111111",
		218230 to 218234 => "11111111",
		218355 to 218359 => "11111111",
		218480 to 218484 => "11111111",
		218605 to 218609 => "11111111",
		219254 to 219258 => "11111111",
		219379 to 219383 => "11111111",
		219504 to 219508 => "11111111",
		219629 to 219633 => "11111111",
		220278 to 220282 => "11111111",
		220403 to 220407 => "11111111",
		220528 to 220532 => "11111111",
		220653 to 220657 => "11111111",
		221302 to 221306 => "11111111",
		221427 to 221431 => "11111111",
		221552 to 221556 => "11111111",
		221677 to 221681 => "11111111",
		222326 to 222330 => "11111111",
		222451 to 222455 => "11111111",
		222576 to 222580 => "11111111",
		222701 to 222705 => "11111111",
		223350 to 223354 => "11111111",
		223475 to 223479 => "11111111",
		223600 to 223604 => "11111111",
		223725 to 223729 => "11111111",
		224374 to 224378 => "11111111",
		224499 to 224503 => "11111111",
		224624 to 224628 => "11111111",
		224749 to 224753 => "11111111",
		225398 to 225402 => "11111111",
		225523 to 225527 => "11111111",
		225648 to 225652 => "11111111",
		225773 to 225777 => "11111111",
		226422 to 226426 => "11111111",
		226547 to 226551 => "11111111",
		226672 to 226676 => "11111111",
		226797 to 226801 => "11111111",
		227446 to 227450 => "11111111",
		227571 to 227575 => "11111111",
		227696 to 227700 => "11111111",
		227821 to 227825 => "11111111",
		228470 to 228474 => "11111111",
		228595 to 228599 => "11111111",
		228720 to 228724 => "11111111",
		228845 to 228849 => "11111111",
		229494 to 229498 => "11111111",
		229619 to 229623 => "11111111",
		229744 to 229748 => "11111111",
		229869 to 229873 => "11111111",
		230518 to 230522 => "11111111",
		230643 to 230647 => "11111111",
		230768 to 230772 => "11111111",
		230893 to 230897 => "11111111",
		231542 to 231546 => "11111111",
		231667 to 231671 => "11111111",
		231792 to 231796 => "11111111",
		231917 to 231921 => "11111111",
		232566 to 232570 => "11111111",
		232691 to 232695 => "11111111",
		232816 to 232820 => "11111111",
		232941 to 232945 => "11111111",
		233590 to 233594 => "11111111",
		233715 to 233719 => "11111111",
		233840 to 233844 => "11111111",
		233965 to 233969 => "11111111",
		234614 to 234618 => "11111111",
		234739 to 234743 => "11111111",
		234864 to 234868 => "11111111",
		234989 to 234993 => "11111111",
		235638 to 235642 => "11111111",
		235763 to 235767 => "11111111",
		235888 to 235892 => "11111111",
		236013 to 236017 => "11111111",
		236662 to 236666 => "11111111",
		236787 to 236791 => "11111111",
		236912 to 236916 => "11111111",
		237037 to 237041 => "11111111",
		237686 to 237690 => "11111111",
		237811 to 237815 => "11111111",
		237936 to 237940 => "11111111",
		238061 to 238065 => "11111111",
		238710 to 238714 => "11111111",
		238835 to 238839 => "11111111",
		238960 to 238964 => "11111111",
		239085 to 239089 => "11111111",
		239734 to 239738 => "11111111",
		239859 to 239863 => "11111111",
		239984 to 239988 => "11111111",
		240109 to 240113 => "11111111",
		240758 to 240762 => "11111111",
		240883 to 240887 => "11111111",
		241008 to 241012 => "11111111",
		241133 to 241137 => "11111111",
		241782 to 241786 => "11111111",
		241907 to 241911 => "11111111",
		242032 to 242036 => "11111111",
		242157 to 242161 => "11111111",
		242806 to 242810 => "11111111",
		242931 to 242935 => "11111111",
		243056 to 243060 => "11111111",
		243181 to 243185 => "11111111",
		243830 to 243834 => "11111111",
		243955 to 243959 => "11111111",
		244080 to 244084 => "11111111",
		244205 to 244209 => "11111111",
		244854 to 244858 => "11111111",
		244979 to 244983 => "11111111",
		245104 to 245108 => "11111111",
		245229 to 245233 => "11111111",
		245878 to 245882 => "11111111",
		246003 to 246007 => "11111111",
		246128 to 246132 => "11111111",
		246253 to 246257 => "11111111",
		246902 to 246906 => "11111111",
		247027 to 247031 => "11111111",
		247152 to 247156 => "11111111",
		247277 to 247281 => "11111111",
		247926 to 247930 => "11111111",
		248051 to 248055 => "11111111",
		248176 to 248180 => "11111111",
		248301 to 248305 => "11111111",
		248950 to 248954 => "11111111",
		249075 to 249079 => "11111111",
		249200 to 249204 => "11111111",
		249325 to 249329 => "11111111",
		249974 to 249978 => "11111111",
		250099 to 250103 => "11111111",
		250224 to 250228 => "11111111",
		250349 to 250353 => "11111111",
		250998 to 251002 => "11111111",
		251123 to 251127 => "11111111",
		251248 to 251252 => "11111111",
		251373 to 251377 => "11111111",
		252022 to 252026 => "11111111",
		252147 to 252151 => "11111111",
		252272 to 252276 => "11111111",
		252397 to 252401 => "11111111",
		253046 to 253050 => "11111111",
		253171 to 253175 => "11111111",
		253296 to 253300 => "11111111",
		253421 to 253425 => "11111111",
		254070 to 254074 => "11111111",
		254195 to 254199 => "11111111",
		254320 to 254324 => "11111111",
		254445 to 254449 => "11111111",
		255094 to 255098 => "11111111",
		255219 to 255223 => "11111111",
		255344 to 255348 => "11111111",
		255469 to 255473 => "11111111",
		256118 to 256122 => "11111111",
		256243 to 256247 => "11111111",
		256368 to 256372 => "11111111",
		256493 to 256497 => "11111111",
		257142 to 257146 => "11111111",
		257267 to 257271 => "11111111",
		257392 to 257396 => "11111111",
		257517 to 257521 => "11111111",
		258166 to 258170 => "11111111",
		258291 to 258295 => "11111111",
		258416 to 258420 => "11111111",
		258541 to 258545 => "11111111",
		259190 to 259194 => "11111111",
		259315 to 259319 => "11111111",
		259440 to 259444 => "11111111",
		259565 to 259569 => "11111111",
		260214 to 260218 => "11111111",
		260339 to 260343 => "11111111",
		260464 to 260468 => "11111111",
		260589 to 260593 => "11111111",
		261238 to 261242 => "11111111",
		261363 to 261367 => "11111111",
		261488 to 261492 => "11111111",
		261613 to 261617 => "11111111",
		262262 to 262266 => "11111111",
		262387 to 262391 => "11111111",
		262512 to 262516 => "11111111",
		262637 to 262641 => "11111111",
		263286 to 263290 => "11111111",
		263411 to 263415 => "11111111",
		263536 to 263540 => "11111111",
		263661 to 263665 => "11111111",
		264310 to 264314 => "11111111",
		264435 to 264439 => "11111111",
		264560 to 264564 => "11111111",
		264685 to 264689 => "11111111",
		265334 to 265338 => "11111111",
		265459 to 265463 => "11111111",
		265584 to 265588 => "11111111",
		265709 to 265713 => "11111111",
		266358 to 266362 => "11111111",
		266483 to 266487 => "11111111",
		266608 to 266612 => "11111111",
		266733 to 266737 => "11111111",
		267382 to 267386 => "11111111",
		267507 to 267511 => "11111111",
		267632 to 267636 => "11111111",
		267757 to 267761 => "11111111",
		268406 to 268410 => "11111111",
		268531 to 268535 => "11111111",
		268656 to 268660 => "11111111",
		268781 to 268785 => "11111111",
		269430 to 269434 => "11111111",
		269555 to 269559 => "11111111",
		269680 to 269684 => "11111111",
		269805 to 269809 => "11111111",
		270454 to 270458 => "11111111",
		270579 to 270583 => "11111111",
		270704 to 270708 => "11111111",
		270829 to 270833 => "11111111",
		271478 to 271482 => "11111111",
		271603 to 271607 => "11111111",
		271728 to 271732 => "11111111",
		271853 to 271857 => "11111111",
		272502 to 272506 => "11111111",
		272627 to 272631 => "11111111",
		272752 to 272756 => "11111111",
		272877 to 272881 => "11111111",
		273526 to 273530 => "11111111",
		273651 to 273655 => "11111111",
		273776 to 273780 => "11111111",
		273901 to 273905 => "11111111",
		274550 to 274554 => "11111111",
		274675 to 274679 => "11111111",
		274800 to 274804 => "11111111",
		274925 to 274929 => "11111111",
		275574 to 275578 => "11111111",
		275699 to 275703 => "11111111",
		275824 to 275828 => "11111111",
		275949 to 275953 => "11111111",
		276598 to 276602 => "11111111",
		276723 to 276727 => "11111111",
		276848 to 276852 => "11111111",
		276973 to 276977 => "11111111",
		277622 to 277626 => "11111111",
		277747 to 277751 => "11111111",
		277872 to 277876 => "11111111",
		277997 to 278001 => "11111111",
		278646 to 278650 => "11111111",
		278771 to 278775 => "11111111",
		278896 to 278900 => "11111111",
		279021 to 279025 => "11111111",
		279670 to 279674 => "11111111",
		279795 to 279799 => "11111111",
		279920 to 279924 => "11111111",
		280045 to 280049 => "11111111",
		280694 to 280698 => "11111111",
		280819 to 280823 => "11111111",
		280944 to 280948 => "11111111",
		281069 to 281073 => "11111111",
		281718 to 281722 => "11111111",
		281843 to 281847 => "11111111",
		281968 to 281972 => "11111111",
		282093 to 282097 => "11111111",
		282742 to 282746 => "11111111",
		282867 to 282871 => "11111111",
		282992 to 282996 => "11111111",
		283117 to 283121 => "11111111",
		283766 to 283770 => "11111111",
		283891 to 283895 => "11111111",
		284016 to 284020 => "11111111",
		284141 to 284145 => "11111111",
		284790 to 284794 => "11111111",
		284915 to 284919 => "11111111",
		285040 to 285044 => "11111111",
		285165 to 285169 => "11111111",
		285814 to 285818 => "11111111",
		285939 to 285943 => "11111111",
		286064 to 286068 => "11111111",
		286189 to 286193 => "11111111",
		286838 to 286842 => "11111111",
		286963 to 286967 => "11111111",
		287088 to 287092 => "11111111",
		287213 to 287217 => "11111111",
		287862 to 287866 => "11111111",
		287987 to 287991 => "11111111",
		288112 to 288116 => "11111111",
		288237 to 288241 => "11111111",
		288886 to 288890 => "11111111",
		289011 to 289015 => "11111111",
		289136 to 289140 => "11111111",
		289261 to 289265 => "11111111",
		289910 to 289914 => "11111111",
		290035 to 290039 => "11111111",
		290160 to 290164 => "11111111",
		290285 to 290289 => "11111111",
		290934 to 290938 => "11111111",
		291059 to 291063 => "11111111",
		291184 to 291188 => "11111111",
		291309 to 291313 => "11111111",
		291958 to 291962 => "11111111",
		292083 to 292087 => "11111111",
		292208 to 292212 => "11111111",
		292333 to 292337 => "11111111",
		292982 to 292986 => "11111111",
		293107 to 293111 => "11111111",
		293232 to 293236 => "11111111",
		293357 to 293361 => "11111111",
		294006 to 294010 => "11111111",
		294131 to 294135 => "11111111",
		294256 to 294260 => "11111111",
		294381 to 294385 => "11111111",
		295030 to 295034 => "11111111",
		295155 to 295159 => "11111111",
		295280 to 295284 => "11111111",
		295405 to 295409 => "11111111",
		296054 to 296058 => "11111111",
		296179 to 296183 => "11111111",
		296304 to 296308 => "11111111",
		296429 to 296433 => "11111111",
		297078 to 297082 => "11111111",
		297203 to 297207 => "11111111",
		297328 to 297332 => "11111111",
		297453 to 297457 => "11111111",
		298102 to 298106 => "11111111",
		298227 to 298231 => "11111111",
		298352 to 298356 => "11111111",
		298477 to 298481 => "11111111",
		299126 to 299130 => "11111111",
		299251 to 299255 => "11111111",
		299376 to 299380 => "11111111",
		299501 to 299505 => "11111111",
		300150 to 300154 => "11111111",
		300275 to 300279 => "11111111",
		300400 to 300404 => "11111111",
		300525 to 300529 => "11111111",
		301174 to 301178 => "11111111",
		301299 to 301303 => "11111111",
		301424 to 301428 => "11111111",
		301549 to 301553 => "11111111",
		302198 to 302202 => "11111111",
		302323 to 302327 => "11111111",
		302448 to 302452 => "11111111",
		302573 to 302577 => "11111111",
		303222 to 303226 => "11111111",
		303347 to 303351 => "11111111",
		303472 to 303476 => "11111111",
		303597 to 303601 => "11111111",
		304246 to 304250 => "11111111",
		304371 to 304375 => "11111111",
		304496 to 304500 => "11111111",
		304621 to 304625 => "11111111",
		305270 to 305649 => "11111111",
		306294 to 306673 => "11111111",
		307318 to 307697 => "11111111",
		308342 to 308721 => "11111111",
		309366 to 309745 => "11111111",
		310390 to 310394 => "11111111",
		310515 to 310519 => "11111111",
		310640 to 310644 => "11111111",
		310765 to 310769 => "11111111",
		311414 to 311418 => "11111111",
		311539 to 311543 => "11111111",
		311664 to 311668 => "11111111",
		311789 to 311793 => "11111111",
		312438 to 312442 => "11111111",
		312563 to 312567 => "11111111",
		312688 to 312692 => "11111111",
		312813 to 312817 => "11111111",
		313462 to 313466 => "11111111",
		313587 to 313591 => "11111111",
		313712 to 313716 => "11111111",
		313837 to 313841 => "11111111",
		314486 to 314490 => "11111111",
		314611 to 314615 => "11111111",
		314736 to 314740 => "11111111",
		314861 to 314865 => "11111111",
		315510 to 315514 => "11111111",
		315635 to 315639 => "11111111",
		315760 to 315764 => "11111111",
		315885 to 315889 => "11111111",
		316534 to 316538 => "11111111",
		316659 to 316663 => "11111111",
		316784 to 316788 => "11111111",
		316909 to 316913 => "11111111",
		317558 to 317562 => "11111111",
		317683 to 317687 => "11111111",
		317808 to 317812 => "11111111",
		317933 to 317937 => "11111111",
		318582 to 318586 => "11111111",
		318707 to 318711 => "11111111",
		318832 to 318836 => "11111111",
		318957 to 318961 => "11111111",
		319606 to 319610 => "11111111",
		319731 to 319735 => "11111111",
		319856 to 319860 => "11111111",
		319981 to 319985 => "11111111",
		320630 to 320634 => "11111111",
		320755 to 320759 => "11111111",
		320880 to 320884 => "11111111",
		321005 to 321009 => "11111111",
		321654 to 321658 => "11111111",
		321779 to 321783 => "11111111",
		321904 to 321908 => "11111111",
		322029 to 322033 => "11111111",
		322678 to 322682 => "11111111",
		322803 to 322807 => "11111111",
		322928 to 322932 => "11111111",
		323053 to 323057 => "11111111",
		323702 to 323706 => "11111111",
		323827 to 323831 => "11111111",
		323952 to 323956 => "11111111",
		324077 to 324081 => "11111111",
		324726 to 324730 => "11111111",
		324851 to 324855 => "11111111",
		324976 to 324980 => "11111111",
		325101 to 325105 => "11111111",
		325750 to 325754 => "11111111",
		325875 to 325879 => "11111111",
		326000 to 326004 => "11111111",
		326125 to 326129 => "11111111",
		326774 to 326778 => "11111111",
		326899 to 326903 => "11111111",
		327024 to 327028 => "11111111",
		327149 to 327153 => "11111111",
		327798 to 327802 => "11111111",
		327923 to 327927 => "11111111",
		328048 to 328052 => "11111111",
		328173 to 328177 => "11111111",
		328822 to 328826 => "11111111",
		328947 to 328951 => "11111111",
		329072 to 329076 => "11111111",
		329197 to 329201 => "11111111",
		329846 to 329850 => "11111111",
		329971 to 329975 => "11111111",
		330096 to 330100 => "11111111",
		330221 to 330225 => "11111111",
		330870 to 330874 => "11111111",
		330995 to 330999 => "11111111",
		331120 to 331124 => "11111111",
		331245 to 331249 => "11111111",
		331894 to 331898 => "11111111",
		332019 to 332023 => "11111111",
		332144 to 332148 => "11111111",
		332269 to 332273 => "11111111",
		332918 to 332922 => "11111111",
		333043 to 333047 => "11111111",
		333168 to 333172 => "11111111",
		333293 to 333297 => "11111111",
		333942 to 333946 => "11111111",
		334067 to 334071 => "11111111",
		334192 to 334196 => "11111111",
		334317 to 334321 => "11111111",
		334966 to 334970 => "11111111",
		335091 to 335095 => "11111111",
		335216 to 335220 => "11111111",
		335341 to 335345 => "11111111",
		335990 to 335994 => "11111111",
		336115 to 336119 => "11111111",
		336240 to 336244 => "11111111",
		336365 to 336369 => "11111111",
		337014 to 337018 => "11111111",
		337139 to 337143 => "11111111",
		337264 to 337268 => "11111111",
		337389 to 337393 => "11111111",
		338038 to 338042 => "11111111",
		338163 to 338167 => "11111111",
		338288 to 338292 => "11111111",
		338413 to 338417 => "11111111",
		339062 to 339066 => "11111111",
		339187 to 339191 => "11111111",
		339312 to 339316 => "11111111",
		339437 to 339441 => "11111111",
		340086 to 340090 => "11111111",
		340211 to 340215 => "11111111",
		340336 to 340340 => "11111111",
		340461 to 340465 => "11111111",
		341110 to 341114 => "11111111",
		341235 to 341239 => "11111111",
		341360 to 341364 => "11111111",
		341485 to 341489 => "11111111",
		342134 to 342138 => "11111111",
		342259 to 342263 => "11111111",
		342384 to 342388 => "11111111",
		342509 to 342513 => "11111111",
		343158 to 343162 => "11111111",
		343283 to 343287 => "11111111",
		343408 to 343412 => "11111111",
		343533 to 343537 => "11111111",
		344182 to 344186 => "11111111",
		344307 to 344311 => "11111111",
		344432 to 344436 => "11111111",
		344557 to 344561 => "11111111",
		345206 to 345210 => "11111111",
		345331 to 345335 => "11111111",
		345456 to 345460 => "11111111",
		345581 to 345585 => "11111111",
		346230 to 346234 => "11111111",
		346355 to 346359 => "11111111",
		346480 to 346484 => "11111111",
		346605 to 346609 => "11111111",
		347254 to 347258 => "11111111",
		347379 to 347383 => "11111111",
		347504 to 347508 => "11111111",
		347629 to 347633 => "11111111",
		348278 to 348282 => "11111111",
		348403 to 348407 => "11111111",
		348528 to 348532 => "11111111",
		348653 to 348657 => "11111111",
		349302 to 349306 => "11111111",
		349427 to 349431 => "11111111",
		349552 to 349556 => "11111111",
		349677 to 349681 => "11111111",
		350326 to 350330 => "11111111",
		350451 to 350455 => "11111111",
		350576 to 350580 => "11111111",
		350701 to 350705 => "11111111",
		351350 to 351354 => "11111111",
		351475 to 351479 => "11111111",
		351600 to 351604 => "11111111",
		351725 to 351729 => "11111111",
		352374 to 352378 => "11111111",
		352499 to 352503 => "11111111",
		352624 to 352628 => "11111111",
		352749 to 352753 => "11111111",
		353398 to 353402 => "11111111",
		353523 to 353527 => "11111111",
		353648 to 353652 => "11111111",
		353773 to 353777 => "11111111",
		354422 to 354426 => "11111111",
		354547 to 354551 => "11111111",
		354672 to 354676 => "11111111",
		354797 to 354801 => "11111111",
		355446 to 355450 => "11111111",
		355571 to 355575 => "11111111",
		355696 to 355700 => "11111111",
		355821 to 355825 => "11111111",
		356470 to 356474 => "11111111",
		356595 to 356599 => "11111111",
		356720 to 356724 => "11111111",
		356845 to 356849 => "11111111",
		357494 to 357498 => "11111111",
		357619 to 357623 => "11111111",
		357744 to 357748 => "11111111",
		357869 to 357873 => "11111111",
		358518 to 358522 => "11111111",
		358643 to 358647 => "11111111",
		358768 to 358772 => "11111111",
		358893 to 358897 => "11111111",
		359542 to 359546 => "11111111",
		359667 to 359671 => "11111111",
		359792 to 359796 => "11111111",
		359917 to 359921 => "11111111",
		360566 to 360570 => "11111111",
		360691 to 360695 => "11111111",
		360816 to 360820 => "11111111",
		360941 to 360945 => "11111111",
		361590 to 361594 => "11111111",
		361715 to 361719 => "11111111",
		361840 to 361844 => "11111111",
		361965 to 361969 => "11111111",
		362614 to 362618 => "11111111",
		362739 to 362743 => "11111111",
		362864 to 362868 => "11111111",
		362989 to 362993 => "11111111",
		363638 to 363642 => "11111111",
		363763 to 363767 => "11111111",
		363888 to 363892 => "11111111",
		364013 to 364017 => "11111111",
		364662 to 364666 => "11111111",
		364787 to 364791 => "11111111",
		364912 to 364916 => "11111111",
		365037 to 365041 => "11111111",
		365686 to 365690 => "11111111",
		365811 to 365815 => "11111111",
		365936 to 365940 => "11111111",
		366061 to 366065 => "11111111",
		366710 to 366714 => "11111111",
		366835 to 366839 => "11111111",
		366960 to 366964 => "11111111",
		367085 to 367089 => "11111111",
		367734 to 367738 => "11111111",
		367859 to 367863 => "11111111",
		367984 to 367988 => "11111111",
		368109 to 368113 => "11111111",
		368758 to 368762 => "11111111",
		368883 to 368887 => "11111111",
		369008 to 369012 => "11111111",
		369133 to 369137 => "11111111",
		369782 to 369786 => "11111111",
		369907 to 369911 => "11111111",
		370032 to 370036 => "11111111",
		370157 to 370161 => "11111111",
		370806 to 370810 => "11111111",
		370931 to 370935 => "11111111",
		371056 to 371060 => "11111111",
		371181 to 371185 => "11111111",
		371830 to 371834 => "11111111",
		371955 to 371959 => "11111111",
		372080 to 372084 => "11111111",
		372205 to 372209 => "11111111",
		372854 to 372858 => "11111111",
		372979 to 372983 => "11111111",
		373104 to 373108 => "11111111",
		373229 to 373233 => "11111111",
		373878 to 373882 => "11111111",
		374003 to 374007 => "11111111",
		374128 to 374132 => "11111111",
		374253 to 374257 => "11111111",
		374902 to 374906 => "11111111",
		375027 to 375031 => "11111111",
		375152 to 375156 => "11111111",
		375277 to 375281 => "11111111",
		375926 to 375930 => "11111111",
		376051 to 376055 => "11111111",
		376176 to 376180 => "11111111",
		376301 to 376305 => "11111111",
		376950 to 376954 => "11111111",
		377075 to 377079 => "11111111",
		377200 to 377204 => "11111111",
		377325 to 377329 => "11111111",
		377974 to 377978 => "11111111",
		378099 to 378103 => "11111111",
		378224 to 378228 => "11111111",
		378349 to 378353 => "11111111",
		378998 to 379002 => "11111111",
		379123 to 379127 => "11111111",
		379248 to 379252 => "11111111",
		379373 to 379377 => "11111111",
		380022 to 380026 => "11111111",
		380147 to 380151 => "11111111",
		380272 to 380276 => "11111111",
		380397 to 380401 => "11111111",
		381046 to 381050 => "11111111",
		381171 to 381175 => "11111111",
		381296 to 381300 => "11111111",
		381421 to 381425 => "11111111",
		382070 to 382074 => "11111111",
		382195 to 382199 => "11111111",
		382320 to 382324 => "11111111",
		382445 to 382449 => "11111111",
		383094 to 383098 => "11111111",
		383219 to 383223 => "11111111",
		383344 to 383348 => "11111111",
		383469 to 383473 => "11111111",
		384118 to 384122 => "11111111",
		384243 to 384247 => "11111111",
		384368 to 384372 => "11111111",
		384493 to 384497 => "11111111",
		385142 to 385146 => "11111111",
		385267 to 385271 => "11111111",
		385392 to 385396 => "11111111",
		385517 to 385521 => "11111111",
		386166 to 386170 => "11111111",
		386291 to 386295 => "11111111",
		386416 to 386420 => "11111111",
		386541 to 386545 => "11111111",
		387190 to 387194 => "11111111",
		387315 to 387319 => "11111111",
		387440 to 387444 => "11111111",
		387565 to 387569 => "11111111",
		388214 to 388218 => "11111111",
		388339 to 388343 => "11111111",
		388464 to 388468 => "11111111",
		388589 to 388593 => "11111111",
		389238 to 389242 => "11111111",
		389363 to 389367 => "11111111",
		389488 to 389492 => "11111111",
		389613 to 389617 => "11111111",
		390262 to 390266 => "11111111",
		390387 to 390391 => "11111111",
		390512 to 390516 => "11111111",
		390637 to 390641 => "11111111",
		391286 to 391290 => "11111111",
		391411 to 391415 => "11111111",
		391536 to 391540 => "11111111",
		391661 to 391665 => "11111111",
		392310 to 392314 => "11111111",
		392435 to 392439 => "11111111",
		392560 to 392564 => "11111111",
		392685 to 392689 => "11111111",
		393334 to 393338 => "11111111",
		393459 to 393463 => "11111111",
		393584 to 393588 => "11111111",
		393709 to 393713 => "11111111",
		394358 to 394362 => "11111111",
		394483 to 394487 => "11111111",
		394608 to 394612 => "11111111",
		394733 to 394737 => "11111111",
		395382 to 395386 => "11111111",
		395507 to 395511 => "11111111",
		395632 to 395636 => "11111111",
		395757 to 395761 => "11111111",
		396406 to 396410 => "11111111",
		396531 to 396535 => "11111111",
		396656 to 396660 => "11111111",
		396781 to 396785 => "11111111",
		397430 to 397434 => "11111111",
		397555 to 397559 => "11111111",
		397680 to 397684 => "11111111",
		397805 to 397809 => "11111111",
		398454 to 398458 => "11111111",
		398579 to 398583 => "11111111",
		398704 to 398708 => "11111111",
		398829 to 398833 => "11111111",
		399478 to 399482 => "11111111",
		399603 to 399607 => "11111111",
		399728 to 399732 => "11111111",
		399853 to 399857 => "11111111",
		400502 to 400506 => "11111111",
		400627 to 400631 => "11111111",
		400752 to 400756 => "11111111",
		400877 to 400881 => "11111111",
		401526 to 401530 => "11111111",
		401651 to 401655 => "11111111",
		401776 to 401780 => "11111111",
		401901 to 401905 => "11111111",
		402550 to 402554 => "11111111",
		402675 to 402679 => "11111111",
		402800 to 402804 => "11111111",
		402925 to 402929 => "11111111",
		403574 to 403578 => "11111111",
		403699 to 403703 => "11111111",
		403824 to 403828 => "11111111",
		403949 to 403953 => "11111111",
		404598 to 404602 => "11111111",
		404723 to 404727 => "11111111",
		404848 to 404852 => "11111111",
		404973 to 404977 => "11111111",
		405622 to 405626 => "11111111",
		405747 to 405751 => "11111111",
		405872 to 405876 => "11111111",
		405997 to 406001 => "11111111",
		406646 to 406650 => "11111111",
		406771 to 406775 => "11111111",
		406896 to 406900 => "11111111",
		407021 to 407025 => "11111111",
		407670 to 407674 => "11111111",
		407795 to 407799 => "11111111",
		407920 to 407924 => "11111111",
		408045 to 408049 => "11111111",
		408694 to 408698 => "11111111",
		408819 to 408823 => "11111111",
		408944 to 408948 => "11111111",
		409069 to 409073 => "11111111",
		409718 to 409722 => "11111111",
		409843 to 409847 => "11111111",
		409968 to 409972 => "11111111",
		410093 to 410097 => "11111111",
		410742 to 410746 => "11111111",
		410867 to 410871 => "11111111",
		410992 to 410996 => "11111111",
		411117 to 411121 => "11111111",
		411766 to 411770 => "11111111",
		411891 to 411895 => "11111111",
		412016 to 412020 => "11111111",
		412141 to 412145 => "11111111",
		412790 to 412794 => "11111111",
		412915 to 412919 => "11111111",
		413040 to 413044 => "11111111",
		413165 to 413169 => "11111111",
		413814 to 413818 => "11111111",
		413939 to 413943 => "11111111",
		414064 to 414068 => "11111111",
		414189 to 414193 => "11111111",
		414838 to 414842 => "11111111",
		414963 to 414967 => "11111111",
		415088 to 415092 => "11111111",
		415213 to 415217 => "11111111",
		415862 to 415866 => "11111111",
		415987 to 415991 => "11111111",
		416112 to 416116 => "11111111",
		416237 to 416241 => "11111111",
		416886 to 416890 => "11111111",
		417011 to 417015 => "11111111",
		417136 to 417140 => "11111111",
		417261 to 417265 => "11111111",
		417910 to 417914 => "11111111",
		418035 to 418039 => "11111111",
		418160 to 418164 => "11111111",
		418285 to 418289 => "11111111",
		418934 to 418938 => "11111111",
		419059 to 419063 => "11111111",
		419184 to 419188 => "11111111",
		419309 to 419313 => "11111111",
		419958 to 419962 => "11111111",
		420083 to 420087 => "11111111",
		420208 to 420212 => "11111111",
		420333 to 420337 => "11111111",
		420982 to 420986 => "11111111",
		421107 to 421111 => "11111111",
		421232 to 421236 => "11111111",
		421357 to 421361 => "11111111",
		422006 to 422010 => "11111111",
		422131 to 422135 => "11111111",
		422256 to 422260 => "11111111",
		422381 to 422385 => "11111111",
		423030 to 423034 => "11111111",
		423155 to 423159 => "11111111",
		423280 to 423284 => "11111111",
		423405 to 423409 => "11111111",
		424054 to 424058 => "11111111",
		424179 to 424183 => "11111111",
		424304 to 424308 => "11111111",
		424429 to 424433 => "11111111",
		425078 to 425082 => "11111111",
		425203 to 425207 => "11111111",
		425328 to 425332 => "11111111",
		425453 to 425457 => "11111111",
		426102 to 426106 => "11111111",
		426227 to 426231 => "11111111",
		426352 to 426356 => "11111111",
		426477 to 426481 => "11111111",
		427126 to 427130 => "11111111",
		427251 to 427255 => "11111111",
		427376 to 427380 => "11111111",
		427501 to 427505 => "11111111",
		428150 to 428154 => "11111111",
		428275 to 428279 => "11111111",
		428400 to 428404 => "11111111",
		428525 to 428529 => "11111111",
		429174 to 429178 => "11111111",
		429299 to 429303 => "11111111",
		429424 to 429428 => "11111111",
		429549 to 429553 => "11111111",
		430198 to 430202 => "11111111",
		430323 to 430327 => "11111111",
		430448 to 430452 => "11111111",
		430573 to 430577 => "11111111",
		431222 to 431226 => "11111111",
		431347 to 431351 => "11111111",
		431472 to 431476 => "11111111",
		431597 to 431601 => "11111111",
		432246 to 432250 => "11111111",
		432371 to 432375 => "11111111",
		432496 to 432500 => "11111111",
		432621 to 432625 => "11111111",
		433270 to 433649 => "11111111",
		434294 to 434673 => "11111111",
		435318 to 435697 => "11111111",
		436342 to 436721 => "11111111",
		437366 to 437745 => "11111111",
