		8200 to 8293 => "11111111",
		9224 to 9224 => "11111111",
		9255 to 9255 => "11111111",
		9286 to 9286 => "11111111",
		9317 to 9317 => "11111111",
		10248 to 10248 => "11111111",
		10279 to 10279 => "11111111",
		10310 to 10310 => "11111111",
		10341 to 10341 => "11111111",
		11272 to 11272 => "11111111",
		11303 to 11303 => "11111111",
		11334 to 11334 => "11111111",
		11365 to 11365 => "11111111",
		12296 to 12296 => "11111111",
		12327 to 12327 => "11111111",
		12358 to 12358 => "11111111",
		12389 to 12389 => "11111111",
		13320 to 13320 => "11111111",
		13351 to 13351 => "11111111",
		13382 to 13382 => "11111111",
		13413 to 13413 => "11111111",
		14344 to 14344 => "11111111",
		14375 to 14375 => "11111111",
		14406 to 14406 => "11111111",
		14437 to 14437 => "11111111",
		15368 to 15368 => "11111111",
		15399 to 15399 => "11111111",
		15430 to 15430 => "11111111",
		15461 to 15461 => "11111111",
		16392 to 16392 => "11111111",
		16423 to 16423 => "11111111",
		16454 to 16454 => "11111111",
		16485 to 16485 => "11111111",
		17416 to 17416 => "11111111",
		17447 to 17447 => "11111111",
		17478 to 17478 => "11111111",
		17509 to 17509 => "11111111",
		18440 to 18440 => "11111111",
		18471 to 18471 => "11111111",
		18502 to 18502 => "11111111",
		18533 to 18533 => "11111111",
		19464 to 19464 => "11111111",
		19495 to 19495 => "11111111",
		19526 to 19526 => "11111111",
		19557 to 19557 => "11111111",
		20488 to 20488 => "11111111",
		20519 to 20519 => "11111111",
		20550 to 20550 => "11111111",
		20581 to 20581 => "11111111",
		21512 to 21512 => "11111111",
		21543 to 21543 => "11111111",
		21574 to 21574 => "11111111",
		21605 to 21605 => "11111111",
		22536 to 22536 => "11111111",
		22567 to 22567 => "11111111",
		22598 to 22598 => "11111111",
		22629 to 22629 => "11111111",
		23560 to 23560 => "11111111",
		23591 to 23591 => "11111111",
		23622 to 23622 => "11111111",
		23653 to 23653 => "11111111",
		24584 to 24584 => "11111111",
		24615 to 24615 => "11111111",
		24646 to 24646 => "11111111",
		24677 to 24677 => "11111111",
		25608 to 25608 => "11111111",
		25639 to 25639 => "11111111",
		25670 to 25670 => "11111111",
		25701 to 25701 => "11111111",
		26632 to 26632 => "11111111",
		26663 to 26663 => "11111111",
		26694 to 26694 => "11111111",
		26725 to 26725 => "11111111",
		27656 to 27656 => "11111111",
		27687 to 27687 => "11111111",
		27718 to 27718 => "11111111",
		27749 to 27749 => "11111111",
		28680 to 28680 => "11111111",
		28711 to 28711 => "11111111",
		28742 to 28742 => "11111111",
		28773 to 28773 => "11111111",
		29704 to 29704 => "11111111",
		29735 to 29735 => "11111111",
		29766 to 29766 => "11111111",
		29797 to 29797 => "11111111",
		30728 to 30728 => "11111111",
		30759 to 30759 => "11111111",
		30790 to 30790 => "11111111",
		30821 to 30821 => "11111111",
		31752 to 31752 => "11111111",
		31783 to 31783 => "11111111",
		31814 to 31814 => "11111111",
		31845 to 31845 => "11111111",
		32776 to 32776 => "11111111",
		32807 to 32807 => "11111111",
		32838 to 32838 => "11111111",
		32869 to 32869 => "11111111",
		33800 to 33800 => "11111111",
		33831 to 33831 => "11111111",
		33862 to 33862 => "11111111",
		33893 to 33893 => "11111111",
		34824 to 34824 => "11111111",
		34855 to 34855 => "11111111",
		34886 to 34886 => "11111111",
		34917 to 34917 => "11111111",
		35848 to 35848 => "11111111",
		35879 to 35879 => "11111111",
		35910 to 35910 => "11111111",
		35941 to 35941 => "11111111",
		36872 to 36872 => "11111111",
		36903 to 36903 => "11111111",
		36934 to 36934 => "11111111",
		36965 to 36965 => "11111111",
		37896 to 37896 => "11111111",
		37927 to 37927 => "11111111",
		37958 to 37958 => "11111111",
		37989 to 37989 => "11111111",
		38920 to 38920 => "11111111",
		38951 to 38951 => "11111111",
		38982 to 38982 => "11111111",
		39013 to 39013 => "11111111",
		39944 to 40037 => "11111111",
		40968 to 40968 => "11111111",
		40999 to 40999 => "11111111",
		41030 to 41030 => "11111111",
		41061 to 41061 => "11111111",
		41992 to 41992 => "11111111",
		42023 to 42023 => "11111111",
		42054 to 42054 => "11111111",
		42085 to 42085 => "11111111",
		43016 to 43016 => "11111111",
		43047 to 43047 => "11111111",
		43078 to 43078 => "11111111",
		43109 to 43109 => "11111111",
		44040 to 44040 => "11111111",
		44071 to 44071 => "11111111",
		44102 to 44102 => "11111111",
		44133 to 44133 => "11111111",
		45064 to 45064 => "11111111",
		45095 to 45095 => "11111111",
		45126 to 45126 => "11111111",
		45157 to 45157 => "11111111",
		46088 to 46088 => "11111111",
		46119 to 46119 => "11111111",
		46150 to 46150 => "11111111",
		46181 to 46181 => "11111111",
		47112 to 47112 => "11111111",
		47143 to 47143 => "11111111",
		47174 to 47174 => "11111111",
		47205 to 47205 => "11111111",
		48136 to 48136 => "11111111",
		48167 to 48167 => "11111111",
		48198 to 48198 => "11111111",
		48229 to 48229 => "11111111",
		49160 to 49160 => "11111111",
		49191 to 49191 => "11111111",
		49222 to 49222 => "11111111",
		49253 to 49253 => "11111111",
		50184 to 50184 => "11111111",
		50215 to 50215 => "11111111",
		50246 to 50246 => "11111111",
		50277 to 50277 => "11111111",
		51208 to 51208 => "11111111",
		51239 to 51239 => "11111111",
		51270 to 51270 => "11111111",
		51301 to 51301 => "11111111",
		52232 to 52232 => "11111111",
		52263 to 52263 => "11111111",
		52294 to 52294 => "11111111",
		52325 to 52325 => "11111111",
		53256 to 53256 => "11111111",
		53287 to 53287 => "11111111",
		53318 to 53318 => "11111111",
		53349 to 53349 => "11111111",
		54280 to 54280 => "11111111",
		54311 to 54311 => "11111111",
		54342 to 54342 => "11111111",
		54373 to 54373 => "11111111",
		55304 to 55304 => "11111111",
		55335 to 55335 => "11111111",
		55366 to 55366 => "11111111",
		55397 to 55397 => "11111111",
		56328 to 56328 => "11111111",
		56359 to 56359 => "11111111",
		56390 to 56390 => "11111111",
		56421 to 56421 => "11111111",
		57352 to 57352 => "11111111",
		57383 to 57383 => "11111111",
		57414 to 57414 => "11111111",
		57445 to 57445 => "11111111",
		58376 to 58376 => "11111111",
		58407 to 58407 => "11111111",
		58438 to 58438 => "11111111",
		58469 to 58469 => "11111111",
		59400 to 59400 => "11111111",
		59431 to 59431 => "11111111",
		59462 to 59462 => "11111111",
		59493 to 59493 => "11111111",
		60424 to 60424 => "11111111",
		60455 to 60455 => "11111111",
		60486 to 60486 => "11111111",
		60517 to 60517 => "11111111",
		61448 to 61448 => "11111111",
		61479 to 61479 => "11111111",
		61510 to 61510 => "11111111",
		61541 to 61541 => "11111111",
		62472 to 62472 => "11111111",
		62503 to 62503 => "11111111",
		62534 to 62534 => "11111111",
		62565 to 62565 => "11111111",
		63496 to 63496 => "11111111",
		63527 to 63527 => "11111111",
		63558 to 63558 => "11111111",
		63589 to 63589 => "11111111",
		64520 to 64520 => "11111111",
		64551 to 64551 => "11111111",
		64582 to 64582 => "11111111",
		64613 to 64613 => "11111111",
		65544 to 65544 => "11111111",
		65575 to 65575 => "11111111",
		65606 to 65606 => "11111111",
		65637 to 65637 => "11111111",
		66568 to 66568 => "11111111",
		66599 to 66599 => "11111111",
		66630 to 66630 => "11111111",
		66661 to 66661 => "11111111",
		67592 to 67592 => "11111111",
		67623 to 67623 => "11111111",
		67654 to 67654 => "11111111",
		67685 to 67685 => "11111111",
		68616 to 68616 => "11111111",
		68647 to 68647 => "11111111",
		68678 to 68678 => "11111111",
		68709 to 68709 => "11111111",
		69640 to 69640 => "11111111",
		69671 to 69671 => "11111111",
		69702 to 69702 => "11111111",
		69733 to 69733 => "11111111",
		70664 to 70664 => "11111111",
		70695 to 70695 => "11111111",
		70726 to 70726 => "11111111",
		70757 to 70757 => "11111111",
		71688 to 71781 => "11111111",
		72712 to 72712 => "11111111",
		72743 to 72743 => "11111111",
		72774 to 72774 => "11111111",
		72805 to 72805 => "11111111",
		73736 to 73736 => "11111111",
		73767 to 73767 => "11111111",
		73798 to 73798 => "11111111",
		73829 to 73829 => "11111111",
		74760 to 74760 => "11111111",
		74791 to 74791 => "11111111",
		74822 to 74822 => "11111111",
		74853 to 74853 => "11111111",
		75784 to 75784 => "11111111",
		75815 to 75815 => "11111111",
		75846 to 75846 => "11111111",
		75877 to 75877 => "11111111",
		76808 to 76808 => "11111111",
		76839 to 76839 => "11111111",
		76870 to 76870 => "11111111",
		76901 to 76901 => "11111111",
		77832 to 77832 => "11111111",
		77863 to 77863 => "11111111",
		77894 to 77894 => "11111111",
		77925 to 77925 => "11111111",
		78856 to 78856 => "11111111",
		78887 to 78887 => "11111111",
		78918 to 78918 => "11111111",
		78949 to 78949 => "11111111",
		79880 to 79880 => "11111111",
		79911 to 79911 => "11111111",
		79942 to 79942 => "11111111",
		79973 to 79973 => "11111111",
		80904 to 80904 => "11111111",
		80935 to 80935 => "11111111",
		80966 to 80966 => "11111111",
		80997 to 80997 => "11111111",
		81928 to 81928 => "11111111",
		81959 to 81959 => "11111111",
		81990 to 81990 => "11111111",
		82021 to 82021 => "11111111",
		82952 to 82952 => "11111111",
		82983 to 82983 => "11111111",
		83014 to 83014 => "11111111",
		83045 to 83045 => "11111111",
		83976 to 83976 => "11111111",
		84007 to 84007 => "11111111",
		84038 to 84038 => "11111111",
		84069 to 84069 => "11111111",
		85000 to 85000 => "11111111",
		85031 to 85031 => "11111111",
		85062 to 85062 => "11111111",
		85093 to 85093 => "11111111",
		86024 to 86024 => "11111111",
		86055 to 86055 => "11111111",
		86086 to 86086 => "11111111",
		86117 to 86117 => "11111111",
		87048 to 87048 => "11111111",
		87079 to 87079 => "11111111",
		87110 to 87110 => "11111111",
		87141 to 87141 => "11111111",
		88072 to 88072 => "11111111",
		88103 to 88103 => "11111111",
		88134 to 88134 => "11111111",
		88165 to 88165 => "11111111",
		89096 to 89096 => "11111111",
		89127 to 89127 => "11111111",
		89158 to 89158 => "11111111",
		89189 to 89189 => "11111111",
		90120 to 90120 => "11111111",
		90151 to 90151 => "11111111",
		90182 to 90182 => "11111111",
		90213 to 90213 => "11111111",
		91144 to 91144 => "11111111",
		91175 to 91175 => "11111111",
		91206 to 91206 => "11111111",
		91237 to 91237 => "11111111",
		92168 to 92168 => "11111111",
		92199 to 92199 => "11111111",
		92230 to 92230 => "11111111",
		92261 to 92261 => "11111111",
		93192 to 93192 => "11111111",
		93223 to 93223 => "11111111",
		93254 to 93254 => "11111111",
		93285 to 93285 => "11111111",
		94216 to 94216 => "11111111",
		94247 to 94247 => "11111111",
		94278 to 94278 => "11111111",
		94309 to 94309 => "11111111",
		95240 to 95240 => "11111111",
		95271 to 95271 => "11111111",
		95302 to 95302 => "11111111",
		95333 to 95333 => "11111111",
		96264 to 96264 => "11111111",
		96295 to 96295 => "11111111",
		96326 to 96326 => "11111111",
		96357 to 96357 => "11111111",
		97288 to 97288 => "11111111",
		97319 to 97319 => "11111111",
		97350 to 97350 => "11111111",
		97381 to 97381 => "11111111",
		98312 to 98312 => "11111111",
		98343 to 98343 => "11111111",
		98374 to 98374 => "11111111",
		98405 to 98405 => "11111111",
		99336 to 99336 => "11111111",
		99367 to 99367 => "11111111",
		99398 to 99398 => "11111111",
		99429 to 99429 => "11111111",
		100360 to 100360 => "11111111",
		100391 to 100391 => "11111111",
		100422 to 100422 => "11111111",
		100453 to 100453 => "11111111",
		101384 to 101384 => "11111111",
		101415 to 101415 => "11111111",
		101446 to 101446 => "11111111",
		101477 to 101477 => "11111111",
		102408 to 102408 => "11111111",
		102439 to 102439 => "11111111",
		102470 to 102470 => "11111111",
		102501 to 102501 => "11111111",
		103432 to 103525 => "11111111",
