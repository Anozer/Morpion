		9225 to 9274 => "11111111",
		10249 to 10298 => "11111111",
		11273 to 11322 => "11111111",
		12297 to 12346 => "11111111",
		13321 to 13370 => "11111111",
		14345 to 14349 => "11111111",
		14360 to 14364 => "11111111",
		14375 to 14379 => "11111111",
		14390 to 14394 => "11111111",
		15369 to 15373 => "11111111",
		15384 to 15388 => "11111111",
		15399 to 15403 => "11111111",
		15414 to 15418 => "11111111",
		16393 to 16397 => "11111111",
		16408 to 16412 => "11111111",
		16423 to 16427 => "11111111",
		16438 to 16442 => "11111111",
		17417 to 17421 => "11111111",
		17432 to 17436 => "11111111",
		17447 to 17451 => "11111111",
		17462 to 17466 => "11111111",
		18441 to 18445 => "11111111",
		18456 to 18460 => "11111111",
		18471 to 18475 => "11111111",
		18486 to 18490 => "11111111",
		19465 to 19469 => "11111111",
		19480 to 19484 => "11111111",
		19495 to 19499 => "11111111",
		19510 to 19514 => "11111111",
		20489 to 20493 => "11111111",
		20504 to 20508 => "11111111",
		20519 to 20523 => "11111111",
		20534 to 20538 => "11111111",
		21513 to 21517 => "11111111",
		21528 to 21532 => "11111111",
		21543 to 21547 => "11111111",
		21558 to 21562 => "11111111",
		22537 to 22541 => "11111111",
		22552 to 22556 => "11111111",
		22567 to 22571 => "11111111",
		22582 to 22586 => "11111111",
		23561 to 23565 => "11111111",
		23576 to 23580 => "11111111",
		23591 to 23595 => "11111111",
		23606 to 23610 => "11111111",
		24585 to 24634 => "11111111",
		25609 to 25658 => "11111111",
		26633 to 26682 => "11111111",
		27657 to 27706 => "11111111",
		28681 to 28730 => "11111111",
		29705 to 29709 => "11111111",
		29720 to 29724 => "11111111",
		29735 to 29739 => "11111111",
		29750 to 29754 => "11111111",
		30729 to 30733 => "11111111",
		30744 to 30748 => "11111111",
		30759 to 30763 => "11111111",
		30774 to 30778 => "11111111",
		31753 to 31757 => "11111111",
		31768 to 31772 => "11111111",
		31783 to 31787 => "11111111",
		31798 to 31802 => "11111111",
		32777 to 32781 => "11111111",
		32792 to 32796 => "11111111",
		32807 to 32811 => "11111111",
		32822 to 32826 => "11111111",
		33801 to 33805 => "11111111",
		33816 to 33820 => "11111111",
		33831 to 33835 => "11111111",
		33846 to 33850 => "11111111",
		34825 to 34829 => "11111111",
		34840 to 34844 => "11111111",
		34855 to 34859 => "11111111",
		34870 to 34874 => "11111111",
		35849 to 35853 => "11111111",
		35864 to 35868 => "11111111",
		35879 to 35883 => "11111111",
		35894 to 35898 => "11111111",
		36873 to 36877 => "11111111",
		36888 to 36892 => "11111111",
		36903 to 36907 => "11111111",
		36918 to 36922 => "11111111",
		37897 to 37901 => "11111111",
		37912 to 37916 => "11111111",
		37927 to 37931 => "11111111",
		37942 to 37946 => "11111111",
		38921 to 38925 => "11111111",
		38936 to 38940 => "11111111",
		38951 to 38955 => "11111111",
		38966 to 38970 => "11111111",
		39945 to 39994 => "11111111",
		40969 to 41018 => "11111111",
		41993 to 42042 => "11111111",
		43017 to 43066 => "11111111",
		44041 to 44090 => "11111111",
		45065 to 45069 => "11111111",
		45080 to 45084 => "11111111",
		45095 to 45099 => "11111111",
		45110 to 45114 => "11111111",
		46089 to 46093 => "11111111",
		46104 to 46108 => "11111111",
		46119 to 46123 => "11111111",
		46134 to 46138 => "11111111",
		47113 to 47117 => "11111111",
		47128 to 47132 => "11111111",
		47143 to 47147 => "11111111",
		47158 to 47162 => "11111111",
		48137 to 48141 => "11111111",
		48152 to 48156 => "11111111",
		48167 to 48171 => "11111111",
		48182 to 48186 => "11111111",
		49161 to 49165 => "11111111",
		49176 to 49180 => "11111111",
		49191 to 49195 => "11111111",
		49206 to 49210 => "11111111",
		50185 to 50189 => "11111111",
		50200 to 50204 => "11111111",
		50215 to 50219 => "11111111",
		50230 to 50234 => "11111111",
		51209 to 51213 => "11111111",
		51224 to 51228 => "11111111",
		51239 to 51243 => "11111111",
		51254 to 51258 => "11111111",
		52233 to 52237 => "11111111",
		52248 to 52252 => "11111111",
		52263 to 52267 => "11111111",
		52278 to 52282 => "11111111",
		53257 to 53261 => "11111111",
		53272 to 53276 => "11111111",
		53287 to 53291 => "11111111",
		53302 to 53306 => "11111111",
		54281 to 54285 => "11111111",
		54296 to 54300 => "11111111",
		54311 to 54315 => "11111111",
		54326 to 54330 => "11111111",
		55305 to 55354 => "11111111",
		56329 to 56378 => "11111111",
		57353 to 57402 => "11111111",
		58377 to 58426 => "11111111",
		59401 to 59450 => "11111111",
