		6939 => x"FF",
		6940 => x"FF",
		6941 => x"FF",
		6942 => x"FF",
		6943 => x"FF",
		6944 => x"FF",
		6945 => x"FF",
		6946 => x"FF",
		6947 => x"FF",
		6948 => x"FF",
		6949 => x"FF",
		6950 => x"FF",
		6951 => x"FF",
		6952 => x"FF",
		6953 => x"FF",
		6954 => x"FF",
		6955 => x"FF",
		6956 => x"FF",
		6957 => x"FF",
		6958 => x"FF",
		6959 => x"FF",
		6960 => x"FF",
		6961 => x"FF",
		6962 => x"FF",
		6963 => x"FF",
		6964 => x"FF",
		6965 => x"FF",
		6966 => x"FF",
		6967 => x"FF",
		6968 => x"FF",
		6969 => x"FF",
		6970 => x"FF",
		6971 => x"FF",
		6972 => x"FF",
		6973 => x"FF",
		6974 => x"FF",
		6975 => x"FF",
		6976 => x"FF",
		6977 => x"FF",
		6978 => x"FF",
		6979 => x"FF",
		6980 => x"FF",
		6981 => x"FF",
		6982 => x"FF",
		6983 => x"FF",
		6984 => x"FF",
		6985 => x"FF",
		6986 => x"FF",
		6987 => x"FF",
		6988 => x"FF",
		6989 => x"FF",
		6990 => x"FF",
		6991 => x"FF",
		6992 => x"FF",
		6993 => x"FF",
		6994 => x"FF",
		6995 => x"FF",
		6996 => x"FF",
		6997 => x"FF",
		6998 => x"FF",
		6999 => x"FF",
		7000 => x"FF",
		7001 => x"FF",
		7002 => x"FF",
		7003 => x"FF",
		7004 => x"FF",
		7005 => x"FF",
		7006 => x"FF",
		7007 => x"FF",
		7008 => x"FF",
		7009 => x"FF",
		7010 => x"FF",
		7011 => x"FF",
		7012 => x"FF",
		7013 => x"FF",
		7014 => x"FF",
		7015 => x"FF",
		7016 => x"FF",
		7017 => x"FF",
		7018 => x"FF",
		7019 => x"FF",
		7020 => x"FF",
		7021 => x"FF",
		7022 => x"FF",
		7023 => x"FF",
		7024 => x"FF",
		7025 => x"FF",
		7026 => x"FF",
		7027 => x"FF",
		7028 => x"FF",
		7029 => x"FF",
		7030 => x"FF",
		7031 => x"FF",
		7032 => x"FF",
		7033 => x"FF",
		7034 => x"FF",
		7035 => x"FF",
		7036 => x"FF",
		7037 => x"FF",
		7038 => x"FF",
		7039 => x"FF",
		7040 => x"FF",
		7041 => x"FF",
		7042 => x"FF",
		7043 => x"FF",
		7044 => x"FF",
		7045 => x"FF",
		7046 => x"FF",
		7047 => x"FF",
		7048 => x"FF",
		7049 => x"FF",
		7050 => x"FF",
		7051 => x"FF",
		7052 => x"FF",
		7053 => x"FF",
		7054 => x"FF",
		7055 => x"FF",
		7056 => x"FF",
		7057 => x"FF",
		7058 => x"FF",
		7059 => x"FF",
		7060 => x"FF",
		7061 => x"FF",
		7062 => x"FF",
		7063 => x"FF",
		7064 => x"FF",
		7065 => x"FF",
		7066 => x"FF",
		7067 => x"FF",
		7068 => x"FF",
		7069 => x"FF",
		7070 => x"FF",
		7071 => x"FF",
		7072 => x"FF",
		7073 => x"FF",
		7074 => x"FF",
		7075 => x"FF",
		7076 => x"FF",
		7077 => x"FF",
		7078 => x"FF",
		7079 => x"FF",
		7080 => x"FF",
		7081 => x"FF",
		7082 => x"FF",
		7083 => x"FF",
		7084 => x"FF",
		7085 => x"FF",
		7086 => x"FF",
		7087 => x"FF",
		7088 => x"FF",
		7089 => x"FF",
		7090 => x"FF",
		7091 => x"FF",
		7092 => x"FF",
		7093 => x"FF",
		7094 => x"FF",
		7095 => x"FF",
		7096 => x"FF",
		7097 => x"FF",
		7098 => x"FF",
		7099 => x"FF",
		7100 => x"FF",
		7101 => x"FF",
		7102 => x"FF",
		7103 => x"FF",
		7104 => x"FF",
		7105 => x"FF",
		7106 => x"FF",
		7107 => x"FF",
		7108 => x"FF",
		7109 => x"FF",
		7110 => x"FF",
		7111 => x"FF",
		7112 => x"FF",
		7113 => x"FF",
		7114 => x"FF",
		7115 => x"FF",
		7116 => x"FF",
		7117 => x"FF",
		7118 => x"FF",
		7119 => x"FF",
		7120 => x"FF",
		7121 => x"FF",
		7122 => x"FF",
		7123 => x"FF",
		7124 => x"FF",
		7125 => x"FF",
		7126 => x"FF",
		7127 => x"FF",
		7128 => x"FF",
		7129 => x"FF",
		7130 => x"FF",
		7195 => x"FF",
		7196 => x"FF",
		7197 => x"FF",
		7198 => x"FF",
		7199 => x"FF",
		7200 => x"FF",
		7201 => x"FF",
		7202 => x"FF",
		7203 => x"FF",
		7204 => x"FF",
		7205 => x"FF",
		7206 => x"FF",
		7207 => x"FF",
		7208 => x"FF",
		7209 => x"FF",
		7210 => x"FF",
		7211 => x"FF",
		7212 => x"FF",
		7213 => x"FF",
		7214 => x"FF",
		7215 => x"FF",
		7216 => x"FF",
		7217 => x"FF",
		7218 => x"FF",
		7219 => x"FF",
		7220 => x"FF",
		7221 => x"FF",
		7222 => x"FF",
		7223 => x"FF",
		7224 => x"FF",
		7225 => x"FF",
		7226 => x"FF",
		7227 => x"FF",
		7228 => x"FF",
		7229 => x"FF",
		7230 => x"FF",
		7231 => x"FF",
		7232 => x"FF",
		7233 => x"FF",
		7234 => x"FF",
		7235 => x"FF",
		7236 => x"FF",
		7237 => x"FF",
		7238 => x"FF",
		7239 => x"FF",
		7240 => x"FF",
		7241 => x"FF",
		7242 => x"FF",
		7243 => x"FF",
		7244 => x"FF",
		7245 => x"FF",
		7246 => x"FF",
		7247 => x"FF",
		7248 => x"FF",
		7249 => x"FF",
		7250 => x"FF",
		7251 => x"FF",
		7252 => x"FF",
		7253 => x"FF",
		7254 => x"FF",
		7255 => x"FF",
		7256 => x"FF",
		7257 => x"FF",
		7258 => x"FF",
		7259 => x"FF",
		7260 => x"FF",
		7261 => x"FF",
		7262 => x"FF",
		7263 => x"FF",
		7264 => x"FF",
		7265 => x"FF",
		7266 => x"FF",
		7267 => x"FF",
		7268 => x"FF",
		7269 => x"FF",
		7270 => x"FF",
		7271 => x"FF",
		7272 => x"FF",
		7273 => x"FF",
		7274 => x"FF",
		7275 => x"FF",
		7276 => x"FF",
		7277 => x"FF",
		7278 => x"FF",
		7279 => x"FF",
		7280 => x"FF",
		7281 => x"FF",
		7282 => x"FF",
		7283 => x"FF",
		7284 => x"FF",
		7285 => x"FF",
		7286 => x"FF",
		7287 => x"FF",
		7288 => x"FF",
		7289 => x"FF",
		7290 => x"FF",
		7291 => x"FF",
		7292 => x"FF",
		7293 => x"FF",
		7294 => x"FF",
		7295 => x"FF",
		7296 => x"FF",
		7297 => x"FF",
		7298 => x"FF",
		7299 => x"FF",
		7300 => x"FF",
		7301 => x"FF",
		7302 => x"FF",
		7303 => x"FF",
		7304 => x"FF",
		7305 => x"FF",
		7306 => x"FF",
		7307 => x"FF",
		7308 => x"FF",
		7309 => x"FF",
		7310 => x"FF",
		7311 => x"FF",
		7312 => x"FF",
		7313 => x"FF",
		7314 => x"FF",
		7315 => x"FF",
		7316 => x"FF",
		7317 => x"FF",
		7318 => x"FF",
		7319 => x"FF",
		7320 => x"FF",
		7321 => x"FF",
		7322 => x"FF",
		7323 => x"FF",
		7324 => x"FF",
		7325 => x"FF",
		7326 => x"FF",
		7327 => x"FF",
		7328 => x"FF",
		7329 => x"FF",
		7330 => x"FF",
		7331 => x"FF",
		7332 => x"FF",
		7333 => x"FF",
		7334 => x"FF",
		7335 => x"FF",
		7336 => x"FF",
		7337 => x"FF",
		7338 => x"FF",
		7339 => x"FF",
		7340 => x"FF",
		7341 => x"FF",
		7342 => x"FF",
		7343 => x"FF",
		7344 => x"FF",
		7345 => x"FF",
		7346 => x"FF",
		7347 => x"FF",
		7348 => x"FF",
		7349 => x"FF",
		7350 => x"FF",
		7351 => x"FF",
		7352 => x"FF",
		7353 => x"FF",
		7354 => x"FF",
		7355 => x"FF",
		7356 => x"FF",
		7357 => x"FF",
		7358 => x"FF",
		7359 => x"FF",
		7360 => x"FF",
		7361 => x"FF",
		7362 => x"FF",
		7363 => x"FF",
		7364 => x"FF",
		7365 => x"FF",
		7366 => x"FF",
		7367 => x"FF",
		7368 => x"FF",
		7369 => x"FF",
		7370 => x"FF",
		7371 => x"FF",
		7372 => x"FF",
		7373 => x"FF",
		7374 => x"FF",
		7375 => x"FF",
		7376 => x"FF",
		7377 => x"FF",
		7378 => x"FF",
		7379 => x"FF",
		7380 => x"FF",
		7381 => x"FF",
		7382 => x"FF",
		7383 => x"FF",
		7384 => x"FF",
		7385 => x"FF",
		7386 => x"FF",
		7451 => x"FF",
		7452 => x"FF",
		7453 => x"FF",
		7454 => x"FF",
		7455 => x"FF",
		7456 => x"FF",
		7457 => x"FF",
		7458 => x"FF",
		7459 => x"FF",
		7460 => x"FF",
		7461 => x"FF",
		7462 => x"FF",
		7463 => x"FF",
		7464 => x"FF",
		7465 => x"FF",
		7466 => x"FF",
		7467 => x"FF",
		7468 => x"FF",
		7469 => x"FF",
		7470 => x"FF",
		7471 => x"FF",
		7472 => x"FF",
		7473 => x"FF",
		7474 => x"FF",
		7475 => x"FF",
		7476 => x"FF",
		7477 => x"FF",
		7478 => x"FF",
		7479 => x"FF",
		7480 => x"FF",
		7481 => x"FF",
		7482 => x"FF",
		7483 => x"FF",
		7484 => x"FF",
		7485 => x"FF",
		7486 => x"FF",
		7487 => x"FF",
		7488 => x"FF",
		7489 => x"FF",
		7490 => x"FF",
		7491 => x"FF",
		7492 => x"FF",
		7493 => x"FF",
		7494 => x"FF",
		7495 => x"FF",
		7496 => x"FF",
		7497 => x"FF",
		7498 => x"FF",
		7499 => x"FF",
		7500 => x"FF",
		7501 => x"FF",
		7502 => x"FF",
		7503 => x"FF",
		7504 => x"FF",
		7505 => x"FF",
		7506 => x"FF",
		7507 => x"FF",
		7508 => x"FF",
		7509 => x"FF",
		7510 => x"FF",
		7511 => x"FF",
		7512 => x"FF",
		7513 => x"FF",
		7514 => x"FF",
		7515 => x"FF",
		7516 => x"FF",
		7517 => x"FF",
		7518 => x"FF",
		7519 => x"FF",
		7520 => x"FF",
		7521 => x"FF",
		7522 => x"FF",
		7523 => x"FF",
		7524 => x"FF",
		7525 => x"FF",
		7526 => x"FF",
		7527 => x"FF",
		7528 => x"FF",
		7529 => x"FF",
		7530 => x"FF",
		7531 => x"FF",
		7532 => x"FF",
		7533 => x"FF",
		7534 => x"FF",
		7535 => x"FF",
		7536 => x"FF",
		7537 => x"FF",
		7538 => x"FF",
		7539 => x"FF",
		7540 => x"FF",
		7541 => x"FF",
		7542 => x"FF",
		7543 => x"FF",
		7544 => x"FF",
		7545 => x"FF",
		7546 => x"FF",
		7547 => x"FF",
		7548 => x"FF",
		7549 => x"FF",
		7550 => x"FF",
		7551 => x"FF",
		7552 => x"FF",
		7553 => x"FF",
		7554 => x"FF",
		7555 => x"FF",
		7556 => x"FF",
		7557 => x"FF",
		7558 => x"FF",
		7559 => x"FF",
		7560 => x"FF",
		7561 => x"FF",
		7562 => x"FF",
		7563 => x"FF",
		7564 => x"FF",
		7565 => x"FF",
		7566 => x"FF",
		7567 => x"FF",
		7568 => x"FF",
		7569 => x"FF",
		7570 => x"FF",
		7571 => x"FF",
		7572 => x"FF",
		7573 => x"FF",
		7574 => x"FF",
		7575 => x"FF",
		7576 => x"FF",
		7577 => x"FF",
		7578 => x"FF",
		7579 => x"FF",
		7580 => x"FF",
		7581 => x"FF",
		7582 => x"FF",
		7583 => x"FF",
		7584 => x"FF",
		7585 => x"FF",
		7586 => x"FF",
		7587 => x"FF",
		7588 => x"FF",
		7589 => x"FF",
		7590 => x"FF",
		7591 => x"FF",
		7592 => x"FF",
		7593 => x"FF",
		7594 => x"FF",
		7595 => x"FF",
		7596 => x"FF",
		7597 => x"FF",
		7598 => x"FF",
		7599 => x"FF",
		7600 => x"FF",
		7601 => x"FF",
		7602 => x"FF",
		7603 => x"FF",
		7604 => x"FF",
		7605 => x"FF",
		7606 => x"FF",
		7607 => x"FF",
		7608 => x"FF",
		7609 => x"FF",
		7610 => x"FF",
		7611 => x"FF",
		7612 => x"FF",
		7613 => x"FF",
		7614 => x"FF",
		7615 => x"FF",
		7616 => x"FF",
		7617 => x"FF",
		7618 => x"FF",
		7619 => x"FF",
		7620 => x"FF",
		7621 => x"FF",
		7622 => x"FF",
		7623 => x"FF",
		7624 => x"FF",
		7625 => x"FF",
		7626 => x"FF",
		7627 => x"FF",
		7628 => x"FF",
		7629 => x"FF",
		7630 => x"FF",
		7631 => x"FF",
		7632 => x"FF",
		7633 => x"FF",
		7634 => x"FF",
		7635 => x"FF",
		7636 => x"FF",
		7637 => x"FF",
		7638 => x"FF",
		7639 => x"FF",
		7640 => x"FF",
		7641 => x"FF",
		7642 => x"FF",
		7707 => x"FF",
		7708 => x"FF",
		7709 => x"FF",
		7770 => x"FF",
		7771 => x"FF",
		7772 => x"FF",
		7833 => x"FF",
		7834 => x"FF",
		7835 => x"FF",
		7896 => x"FF",
		7897 => x"FF",
		7898 => x"FF",
		7963 => x"FF",
		7964 => x"FF",
		7965 => x"FF",
		8026 => x"FF",
		8027 => x"FF",
		8028 => x"FF",
		8089 => x"FF",
		8090 => x"FF",
		8091 => x"FF",
		8152 => x"FF",
		8153 => x"FF",
		8154 => x"FF",
		8219 => x"FF",
		8220 => x"FF",
		8221 => x"FF",
		8282 => x"FF",
		8283 => x"FF",
		8284 => x"FF",
		8345 => x"FF",
		8346 => x"FF",
		8347 => x"FF",
		8408 => x"FF",
		8409 => x"FF",
		8410 => x"FF",
		8475 => x"FF",
		8476 => x"FF",
		8477 => x"FF",
		8538 => x"FF",
		8539 => x"FF",
		8540 => x"FF",
		8601 => x"FF",
		8602 => x"FF",
		8603 => x"FF",
		8664 => x"FF",
		8665 => x"FF",
		8666 => x"FF",
		8731 => x"FF",
		8732 => x"FF",
		8733 => x"FF",
		8794 => x"FF",
		8795 => x"FF",
		8796 => x"FF",
		8857 => x"FF",
		8858 => x"FF",
		8859 => x"FF",
		8920 => x"FF",
		8921 => x"FF",
		8922 => x"FF",
		8987 => x"FF",
		8988 => x"FF",
		8989 => x"FF",
		9050 => x"FF",
		9051 => x"FF",
		9052 => x"FF",
		9113 => x"FF",
		9114 => x"FF",
		9115 => x"FF",
		9176 => x"FF",
		9177 => x"FF",
		9178 => x"FF",
		9243 => x"FF",
		9244 => x"FF",
		9245 => x"FF",
		9306 => x"FF",
		9307 => x"FF",
		9308 => x"FF",
		9369 => x"FF",
		9370 => x"FF",
		9371 => x"FF",
		9432 => x"FF",
		9433 => x"FF",
		9434 => x"FF",
		9499 => x"FF",
		9500 => x"FF",
		9501 => x"FF",
		9562 => x"FF",
		9563 => x"FF",
		9564 => x"FF",
		9625 => x"FF",
		9626 => x"FF",
		9627 => x"FF",
		9688 => x"FF",
		9689 => x"FF",
		9690 => x"FF",
		9755 => x"FF",
		9756 => x"FF",
		9757 => x"FF",
		9818 => x"FF",
		9819 => x"FF",
		9820 => x"FF",
		9881 => x"FF",
		9882 => x"FF",
		9883 => x"FF",
		9944 => x"FF",
		9945 => x"FF",
		9946 => x"FF",
		10011 => x"FF",
		10012 => x"FF",
		10013 => x"FF",
		10074 => x"FF",
		10075 => x"FF",
		10076 => x"FF",
		10137 => x"FF",
		10138 => x"FF",
		10139 => x"FF",
		10200 => x"FF",
		10201 => x"FF",
		10202 => x"FF",
		10267 => x"FF",
		10268 => x"FF",
		10269 => x"FF",
		10330 => x"FF",
		10331 => x"FF",
		10332 => x"FF",
		10393 => x"FF",
		10394 => x"FF",
		10395 => x"FF",
		10456 => x"FF",
		10457 => x"FF",
		10458 => x"FF",
		10523 => x"FF",
		10524 => x"FF",
		10525 => x"FF",
		10586 => x"FF",
		10587 => x"FF",
		10588 => x"FF",
		10649 => x"FF",
		10650 => x"FF",
		10651 => x"FF",
		10712 => x"FF",
		10713 => x"FF",
		10714 => x"FF",
		10779 => x"FF",
		10780 => x"FF",
		10781 => x"FF",
		10842 => x"FF",
		10843 => x"FF",
		10844 => x"FF",
		10905 => x"FF",
		10906 => x"FF",
		10907 => x"FF",
		10968 => x"FF",
		10969 => x"FF",
		10970 => x"FF",
		11035 => x"FF",
		11036 => x"FF",
		11037 => x"FF",
		11098 => x"FF",
		11099 => x"FF",
		11100 => x"FF",
		11161 => x"FF",
		11162 => x"FF",
		11163 => x"FF",
		11224 => x"FF",
		11225 => x"FF",
		11226 => x"FF",
		11291 => x"FF",
		11292 => x"FF",
		11293 => x"FF",
		11354 => x"FF",
		11355 => x"FF",
		11356 => x"FF",
		11417 => x"FF",
		11418 => x"FF",
		11419 => x"FF",
		11480 => x"FF",
		11481 => x"FF",
		11482 => x"FF",
		11547 => x"FF",
		11548 => x"FF",
		11549 => x"FF",
		11610 => x"FF",
		11611 => x"FF",
		11612 => x"FF",
		11673 => x"FF",
		11674 => x"FF",
		11675 => x"FF",
		11736 => x"FF",
		11737 => x"FF",
		11738 => x"FF",
		11803 => x"FF",
		11804 => x"FF",
		11805 => x"FF",
		11866 => x"FF",
		11867 => x"FF",
		11868 => x"FF",
		11929 => x"FF",
		11930 => x"FF",
		11931 => x"FF",
		11992 => x"FF",
		11993 => x"FF",
		11994 => x"FF",
		12059 => x"FF",
		12060 => x"FF",
		12061 => x"FF",
		12122 => x"FF",
		12123 => x"FF",
		12124 => x"FF",
		12185 => x"FF",
		12186 => x"FF",
		12187 => x"FF",
		12248 => x"FF",
		12249 => x"FF",
		12250 => x"FF",
		12315 => x"FF",
		12316 => x"FF",
		12317 => x"FF",
		12378 => x"FF",
		12379 => x"FF",
		12380 => x"FF",
		12441 => x"FF",
		12442 => x"FF",
		12443 => x"FF",
		12504 => x"FF",
		12505 => x"FF",
		12506 => x"FF",
		12571 => x"FF",
		12572 => x"FF",
		12573 => x"FF",
		12634 => x"FF",
		12635 => x"FF",
		12636 => x"FF",
		12697 => x"FF",
		12698 => x"FF",
		12699 => x"FF",
		12760 => x"FF",
		12761 => x"FF",
		12762 => x"FF",
		12827 => x"FF",
		12828 => x"FF",
		12829 => x"FF",
		12890 => x"FF",
		12891 => x"FF",
		12892 => x"FF",
		12953 => x"FF",
		12954 => x"FF",
		12955 => x"FF",
		13016 => x"FF",
		13017 => x"FF",
		13018 => x"FF",
		13083 => x"FF",
		13084 => x"FF",
		13085 => x"FF",
		13146 => x"FF",
		13147 => x"FF",
		13148 => x"FF",
		13209 => x"FF",
		13210 => x"FF",
		13211 => x"FF",
		13272 => x"FF",
		13273 => x"FF",
		13274 => x"FF",
		13339 => x"FF",
		13340 => x"FF",
		13341 => x"FF",
		13402 => x"FF",
		13403 => x"FF",
		13404 => x"FF",
		13465 => x"FF",
		13466 => x"FF",
		13467 => x"FF",
		13528 => x"FF",
		13529 => x"FF",
		13530 => x"FF",
		13595 => x"FF",
		13596 => x"FF",
		13597 => x"FF",
		13658 => x"FF",
		13659 => x"FF",
		13660 => x"FF",
		13721 => x"FF",
		13722 => x"FF",
		13723 => x"FF",
		13784 => x"FF",
		13785 => x"FF",
		13786 => x"FF",
		13851 => x"FF",
		13852 => x"FF",
		13853 => x"FF",
		13914 => x"FF",
		13915 => x"FF",
		13916 => x"FF",
		13977 => x"FF",
		13978 => x"FF",
		13979 => x"FF",
		14040 => x"FF",
		14041 => x"FF",
		14042 => x"FF",
		14107 => x"FF",
		14108 => x"FF",
		14109 => x"FF",
		14170 => x"FF",
		14171 => x"FF",
		14172 => x"FF",
		14233 => x"FF",
		14234 => x"FF",
		14235 => x"FF",
		14296 => x"FF",
		14297 => x"FF",
		14298 => x"FF",
		14363 => x"FF",
		14364 => x"FF",
		14365 => x"FF",
		14426 => x"FF",
		14427 => x"FF",
		14428 => x"FF",
		14489 => x"FF",
		14490 => x"FF",
		14491 => x"FF",
		14552 => x"FF",
		14553 => x"FF",
		14554 => x"FF",
		14619 => x"FF",
		14620 => x"FF",
		14621 => x"FF",
		14682 => x"FF",
		14683 => x"FF",
		14684 => x"FF",
		14745 => x"FF",
		14746 => x"FF",
		14747 => x"FF",
		14808 => x"FF",
		14809 => x"FF",
		14810 => x"FF",
		14875 => x"FF",
		14876 => x"FF",
		14877 => x"FF",
		14938 => x"FF",
		14939 => x"FF",
		14940 => x"FF",
		15001 => x"FF",
		15002 => x"FF",
		15003 => x"FF",
		15064 => x"FF",
		15065 => x"FF",
		15066 => x"FF",
		15131 => x"FF",
		15132 => x"FF",
		15133 => x"FF",
		15194 => x"FF",
		15195 => x"FF",
		15196 => x"FF",
		15257 => x"FF",
		15258 => x"FF",
		15259 => x"FF",
		15320 => x"FF",
		15321 => x"FF",
		15322 => x"FF",
		15387 => x"FF",
		15388 => x"FF",
		15389 => x"FF",
		15450 => x"FF",
		15451 => x"FF",
		15452 => x"FF",
		15513 => x"FF",
		15514 => x"FF",
		15515 => x"FF",
		15576 => x"FF",
		15577 => x"FF",
		15578 => x"FF",
		15643 => x"FF",
		15644 => x"FF",
		15645 => x"FF",
		15706 => x"FF",
		15707 => x"FF",
		15708 => x"FF",
		15769 => x"FF",
		15770 => x"FF",
		15771 => x"FF",
		15832 => x"FF",
		15833 => x"FF",
		15834 => x"FF",
		15899 => x"FF",
		15900 => x"FF",
		15901 => x"FF",
		15962 => x"FF",
		15963 => x"FF",
		15964 => x"FF",
		16025 => x"FF",
		16026 => x"FF",
		16027 => x"FF",
		16088 => x"FF",
		16089 => x"FF",
		16090 => x"FF",
		16155 => x"FF",
		16156 => x"FF",
		16157 => x"FF",
		16218 => x"FF",
		16219 => x"FF",
		16220 => x"FF",
		16281 => x"FF",
		16282 => x"FF",
		16283 => x"FF",
		16344 => x"FF",
		16345 => x"FF",
		16346 => x"FF",
		16411 => x"FF",
		16412 => x"FF",
		16413 => x"FF",
		16474 => x"FF",
		16475 => x"FF",
		16476 => x"FF",
		16537 => x"FF",
		16538 => x"FF",
		16539 => x"FF",
		16600 => x"FF",
		16601 => x"FF",
		16602 => x"FF",
		16667 => x"FF",
		16668 => x"FF",
		16669 => x"FF",
		16730 => x"FF",
		16731 => x"FF",
		16732 => x"FF",
		16793 => x"FF",
		16794 => x"FF",
		16795 => x"FF",
		16856 => x"FF",
		16857 => x"FF",
		16858 => x"FF",
		16923 => x"FF",
		16924 => x"FF",
		16925 => x"FF",
		16986 => x"FF",
		16987 => x"FF",
		16988 => x"FF",
		17049 => x"FF",
		17050 => x"FF",
		17051 => x"FF",
		17112 => x"FF",
		17113 => x"FF",
		17114 => x"FF",
		17179 => x"FF",
		17180 => x"FF",
		17181 => x"FF",
		17242 => x"FF",
		17243 => x"FF",
		17244 => x"FF",
		17305 => x"FF",
		17306 => x"FF",
		17307 => x"FF",
		17368 => x"FF",
		17369 => x"FF",
		17370 => x"FF",
		17435 => x"FF",
		17436 => x"FF",
		17437 => x"FF",
		17498 => x"FF",
		17499 => x"FF",
		17500 => x"FF",
		17561 => x"FF",
		17562 => x"FF",
		17563 => x"FF",
		17624 => x"FF",
		17625 => x"FF",
		17626 => x"FF",
		17691 => x"FF",
		17692 => x"FF",
		17693 => x"FF",
		17754 => x"FF",
		17755 => x"FF",
		17756 => x"FF",
		17817 => x"FF",
		17818 => x"FF",
		17819 => x"FF",
		17880 => x"FF",
		17881 => x"FF",
		17882 => x"FF",
		17947 => x"FF",
		17948 => x"FF",
		17949 => x"FF",
		18010 => x"FF",
		18011 => x"FF",
		18012 => x"FF",
		18073 => x"FF",
		18074 => x"FF",
		18075 => x"FF",
		18136 => x"FF",
		18137 => x"FF",
		18138 => x"FF",
		18203 => x"FF",
		18204 => x"FF",
		18205 => x"FF",
		18266 => x"FF",
		18267 => x"FF",
		18268 => x"FF",
		18329 => x"FF",
		18330 => x"FF",
		18331 => x"FF",
		18392 => x"FF",
		18393 => x"FF",
		18394 => x"FF",
		18459 => x"FF",
		18460 => x"FF",
		18461 => x"FF",
		18522 => x"FF",
		18523 => x"FF",
		18524 => x"FF",
		18585 => x"FF",
		18586 => x"FF",
		18587 => x"FF",
		18648 => x"FF",
		18649 => x"FF",
		18650 => x"FF",
		18715 => x"FF",
		18716 => x"FF",
		18717 => x"FF",
		18778 => x"FF",
		18779 => x"FF",
		18780 => x"FF",
		18841 => x"FF",
		18842 => x"FF",
		18843 => x"FF",
		18904 => x"FF",
		18905 => x"FF",
		18906 => x"FF",
		18971 => x"FF",
		18972 => x"FF",
		18973 => x"FF",
		19034 => x"FF",
		19035 => x"FF",
		19036 => x"FF",
		19097 => x"FF",
		19098 => x"FF",
		19099 => x"FF",
		19160 => x"FF",
		19161 => x"FF",
		19162 => x"FF",
		19227 => x"FF",
		19228 => x"FF",
		19229 => x"FF",
		19290 => x"FF",
		19291 => x"FF",
		19292 => x"FF",
		19353 => x"FF",
		19354 => x"FF",
		19355 => x"FF",
		19416 => x"FF",
		19417 => x"FF",
		19418 => x"FF",
		19483 => x"FF",
		19484 => x"FF",
		19485 => x"FF",
		19546 => x"FF",
		19547 => x"FF",
		19548 => x"FF",
		19609 => x"FF",
		19610 => x"FF",
		19611 => x"FF",
		19672 => x"FF",
		19673 => x"FF",
		19674 => x"FF",
		19739 => x"FF",
		19740 => x"FF",
		19741 => x"FF",
		19802 => x"FF",
		19803 => x"FF",
		19804 => x"FF",
		19865 => x"FF",
		19866 => x"FF",
		19867 => x"FF",
		19928 => x"FF",
		19929 => x"FF",
		19930 => x"FF",
		19995 => x"FF",
		19996 => x"FF",
		19997 => x"FF",
		20058 => x"FF",
		20059 => x"FF",
		20060 => x"FF",
		20121 => x"FF",
		20122 => x"FF",
		20123 => x"FF",
		20184 => x"FF",
		20185 => x"FF",
		20186 => x"FF",
		20251 => x"FF",
		20252 => x"FF",
		20253 => x"FF",
		20314 => x"FF",
		20315 => x"FF",
		20316 => x"FF",
		20377 => x"FF",
		20378 => x"FF",
		20379 => x"FF",
		20440 => x"FF",
		20441 => x"FF",
		20442 => x"FF",
		20507 => x"FF",
		20508 => x"FF",
		20509 => x"FF",
		20570 => x"FF",
		20571 => x"FF",
		20572 => x"FF",
		20633 => x"FF",
		20634 => x"FF",
		20635 => x"FF",
		20696 => x"FF",
		20697 => x"FF",
		20698 => x"FF",
		20763 => x"FF",
		20764 => x"FF",
		20765 => x"FF",
		20826 => x"FF",
		20827 => x"FF",
		20828 => x"FF",
		20889 => x"FF",
		20890 => x"FF",
		20891 => x"FF",
		20952 => x"FF",
		20953 => x"FF",
		20954 => x"FF",
		21019 => x"FF",
		21020 => x"FF",
		21021 => x"FF",
		21082 => x"FF",
		21083 => x"FF",
		21084 => x"FF",
		21145 => x"FF",
		21146 => x"FF",
		21147 => x"FF",
		21208 => x"FF",
		21209 => x"FF",
		21210 => x"FF",
		21275 => x"FF",
		21276 => x"FF",
		21277 => x"FF",
		21338 => x"FF",
		21339 => x"FF",
		21340 => x"FF",
		21401 => x"FF",
		21402 => x"FF",
		21403 => x"FF",
		21464 => x"FF",
		21465 => x"FF",
		21466 => x"FF",
		21531 => x"FF",
		21532 => x"FF",
		21533 => x"FF",
		21594 => x"FF",
		21595 => x"FF",
		21596 => x"FF",
		21657 => x"FF",
		21658 => x"FF",
		21659 => x"FF",
		21720 => x"FF",
		21721 => x"FF",
		21722 => x"FF",
		21787 => x"FF",
		21788 => x"FF",
		21789 => x"FF",
		21850 => x"FF",
		21851 => x"FF",
		21852 => x"FF",
		21913 => x"FF",
		21914 => x"FF",
		21915 => x"FF",
		21976 => x"FF",
		21977 => x"FF",
		21978 => x"FF",
		22043 => x"FF",
		22044 => x"FF",
		22045 => x"FF",
		22106 => x"FF",
		22107 => x"FF",
		22108 => x"FF",
		22169 => x"FF",
		22170 => x"FF",
		22171 => x"FF",
		22232 => x"FF",
		22233 => x"FF",
		22234 => x"FF",
		22299 => x"FF",
		22300 => x"FF",
		22301 => x"FF",
		22362 => x"FF",
		22363 => x"FF",
		22364 => x"FF",
		22425 => x"FF",
		22426 => x"FF",
		22427 => x"FF",
		22488 => x"FF",
		22489 => x"FF",
		22490 => x"FF",
		22555 => x"FF",
		22556 => x"FF",
		22557 => x"FF",
		22618 => x"FF",
		22619 => x"FF",
		22620 => x"FF",
		22681 => x"FF",
		22682 => x"FF",
		22683 => x"FF",
		22744 => x"FF",
		22745 => x"FF",
		22746 => x"FF",
		22811 => x"FF",
		22812 => x"FF",
		22813 => x"FF",
		22874 => x"FF",
		22875 => x"FF",
		22876 => x"FF",
		22937 => x"FF",
		22938 => x"FF",
		22939 => x"FF",
		23000 => x"FF",
		23001 => x"FF",
		23002 => x"FF",
		23067 => x"FF",
		23068 => x"FF",
		23069 => x"FF",
		23070 => x"FF",
		23071 => x"FF",
		23072 => x"FF",
		23073 => x"FF",
		23074 => x"FF",
		23075 => x"FF",
		23076 => x"FF",
		23077 => x"FF",
		23078 => x"FF",
		23079 => x"FF",
		23080 => x"FF",
		23081 => x"FF",
		23082 => x"FF",
		23083 => x"FF",
		23084 => x"FF",
		23085 => x"FF",
		23086 => x"FF",
		23087 => x"FF",
		23088 => x"FF",
		23089 => x"FF",
		23090 => x"FF",
		23091 => x"FF",
		23092 => x"FF",
		23093 => x"FF",
		23094 => x"FF",
		23095 => x"FF",
		23096 => x"FF",
		23097 => x"FF",
		23098 => x"FF",
		23099 => x"FF",
		23100 => x"FF",
		23101 => x"FF",
		23102 => x"FF",
		23103 => x"FF",
		23104 => x"FF",
		23105 => x"FF",
		23106 => x"FF",
		23107 => x"FF",
		23108 => x"FF",
		23109 => x"FF",
		23110 => x"FF",
		23111 => x"FF",
		23112 => x"FF",
		23113 => x"FF",
		23114 => x"FF",
		23115 => x"FF",
		23116 => x"FF",
		23117 => x"FF",
		23118 => x"FF",
		23119 => x"FF",
		23120 => x"FF",
		23121 => x"FF",
		23122 => x"FF",
		23123 => x"FF",
		23124 => x"FF",
		23125 => x"FF",
		23126 => x"FF",
		23127 => x"FF",
		23128 => x"FF",
		23129 => x"FF",
		23130 => x"FF",
		23131 => x"FF",
		23132 => x"FF",
		23133 => x"FF",
		23134 => x"FF",
		23135 => x"FF",
		23136 => x"FF",
		23137 => x"FF",
		23138 => x"FF",
		23139 => x"FF",
		23140 => x"FF",
		23141 => x"FF",
		23142 => x"FF",
		23143 => x"FF",
		23144 => x"FF",
		23145 => x"FF",
		23146 => x"FF",
		23147 => x"FF",
		23148 => x"FF",
		23149 => x"FF",
		23150 => x"FF",
		23151 => x"FF",
		23152 => x"FF",
		23153 => x"FF",
		23154 => x"FF",
		23155 => x"FF",
		23156 => x"FF",
		23157 => x"FF",
		23158 => x"FF",
		23159 => x"FF",
		23160 => x"FF",
		23161 => x"FF",
		23162 => x"FF",
		23163 => x"FF",
		23164 => x"FF",
		23165 => x"FF",
		23166 => x"FF",
		23167 => x"FF",
		23168 => x"FF",
		23169 => x"FF",
		23170 => x"FF",
		23171 => x"FF",
		23172 => x"FF",
		23173 => x"FF",
		23174 => x"FF",
		23175 => x"FF",
		23176 => x"FF",
		23177 => x"FF",
		23178 => x"FF",
		23179 => x"FF",
		23180 => x"FF",
		23181 => x"FF",
		23182 => x"FF",
		23183 => x"FF",
		23184 => x"FF",
		23185 => x"FF",
		23186 => x"FF",
		23187 => x"FF",
		23188 => x"FF",
		23189 => x"FF",
		23190 => x"FF",
		23191 => x"FF",
		23192 => x"FF",
		23193 => x"FF",
		23194 => x"FF",
		23195 => x"FF",
		23196 => x"FF",
		23197 => x"FF",
		23198 => x"FF",
		23199 => x"FF",
		23200 => x"FF",
		23201 => x"FF",
		23202 => x"FF",
		23203 => x"FF",
		23204 => x"FF",
		23205 => x"FF",
		23206 => x"FF",
		23207 => x"FF",
		23208 => x"FF",
		23209 => x"FF",
		23210 => x"FF",
		23211 => x"FF",
		23212 => x"FF",
		23213 => x"FF",
		23214 => x"FF",
		23215 => x"FF",
		23216 => x"FF",
		23217 => x"FF",
		23218 => x"FF",
		23219 => x"FF",
		23220 => x"FF",
		23221 => x"FF",
		23222 => x"FF",
		23223 => x"FF",
		23224 => x"FF",
		23225 => x"FF",
		23226 => x"FF",
		23227 => x"FF",
		23228 => x"FF",
		23229 => x"FF",
		23230 => x"FF",
		23231 => x"FF",
		23232 => x"FF",
		23233 => x"FF",
		23234 => x"FF",
		23235 => x"FF",
		23236 => x"FF",
		23237 => x"FF",
		23238 => x"FF",
		23239 => x"FF",
		23240 => x"FF",
		23241 => x"FF",
		23242 => x"FF",
		23243 => x"FF",
		23244 => x"FF",
		23245 => x"FF",
		23246 => x"FF",
		23247 => x"FF",
		23248 => x"FF",
		23249 => x"FF",
		23250 => x"FF",
		23251 => x"FF",
		23252 => x"FF",
		23253 => x"FF",
		23254 => x"FF",
		23255 => x"FF",
		23256 => x"FF",
		23257 => x"FF",
		23258 => x"FF",
		23323 => x"FF",
		23324 => x"FF",
		23325 => x"FF",
		23326 => x"FF",
		23327 => x"FF",
		23328 => x"FF",
		23329 => x"FF",
		23330 => x"FF",
		23331 => x"FF",
		23332 => x"FF",
		23333 => x"FF",
		23334 => x"FF",
		23335 => x"FF",
		23336 => x"FF",
		23337 => x"FF",
		23338 => x"FF",
		23339 => x"FF",
		23340 => x"FF",
		23341 => x"FF",
		23342 => x"FF",
		23343 => x"FF",
		23344 => x"FF",
		23345 => x"FF",
		23346 => x"FF",
		23347 => x"FF",
		23348 => x"FF",
		23349 => x"FF",
		23350 => x"FF",
		23351 => x"FF",
		23352 => x"FF",
		23353 => x"FF",
		23354 => x"FF",
		23355 => x"FF",
		23356 => x"FF",
		23357 => x"FF",
		23358 => x"FF",
		23359 => x"FF",
		23360 => x"FF",
		23361 => x"FF",
		23362 => x"FF",
		23363 => x"FF",
		23364 => x"FF",
		23365 => x"FF",
		23366 => x"FF",
		23367 => x"FF",
		23368 => x"FF",
		23369 => x"FF",
		23370 => x"FF",
		23371 => x"FF",
		23372 => x"FF",
		23373 => x"FF",
		23374 => x"FF",
		23375 => x"FF",
		23376 => x"FF",
		23377 => x"FF",
		23378 => x"FF",
		23379 => x"FF",
		23380 => x"FF",
		23381 => x"FF",
		23382 => x"FF",
		23383 => x"FF",
		23384 => x"FF",
		23385 => x"FF",
		23386 => x"FF",
		23387 => x"FF",
		23388 => x"FF",
		23389 => x"FF",
		23390 => x"FF",
		23391 => x"FF",
		23392 => x"FF",
		23393 => x"FF",
		23394 => x"FF",
		23395 => x"FF",
		23396 => x"FF",
		23397 => x"FF",
		23398 => x"FF",
		23399 => x"FF",
		23400 => x"FF",
		23401 => x"FF",
		23402 => x"FF",
		23403 => x"FF",
		23404 => x"FF",
		23405 => x"FF",
		23406 => x"FF",
		23407 => x"FF",
		23408 => x"FF",
		23409 => x"FF",
		23410 => x"FF",
		23411 => x"FF",
		23412 => x"FF",
		23413 => x"FF",
		23414 => x"FF",
		23415 => x"FF",
		23416 => x"FF",
		23417 => x"FF",
		23418 => x"FF",
		23419 => x"FF",
		23420 => x"FF",
		23421 => x"FF",
		23422 => x"FF",
		23423 => x"FF",
		23424 => x"FF",
		23425 => x"FF",
		23426 => x"FF",
		23427 => x"FF",
		23428 => x"FF",
		23429 => x"FF",
		23430 => x"FF",
		23431 => x"FF",
		23432 => x"FF",
		23433 => x"FF",
		23434 => x"FF",
		23435 => x"FF",
		23436 => x"FF",
		23437 => x"FF",
		23438 => x"FF",
		23439 => x"FF",
		23440 => x"FF",
		23441 => x"FF",
		23442 => x"FF",
		23443 => x"FF",
		23444 => x"FF",
		23445 => x"FF",
		23446 => x"FF",
		23447 => x"FF",
		23448 => x"FF",
		23449 => x"FF",
		23450 => x"FF",
		23451 => x"FF",
		23452 => x"FF",
		23453 => x"FF",
		23454 => x"FF",
		23455 => x"FF",
		23456 => x"FF",
		23457 => x"FF",
		23458 => x"FF",
		23459 => x"FF",
		23460 => x"FF",
		23461 => x"FF",
		23462 => x"FF",
		23463 => x"FF",
		23464 => x"FF",
		23465 => x"FF",
		23466 => x"FF",
		23467 => x"FF",
		23468 => x"FF",
		23469 => x"FF",
		23470 => x"FF",
		23471 => x"FF",
		23472 => x"FF",
		23473 => x"FF",
		23474 => x"FF",
		23475 => x"FF",
		23476 => x"FF",
		23477 => x"FF",
		23478 => x"FF",
		23479 => x"FF",
		23480 => x"FF",
		23481 => x"FF",
		23482 => x"FF",
		23483 => x"FF",
		23484 => x"FF",
		23485 => x"FF",
		23486 => x"FF",
		23487 => x"FF",
		23488 => x"FF",
		23489 => x"FF",
		23490 => x"FF",
		23491 => x"FF",
		23492 => x"FF",
		23493 => x"FF",
		23494 => x"FF",
		23495 => x"FF",
		23496 => x"FF",
		23497 => x"FF",
		23498 => x"FF",
		23499 => x"FF",
		23500 => x"FF",
		23501 => x"FF",
		23502 => x"FF",
		23503 => x"FF",
		23504 => x"FF",
		23505 => x"FF",
		23506 => x"FF",
		23507 => x"FF",
		23508 => x"FF",
		23509 => x"FF",
		23510 => x"FF",
		23511 => x"FF",
		23512 => x"FF",
		23513 => x"FF",
		23514 => x"FF",
		23579 => x"FF",
		23580 => x"FF",
		23581 => x"FF",
		23582 => x"FF",
		23583 => x"FF",
		23584 => x"FF",
		23585 => x"FF",
		23586 => x"FF",
		23587 => x"FF",
		23588 => x"FF",
		23589 => x"FF",
		23590 => x"FF",
		23591 => x"FF",
		23592 => x"FF",
		23593 => x"FF",
		23594 => x"FF",
		23595 => x"FF",
		23596 => x"FF",
		23597 => x"FF",
		23598 => x"FF",
		23599 => x"FF",
		23600 => x"FF",
		23601 => x"FF",
		23602 => x"FF",
		23603 => x"FF",
		23604 => x"FF",
		23605 => x"FF",
		23606 => x"FF",
		23607 => x"FF",
		23608 => x"FF",
		23609 => x"FF",
		23610 => x"FF",
		23611 => x"FF",
		23612 => x"FF",
		23613 => x"FF",
		23614 => x"FF",
		23615 => x"FF",
		23616 => x"FF",
		23617 => x"FF",
		23618 => x"FF",
		23619 => x"FF",
		23620 => x"FF",
		23621 => x"FF",
		23622 => x"FF",
		23623 => x"FF",
		23624 => x"FF",
		23625 => x"FF",
		23626 => x"FF",
		23627 => x"FF",
		23628 => x"FF",
		23629 => x"FF",
		23630 => x"FF",
		23631 => x"FF",
		23632 => x"FF",
		23633 => x"FF",
		23634 => x"FF",
		23635 => x"FF",
		23636 => x"FF",
		23637 => x"FF",
		23638 => x"FF",
		23639 => x"FF",
		23640 => x"FF",
		23641 => x"FF",
		23642 => x"FF",
		23643 => x"FF",
		23644 => x"FF",
		23645 => x"FF",
		23646 => x"FF",
		23647 => x"FF",
		23648 => x"FF",
		23649 => x"FF",
		23650 => x"FF",
		23651 => x"FF",
		23652 => x"FF",
		23653 => x"FF",
		23654 => x"FF",
		23655 => x"FF",
		23656 => x"FF",
		23657 => x"FF",
		23658 => x"FF",
		23659 => x"FF",
		23660 => x"FF",
		23661 => x"FF",
		23662 => x"FF",
		23663 => x"FF",
		23664 => x"FF",
		23665 => x"FF",
		23666 => x"FF",
		23667 => x"FF",
		23668 => x"FF",
		23669 => x"FF",
		23670 => x"FF",
		23671 => x"FF",
		23672 => x"FF",
		23673 => x"FF",
		23674 => x"FF",
		23675 => x"FF",
		23676 => x"FF",
		23677 => x"FF",
		23678 => x"FF",
		23679 => x"FF",
		23680 => x"FF",
		23681 => x"FF",
		23682 => x"FF",
		23683 => x"FF",
		23684 => x"FF",
		23685 => x"FF",
		23686 => x"FF",
		23687 => x"FF",
		23688 => x"FF",
		23689 => x"FF",
		23690 => x"FF",
		23691 => x"FF",
		23692 => x"FF",
		23693 => x"FF",
		23694 => x"FF",
		23695 => x"FF",
		23696 => x"FF",
		23697 => x"FF",
		23698 => x"FF",
		23699 => x"FF",
		23700 => x"FF",
		23701 => x"FF",
		23702 => x"FF",
		23703 => x"FF",
		23704 => x"FF",
		23705 => x"FF",
		23706 => x"FF",
		23707 => x"FF",
		23708 => x"FF",
		23709 => x"FF",
		23710 => x"FF",
		23711 => x"FF",
		23712 => x"FF",
		23713 => x"FF",
		23714 => x"FF",
		23715 => x"FF",
		23716 => x"FF",
		23717 => x"FF",
		23718 => x"FF",
		23719 => x"FF",
		23720 => x"FF",
		23721 => x"FF",
		23722 => x"FF",
		23723 => x"FF",
		23724 => x"FF",
		23725 => x"FF",
		23726 => x"FF",
		23727 => x"FF",
		23728 => x"FF",
		23729 => x"FF",
		23730 => x"FF",
		23731 => x"FF",
		23732 => x"FF",
		23733 => x"FF",
		23734 => x"FF",
		23735 => x"FF",
		23736 => x"FF",
		23737 => x"FF",
		23738 => x"FF",
		23739 => x"FF",
		23740 => x"FF",
		23741 => x"FF",
		23742 => x"FF",
		23743 => x"FF",
		23744 => x"FF",
		23745 => x"FF",
		23746 => x"FF",
		23747 => x"FF",
		23748 => x"FF",
		23749 => x"FF",
		23750 => x"FF",
		23751 => x"FF",
		23752 => x"FF",
		23753 => x"FF",
		23754 => x"FF",
		23755 => x"FF",
		23756 => x"FF",
		23757 => x"FF",
		23758 => x"FF",
		23759 => x"FF",
		23760 => x"FF",
		23761 => x"FF",
		23762 => x"FF",
		23763 => x"FF",
		23764 => x"FF",
		23765 => x"FF",
		23766 => x"FF",
		23767 => x"FF",
		23768 => x"FF",
		23769 => x"FF",
		23770 => x"FF",
		23835 => x"FF",
		23836 => x"FF",
		23837 => x"FF",
		23898 => x"FF",
		23899 => x"FF",
		23900 => x"FF",
		23961 => x"FF",
		23962 => x"FF",
		23963 => x"FF",
		24024 => x"FF",
		24025 => x"FF",
		24026 => x"FF",
		24091 => x"FF",
		24092 => x"FF",
		24093 => x"FF",
		24154 => x"FF",
		24155 => x"FF",
		24156 => x"FF",
		24217 => x"FF",
		24218 => x"FF",
		24219 => x"FF",
		24280 => x"FF",
		24281 => x"FF",
		24282 => x"FF",
		24347 => x"FF",
		24348 => x"FF",
		24349 => x"FF",
		24410 => x"FF",
		24411 => x"FF",
		24412 => x"FF",
		24473 => x"FF",
		24474 => x"FF",
		24475 => x"FF",
		24536 => x"FF",
		24537 => x"FF",
		24538 => x"FF",
		24603 => x"FF",
		24604 => x"FF",
		24605 => x"FF",
		24666 => x"FF",
		24667 => x"FF",
		24668 => x"FF",
		24729 => x"FF",
		24730 => x"FF",
		24731 => x"FF",
		24792 => x"FF",
		24793 => x"FF",
		24794 => x"FF",
		24859 => x"FF",
		24860 => x"FF",
		24861 => x"FF",
		24922 => x"FF",
		24923 => x"FF",
		24924 => x"FF",
		24985 => x"FF",
		24986 => x"FF",
		24987 => x"FF",
		25048 => x"FF",
		25049 => x"FF",
		25050 => x"FF",
		25115 => x"FF",
		25116 => x"FF",
		25117 => x"FF",
		25178 => x"FF",
		25179 => x"FF",
		25180 => x"FF",
		25241 => x"FF",
		25242 => x"FF",
		25243 => x"FF",
		25304 => x"FF",
		25305 => x"FF",
		25306 => x"FF",
		25371 => x"FF",
		25372 => x"FF",
		25373 => x"FF",
		25434 => x"FF",
		25435 => x"FF",
		25436 => x"FF",
		25497 => x"FF",
		25498 => x"FF",
		25499 => x"FF",
		25560 => x"FF",
		25561 => x"FF",
		25562 => x"FF",
		25627 => x"FF",
		25628 => x"FF",
		25629 => x"FF",
		25690 => x"FF",
		25691 => x"FF",
		25692 => x"FF",
		25753 => x"FF",
		25754 => x"FF",
		25755 => x"FF",
		25816 => x"FF",
		25817 => x"FF",
		25818 => x"FF",
		25883 => x"FF",
		25884 => x"FF",
		25885 => x"FF",
		25946 => x"FF",
		25947 => x"FF",
		25948 => x"FF",
		26009 => x"FF",
		26010 => x"FF",
		26011 => x"FF",
		26072 => x"FF",
		26073 => x"FF",
		26074 => x"FF",
		26139 => x"FF",
		26140 => x"FF",
		26141 => x"FF",
		26202 => x"FF",
		26203 => x"FF",
		26204 => x"FF",
		26265 => x"FF",
		26266 => x"FF",
		26267 => x"FF",
		26328 => x"FF",
		26329 => x"FF",
		26330 => x"FF",
		26395 => x"FF",
		26396 => x"FF",
		26397 => x"FF",
		26458 => x"FF",
		26459 => x"FF",
		26460 => x"FF",
		26521 => x"FF",
		26522 => x"FF",
		26523 => x"FF",
		26584 => x"FF",
		26585 => x"FF",
		26586 => x"FF",
		26651 => x"FF",
		26652 => x"FF",
		26653 => x"FF",
		26714 => x"FF",
		26715 => x"FF",
		26716 => x"FF",
		26777 => x"FF",
		26778 => x"FF",
		26779 => x"FF",
		26840 => x"FF",
		26841 => x"FF",
		26842 => x"FF",
		26907 => x"FF",
		26908 => x"FF",
		26909 => x"FF",
		26970 => x"FF",
		26971 => x"FF",
		26972 => x"FF",
		27033 => x"FF",
		27034 => x"FF",
		27035 => x"FF",
		27096 => x"FF",
		27097 => x"FF",
		27098 => x"FF",
		27163 => x"FF",
		27164 => x"FF",
		27165 => x"FF",
		27226 => x"FF",
		27227 => x"FF",
		27228 => x"FF",
		27289 => x"FF",
		27290 => x"FF",
		27291 => x"FF",
		27352 => x"FF",
		27353 => x"FF",
		27354 => x"FF",
		27419 => x"FF",
		27420 => x"FF",
		27421 => x"FF",
		27482 => x"FF",
		27483 => x"FF",
		27484 => x"FF",
		27545 => x"FF",
		27546 => x"FF",
		27547 => x"FF",
		27608 => x"FF",
		27609 => x"FF",
		27610 => x"FF",
		27675 => x"FF",
		27676 => x"FF",
		27677 => x"FF",
		27738 => x"FF",
		27739 => x"FF",
		27740 => x"FF",
		27801 => x"FF",
		27802 => x"FF",
		27803 => x"FF",
		27864 => x"FF",
		27865 => x"FF",
		27866 => x"FF",
		27931 => x"FF",
		27932 => x"FF",
		27933 => x"FF",
		27994 => x"FF",
		27995 => x"FF",
		27996 => x"FF",
		28057 => x"FF",
		28058 => x"FF",
		28059 => x"FF",
		28120 => x"FF",
		28121 => x"FF",
		28122 => x"FF",
		28187 => x"FF",
		28188 => x"FF",
		28189 => x"FF",
		28250 => x"FF",
		28251 => x"FF",
		28252 => x"FF",
		28313 => x"FF",
		28314 => x"FF",
		28315 => x"FF",
		28376 => x"FF",
		28377 => x"FF",
		28378 => x"FF",
		28443 => x"FF",
		28444 => x"FF",
		28445 => x"FF",
		28506 => x"FF",
		28507 => x"FF",
		28508 => x"FF",
		28569 => x"FF",
		28570 => x"FF",
		28571 => x"FF",
		28632 => x"FF",
		28633 => x"FF",
		28634 => x"FF",
		28699 => x"FF",
		28700 => x"FF",
		28701 => x"FF",
		28762 => x"FF",
		28763 => x"FF",
		28764 => x"FF",
		28825 => x"FF",
		28826 => x"FF",
		28827 => x"FF",
		28888 => x"FF",
		28889 => x"FF",
		28890 => x"FF",
		28955 => x"FF",
		28956 => x"FF",
		28957 => x"FF",
		29018 => x"FF",
		29019 => x"FF",
		29020 => x"FF",
		29081 => x"FF",
		29082 => x"FF",
		29083 => x"FF",
		29144 => x"FF",
		29145 => x"FF",
		29146 => x"FF",
		29211 => x"FF",
		29212 => x"FF",
		29213 => x"FF",
		29274 => x"FF",
		29275 => x"FF",
		29276 => x"FF",
		29337 => x"FF",
		29338 => x"FF",
		29339 => x"FF",
		29400 => x"FF",
		29401 => x"FF",
		29402 => x"FF",
		29467 => x"FF",
		29468 => x"FF",
		29469 => x"FF",
		29530 => x"FF",
		29531 => x"FF",
		29532 => x"FF",
		29593 => x"FF",
		29594 => x"FF",
		29595 => x"FF",
		29656 => x"FF",
		29657 => x"FF",
		29658 => x"FF",
		29723 => x"FF",
		29724 => x"FF",
		29725 => x"FF",
		29786 => x"FF",
		29787 => x"FF",
		29788 => x"FF",
		29849 => x"FF",
		29850 => x"FF",
		29851 => x"FF",
		29912 => x"FF",
		29913 => x"FF",
		29914 => x"FF",
		29979 => x"FF",
		29980 => x"FF",
		29981 => x"FF",
		30042 => x"FF",
		30043 => x"FF",
		30044 => x"FF",
		30105 => x"FF",
		30106 => x"FF",
		30107 => x"FF",
		30168 => x"FF",
		30169 => x"FF",
		30170 => x"FF",
		30235 => x"FF",
		30236 => x"FF",
		30237 => x"FF",
		30298 => x"FF",
		30299 => x"FF",
		30300 => x"FF",
		30361 => x"FF",
		30362 => x"FF",
		30363 => x"FF",
		30424 => x"FF",
		30425 => x"FF",
		30426 => x"FF",
		30491 => x"FF",
		30492 => x"FF",
		30493 => x"FF",
		30554 => x"FF",
		30555 => x"FF",
		30556 => x"FF",
		30617 => x"FF",
		30618 => x"FF",
		30619 => x"FF",
		30680 => x"FF",
		30681 => x"FF",
		30682 => x"FF",
		30747 => x"FF",
		30748 => x"FF",
		30749 => x"FF",
		30810 => x"FF",
		30811 => x"FF",
		30812 => x"FF",
		30873 => x"FF",
		30874 => x"FF",
		30875 => x"FF",
		30936 => x"FF",
		30937 => x"FF",
		30938 => x"FF",
		31003 => x"FF",
		31004 => x"FF",
		31005 => x"FF",
		31066 => x"FF",
		31067 => x"FF",
		31068 => x"FF",
		31129 => x"FF",
		31130 => x"FF",
		31131 => x"FF",
		31192 => x"FF",
		31193 => x"FF",
		31194 => x"FF",
		31259 => x"FF",
		31260 => x"FF",
		31261 => x"FF",
		31322 => x"FF",
		31323 => x"FF",
		31324 => x"FF",
		31385 => x"FF",
		31386 => x"FF",
		31387 => x"FF",
		31448 => x"FF",
		31449 => x"FF",
		31450 => x"FF",
		31515 => x"FF",
		31516 => x"FF",
		31517 => x"FF",
		31578 => x"FF",
		31579 => x"FF",
		31580 => x"FF",
		31641 => x"FF",
		31642 => x"FF",
		31643 => x"FF",
		31704 => x"FF",
		31705 => x"FF",
		31706 => x"FF",
		31771 => x"FF",
		31772 => x"FF",
		31773 => x"FF",
		31834 => x"FF",
		31835 => x"FF",
		31836 => x"FF",
		31897 => x"FF",
		31898 => x"FF",
		31899 => x"FF",
		31960 => x"FF",
		31961 => x"FF",
		31962 => x"FF",
		32027 => x"FF",
		32028 => x"FF",
		32029 => x"FF",
		32090 => x"FF",
		32091 => x"FF",
		32092 => x"FF",
		32153 => x"FF",
		32154 => x"FF",
		32155 => x"FF",
		32216 => x"FF",
		32217 => x"FF",
		32218 => x"FF",
		32283 => x"FF",
		32284 => x"FF",
		32285 => x"FF",
		32346 => x"FF",
		32347 => x"FF",
		32348 => x"FF",
		32409 => x"FF",
		32410 => x"FF",
		32411 => x"FF",
		32472 => x"FF",
		32473 => x"FF",
		32474 => x"FF",
		32539 => x"FF",
		32540 => x"FF",
		32541 => x"FF",
		32602 => x"FF",
		32603 => x"FF",
		32604 => x"FF",
		32665 => x"FF",
		32666 => x"FF",
		32667 => x"FF",
		32728 => x"FF",
		32729 => x"FF",
		32730 => x"FF",
		32795 => x"FF",
		32796 => x"FF",
		32797 => x"FF",
		32858 => x"FF",
		32859 => x"FF",
		32860 => x"FF",
		32921 => x"FF",
		32922 => x"FF",
		32923 => x"FF",
		32984 => x"FF",
		32985 => x"FF",
		32986 => x"FF",
		33051 => x"FF",
		33052 => x"FF",
		33053 => x"FF",
		33114 => x"FF",
		33115 => x"FF",
		33116 => x"FF",
		33177 => x"FF",
		33178 => x"FF",
		33179 => x"FF",
		33240 => x"FF",
		33241 => x"FF",
		33242 => x"FF",
		33307 => x"FF",
		33308 => x"FF",
		33309 => x"FF",
		33370 => x"FF",
		33371 => x"FF",
		33372 => x"FF",
		33433 => x"FF",
		33434 => x"FF",
		33435 => x"FF",
		33496 => x"FF",
		33497 => x"FF",
		33498 => x"FF",
		33563 => x"FF",
		33564 => x"FF",
		33565 => x"FF",
		33626 => x"FF",
		33627 => x"FF",
		33628 => x"FF",
		33689 => x"FF",
		33690 => x"FF",
		33691 => x"FF",
		33752 => x"FF",
		33753 => x"FF",
		33754 => x"FF",
		33819 => x"FF",
		33820 => x"FF",
		33821 => x"FF",
		33882 => x"FF",
		33883 => x"FF",
		33884 => x"FF",
		33945 => x"FF",
		33946 => x"FF",
		33947 => x"FF",
		34008 => x"FF",
		34009 => x"FF",
		34010 => x"FF",
		34075 => x"FF",
		34076 => x"FF",
		34077 => x"FF",
		34138 => x"FF",
		34139 => x"FF",
		34140 => x"FF",
		34201 => x"FF",
		34202 => x"FF",
		34203 => x"FF",
		34264 => x"FF",
		34265 => x"FF",
		34266 => x"FF",
		34331 => x"FF",
		34332 => x"FF",
		34333 => x"FF",
		34394 => x"FF",
		34395 => x"FF",
		34396 => x"FF",
		34457 => x"FF",
		34458 => x"FF",
		34459 => x"FF",
		34520 => x"FF",
		34521 => x"FF",
		34522 => x"FF",
		34587 => x"FF",
		34588 => x"FF",
		34589 => x"FF",
		34650 => x"FF",
		34651 => x"FF",
		34652 => x"FF",
		34713 => x"FF",
		34714 => x"FF",
		34715 => x"FF",
		34776 => x"FF",
		34777 => x"FF",
		34778 => x"FF",
		34843 => x"FF",
		34844 => x"FF",
		34845 => x"FF",
		34906 => x"FF",
		34907 => x"FF",
		34908 => x"FF",
		34969 => x"FF",
		34970 => x"FF",
		34971 => x"FF",
		35032 => x"FF",
		35033 => x"FF",
		35034 => x"FF",
		35099 => x"FF",
		35100 => x"FF",
		35101 => x"FF",
		35162 => x"FF",
		35163 => x"FF",
		35164 => x"FF",
		35225 => x"FF",
		35226 => x"FF",
		35227 => x"FF",
		35288 => x"FF",
		35289 => x"FF",
		35290 => x"FF",
		35355 => x"FF",
		35356 => x"FF",
		35357 => x"FF",
		35418 => x"FF",
		35419 => x"FF",
		35420 => x"FF",
		35481 => x"FF",
		35482 => x"FF",
		35483 => x"FF",
		35544 => x"FF",
		35545 => x"FF",
		35546 => x"FF",
		35611 => x"FF",
		35612 => x"FF",
		35613 => x"FF",
		35674 => x"FF",
		35675 => x"FF",
		35676 => x"FF",
		35737 => x"FF",
		35738 => x"FF",
		35739 => x"FF",
		35800 => x"FF",
		35801 => x"FF",
		35802 => x"FF",
		35867 => x"FF",
		35868 => x"FF",
		35869 => x"FF",
		35930 => x"FF",
		35931 => x"FF",
		35932 => x"FF",
		35993 => x"FF",
		35994 => x"FF",
		35995 => x"FF",
		36056 => x"FF",
		36057 => x"FF",
		36058 => x"FF",
		36123 => x"FF",
		36124 => x"FF",
		36125 => x"FF",
		36186 => x"FF",
		36187 => x"FF",
		36188 => x"FF",
		36249 => x"FF",
		36250 => x"FF",
		36251 => x"FF",
		36312 => x"FF",
		36313 => x"FF",
		36314 => x"FF",
		36379 => x"FF",
		36380 => x"FF",
		36381 => x"FF",
		36442 => x"FF",
		36443 => x"FF",
		36444 => x"FF",
		36505 => x"FF",
		36506 => x"FF",
		36507 => x"FF",
		36568 => x"FF",
		36569 => x"FF",
		36570 => x"FF",
		36635 => x"FF",
		36636 => x"FF",
		36637 => x"FF",
		36698 => x"FF",
		36699 => x"FF",
		36700 => x"FF",
		36761 => x"FF",
		36762 => x"FF",
		36763 => x"FF",
		36824 => x"FF",
		36825 => x"FF",
		36826 => x"FF",
		36891 => x"FF",
		36892 => x"FF",
		36893 => x"FF",
		36954 => x"FF",
		36955 => x"FF",
		36956 => x"FF",
		37017 => x"FF",
		37018 => x"FF",
		37019 => x"FF",
		37080 => x"FF",
		37081 => x"FF",
		37082 => x"FF",
		37147 => x"FF",
		37148 => x"FF",
		37149 => x"FF",
		37210 => x"FF",
		37211 => x"FF",
		37212 => x"FF",
		37273 => x"FF",
		37274 => x"FF",
		37275 => x"FF",
		37336 => x"FF",
		37337 => x"FF",
		37338 => x"FF",
		37403 => x"FF",
		37404 => x"FF",
		37405 => x"FF",
		37466 => x"FF",
		37467 => x"FF",
		37468 => x"FF",
		37529 => x"FF",
		37530 => x"FF",
		37531 => x"FF",
		37592 => x"FF",
		37593 => x"FF",
		37594 => x"FF",
		37659 => x"FF",
		37660 => x"FF",
		37661 => x"FF",
		37722 => x"FF",
		37723 => x"FF",
		37724 => x"FF",
		37785 => x"FF",
		37786 => x"FF",
		37787 => x"FF",
		37848 => x"FF",
		37849 => x"FF",
		37850 => x"FF",
		37915 => x"FF",
		37916 => x"FF",
		37917 => x"FF",
		37978 => x"FF",
		37979 => x"FF",
		37980 => x"FF",
		38041 => x"FF",
		38042 => x"FF",
		38043 => x"FF",
		38104 => x"FF",
		38105 => x"FF",
		38106 => x"FF",
		38171 => x"FF",
		38172 => x"FF",
		38173 => x"FF",
		38234 => x"FF",
		38235 => x"FF",
		38236 => x"FF",
		38297 => x"FF",
		38298 => x"FF",
		38299 => x"FF",
		38360 => x"FF",
		38361 => x"FF",
		38362 => x"FF",
		38427 => x"FF",
		38428 => x"FF",
		38429 => x"FF",
		38490 => x"FF",
		38491 => x"FF",
		38492 => x"FF",
		38553 => x"FF",
		38554 => x"FF",
		38555 => x"FF",
		38616 => x"FF",
		38617 => x"FF",
		38618 => x"FF",
		38683 => x"FF",
		38684 => x"FF",
		38685 => x"FF",
		38746 => x"FF",
		38747 => x"FF",
		38748 => x"FF",
		38809 => x"FF",
		38810 => x"FF",
		38811 => x"FF",
		38872 => x"FF",
		38873 => x"FF",
		38874 => x"FF",
		38939 => x"FF",
		38940 => x"FF",
		38941 => x"FF",
		39002 => x"FF",
		39003 => x"FF",
		39004 => x"FF",
		39065 => x"FF",
		39066 => x"FF",
		39067 => x"FF",
		39128 => x"FF",
		39129 => x"FF",
		39130 => x"FF",
		39195 => x"FF",
		39196 => x"FF",
		39197 => x"FF",
		39198 => x"FF",
		39199 => x"FF",
		39200 => x"FF",
		39201 => x"FF",
		39202 => x"FF",
		39203 => x"FF",
		39204 => x"FF",
		39205 => x"FF",
		39206 => x"FF",
		39207 => x"FF",
		39208 => x"FF",
		39209 => x"FF",
		39210 => x"FF",
		39211 => x"FF",
		39212 => x"FF",
		39213 => x"FF",
		39214 => x"FF",
		39215 => x"FF",
		39216 => x"FF",
		39217 => x"FF",
		39218 => x"FF",
		39219 => x"FF",
		39220 => x"FF",
		39221 => x"FF",
		39222 => x"FF",
		39223 => x"FF",
		39224 => x"FF",
		39225 => x"FF",
		39226 => x"FF",
		39227 => x"FF",
		39228 => x"FF",
		39229 => x"FF",
		39230 => x"FF",
		39231 => x"FF",
		39232 => x"FF",
		39233 => x"FF",
		39234 => x"FF",
		39235 => x"FF",
		39236 => x"FF",
		39237 => x"FF",
		39238 => x"FF",
		39239 => x"FF",
		39240 => x"FF",
		39241 => x"FF",
		39242 => x"FF",
		39243 => x"FF",
		39244 => x"FF",
		39245 => x"FF",
		39246 => x"FF",
		39247 => x"FF",
		39248 => x"FF",
		39249 => x"FF",
		39250 => x"FF",
		39251 => x"FF",
		39252 => x"FF",
		39253 => x"FF",
		39254 => x"FF",
		39255 => x"FF",
		39256 => x"FF",
		39257 => x"FF",
		39258 => x"FF",
		39259 => x"FF",
		39260 => x"FF",
		39261 => x"FF",
		39262 => x"FF",
		39263 => x"FF",
		39264 => x"FF",
		39265 => x"FF",
		39266 => x"FF",
		39267 => x"FF",
		39268 => x"FF",
		39269 => x"FF",
		39270 => x"FF",
		39271 => x"FF",
		39272 => x"FF",
		39273 => x"FF",
		39274 => x"FF",
		39275 => x"FF",
		39276 => x"FF",
		39277 => x"FF",
		39278 => x"FF",
		39279 => x"FF",
		39280 => x"FF",
		39281 => x"FF",
		39282 => x"FF",
		39283 => x"FF",
		39284 => x"FF",
		39285 => x"FF",
		39286 => x"FF",
		39287 => x"FF",
		39288 => x"FF",
		39289 => x"FF",
		39290 => x"FF",
		39291 => x"FF",
		39292 => x"FF",
		39293 => x"FF",
		39294 => x"FF",
		39295 => x"FF",
		39296 => x"FF",
		39297 => x"FF",
		39298 => x"FF",
		39299 => x"FF",
		39300 => x"FF",
		39301 => x"FF",
		39302 => x"FF",
		39303 => x"FF",
		39304 => x"FF",
		39305 => x"FF",
		39306 => x"FF",
		39307 => x"FF",
		39308 => x"FF",
		39309 => x"FF",
		39310 => x"FF",
		39311 => x"FF",
		39312 => x"FF",
		39313 => x"FF",
		39314 => x"FF",
		39315 => x"FF",
		39316 => x"FF",
		39317 => x"FF",
		39318 => x"FF",
		39319 => x"FF",
		39320 => x"FF",
		39321 => x"FF",
		39322 => x"FF",
		39323 => x"FF",
		39324 => x"FF",
		39325 => x"FF",
		39326 => x"FF",
		39327 => x"FF",
		39328 => x"FF",
		39329 => x"FF",
		39330 => x"FF",
		39331 => x"FF",
		39332 => x"FF",
		39333 => x"FF",
		39334 => x"FF",
		39335 => x"FF",
		39336 => x"FF",
		39337 => x"FF",
		39338 => x"FF",
		39339 => x"FF",
		39340 => x"FF",
		39341 => x"FF",
		39342 => x"FF",
		39343 => x"FF",
		39344 => x"FF",
		39345 => x"FF",
		39346 => x"FF",
		39347 => x"FF",
		39348 => x"FF",
		39349 => x"FF",
		39350 => x"FF",
		39351 => x"FF",
		39352 => x"FF",
		39353 => x"FF",
		39354 => x"FF",
		39355 => x"FF",
		39356 => x"FF",
		39357 => x"FF",
		39358 => x"FF",
		39359 => x"FF",
		39360 => x"FF",
		39361 => x"FF",
		39362 => x"FF",
		39363 => x"FF",
		39364 => x"FF",
		39365 => x"FF",
		39366 => x"FF",
		39367 => x"FF",
		39368 => x"FF",
		39369 => x"FF",
		39370 => x"FF",
		39371 => x"FF",
		39372 => x"FF",
		39373 => x"FF",
		39374 => x"FF",
		39375 => x"FF",
		39376 => x"FF",
		39377 => x"FF",
		39378 => x"FF",
		39379 => x"FF",
		39380 => x"FF",
		39381 => x"FF",
		39382 => x"FF",
		39383 => x"FF",
		39384 => x"FF",
		39385 => x"FF",
		39386 => x"FF",
		39451 => x"FF",
		39452 => x"FF",
		39453 => x"FF",
		39454 => x"FF",
		39455 => x"FF",
		39456 => x"FF",
		39457 => x"FF",
		39458 => x"FF",
		39459 => x"FF",
		39460 => x"FF",
		39461 => x"FF",
		39462 => x"FF",
		39463 => x"FF",
		39464 => x"FF",
		39465 => x"FF",
		39466 => x"FF",
		39467 => x"FF",
		39468 => x"FF",
		39469 => x"FF",
		39470 => x"FF",
		39471 => x"FF",
		39472 => x"FF",
		39473 => x"FF",
		39474 => x"FF",
		39475 => x"FF",
		39476 => x"FF",
		39477 => x"FF",
		39478 => x"FF",
		39479 => x"FF",
		39480 => x"FF",
		39481 => x"FF",
		39482 => x"FF",
		39483 => x"FF",
		39484 => x"FF",
		39485 => x"FF",
		39486 => x"FF",
		39487 => x"FF",
		39488 => x"FF",
		39489 => x"FF",
		39490 => x"FF",
		39491 => x"FF",
		39492 => x"FF",
		39493 => x"FF",
		39494 => x"FF",
		39495 => x"FF",
		39496 => x"FF",
		39497 => x"FF",
		39498 => x"FF",
		39499 => x"FF",
		39500 => x"FF",
		39501 => x"FF",
		39502 => x"FF",
		39503 => x"FF",
		39504 => x"FF",
		39505 => x"FF",
		39506 => x"FF",
		39507 => x"FF",
		39508 => x"FF",
		39509 => x"FF",
		39510 => x"FF",
		39511 => x"FF",
		39512 => x"FF",
		39513 => x"FF",
		39514 => x"FF",
		39515 => x"FF",
		39516 => x"FF",
		39517 => x"FF",
		39518 => x"FF",
		39519 => x"FF",
		39520 => x"FF",
		39521 => x"FF",
		39522 => x"FF",
		39523 => x"FF",
		39524 => x"FF",
		39525 => x"FF",
		39526 => x"FF",
		39527 => x"FF",
		39528 => x"FF",
		39529 => x"FF",
		39530 => x"FF",
		39531 => x"FF",
		39532 => x"FF",
		39533 => x"FF",
		39534 => x"FF",
		39535 => x"FF",
		39536 => x"FF",
		39537 => x"FF",
		39538 => x"FF",
		39539 => x"FF",
		39540 => x"FF",
		39541 => x"FF",
		39542 => x"FF",
		39543 => x"FF",
		39544 => x"FF",
		39545 => x"FF",
		39546 => x"FF",
		39547 => x"FF",
		39548 => x"FF",
		39549 => x"FF",
		39550 => x"FF",
		39551 => x"FF",
		39552 => x"FF",
		39553 => x"FF",
		39554 => x"FF",
		39555 => x"FF",
		39556 => x"FF",
		39557 => x"FF",
		39558 => x"FF",
		39559 => x"FF",
		39560 => x"FF",
		39561 => x"FF",
		39562 => x"FF",
		39563 => x"FF",
		39564 => x"FF",
		39565 => x"FF",
		39566 => x"FF",
		39567 => x"FF",
		39568 => x"FF",
		39569 => x"FF",
		39570 => x"FF",
		39571 => x"FF",
		39572 => x"FF",
		39573 => x"FF",
		39574 => x"FF",
		39575 => x"FF",
		39576 => x"FF",
		39577 => x"FF",
		39578 => x"FF",
		39579 => x"FF",
		39580 => x"FF",
		39581 => x"FF",
		39582 => x"FF",
		39583 => x"FF",
		39584 => x"FF",
		39585 => x"FF",
		39586 => x"FF",
		39587 => x"FF",
		39588 => x"FF",
		39589 => x"FF",
		39590 => x"FF",
		39591 => x"FF",
		39592 => x"FF",
		39593 => x"FF",
		39594 => x"FF",
		39595 => x"FF",
		39596 => x"FF",
		39597 => x"FF",
		39598 => x"FF",
		39599 => x"FF",
		39600 => x"FF",
		39601 => x"FF",
		39602 => x"FF",
		39603 => x"FF",
		39604 => x"FF",
		39605 => x"FF",
		39606 => x"FF",
		39607 => x"FF",
		39608 => x"FF",
		39609 => x"FF",
		39610 => x"FF",
		39611 => x"FF",
		39612 => x"FF",
		39613 => x"FF",
		39614 => x"FF",
		39615 => x"FF",
		39616 => x"FF",
		39617 => x"FF",
		39618 => x"FF",
		39619 => x"FF",
		39620 => x"FF",
		39621 => x"FF",
		39622 => x"FF",
		39623 => x"FF",
		39624 => x"FF",
		39625 => x"FF",
		39626 => x"FF",
		39627 => x"FF",
		39628 => x"FF",
		39629 => x"FF",
		39630 => x"FF",
		39631 => x"FF",
		39632 => x"FF",
		39633 => x"FF",
		39634 => x"FF",
		39635 => x"FF",
		39636 => x"FF",
		39637 => x"FF",
		39638 => x"FF",
		39639 => x"FF",
		39640 => x"FF",
		39641 => x"FF",
		39642 => x"FF",
		39707 => x"FF",
		39708 => x"FF",
		39709 => x"FF",
		39710 => x"FF",
		39711 => x"FF",
		39712 => x"FF",
		39713 => x"FF",
		39714 => x"FF",
		39715 => x"FF",
		39716 => x"FF",
		39717 => x"FF",
		39718 => x"FF",
		39719 => x"FF",
		39720 => x"FF",
		39721 => x"FF",
		39722 => x"FF",
		39723 => x"FF",
		39724 => x"FF",
		39725 => x"FF",
		39726 => x"FF",
		39727 => x"FF",
		39728 => x"FF",
		39729 => x"FF",
		39730 => x"FF",
		39731 => x"FF",
		39732 => x"FF",
		39733 => x"FF",
		39734 => x"FF",
		39735 => x"FF",
		39736 => x"FF",
		39737 => x"FF",
		39738 => x"FF",
		39739 => x"FF",
		39740 => x"FF",
		39741 => x"FF",
		39742 => x"FF",
		39743 => x"FF",
		39744 => x"FF",
		39745 => x"FF",
		39746 => x"FF",
		39747 => x"FF",
		39748 => x"FF",
		39749 => x"FF",
		39750 => x"FF",
		39751 => x"FF",
		39752 => x"FF",
		39753 => x"FF",
		39754 => x"FF",
		39755 => x"FF",
		39756 => x"FF",
		39757 => x"FF",
		39758 => x"FF",
		39759 => x"FF",
		39760 => x"FF",
		39761 => x"FF",
		39762 => x"FF",
		39763 => x"FF",
		39764 => x"FF",
		39765 => x"FF",
		39766 => x"FF",
		39767 => x"FF",
		39768 => x"FF",
		39769 => x"FF",
		39770 => x"FF",
		39771 => x"FF",
		39772 => x"FF",
		39773 => x"FF",
		39774 => x"FF",
		39775 => x"FF",
		39776 => x"FF",
		39777 => x"FF",
		39778 => x"FF",
		39779 => x"FF",
		39780 => x"FF",
		39781 => x"FF",
		39782 => x"FF",
		39783 => x"FF",
		39784 => x"FF",
		39785 => x"FF",
		39786 => x"FF",
		39787 => x"FF",
		39788 => x"FF",
		39789 => x"FF",
		39790 => x"FF",
		39791 => x"FF",
		39792 => x"FF",
		39793 => x"FF",
		39794 => x"FF",
		39795 => x"FF",
		39796 => x"FF",
		39797 => x"FF",
		39798 => x"FF",
		39799 => x"FF",
		39800 => x"FF",
		39801 => x"FF",
		39802 => x"FF",
		39803 => x"FF",
		39804 => x"FF",
		39805 => x"FF",
		39806 => x"FF",
		39807 => x"FF",
		39808 => x"FF",
		39809 => x"FF",
		39810 => x"FF",
		39811 => x"FF",
		39812 => x"FF",
		39813 => x"FF",
		39814 => x"FF",
		39815 => x"FF",
		39816 => x"FF",
		39817 => x"FF",
		39818 => x"FF",
		39819 => x"FF",
		39820 => x"FF",
		39821 => x"FF",
		39822 => x"FF",
		39823 => x"FF",
		39824 => x"FF",
		39825 => x"FF",
		39826 => x"FF",
		39827 => x"FF",
		39828 => x"FF",
		39829 => x"FF",
		39830 => x"FF",
		39831 => x"FF",
		39832 => x"FF",
		39833 => x"FF",
		39834 => x"FF",
		39835 => x"FF",
		39836 => x"FF",
		39837 => x"FF",
		39838 => x"FF",
		39839 => x"FF",
		39840 => x"FF",
		39841 => x"FF",
		39842 => x"FF",
		39843 => x"FF",
		39844 => x"FF",
		39845 => x"FF",
		39846 => x"FF",
		39847 => x"FF",
		39848 => x"FF",
		39849 => x"FF",
		39850 => x"FF",
		39851 => x"FF",
		39852 => x"FF",
		39853 => x"FF",
		39854 => x"FF",
		39855 => x"FF",
		39856 => x"FF",
		39857 => x"FF",
		39858 => x"FF",
		39859 => x"FF",
		39860 => x"FF",
		39861 => x"FF",
		39862 => x"FF",
		39863 => x"FF",
		39864 => x"FF",
		39865 => x"FF",
		39866 => x"FF",
		39867 => x"FF",
		39868 => x"FF",
		39869 => x"FF",
		39870 => x"FF",
		39871 => x"FF",
		39872 => x"FF",
		39873 => x"FF",
		39874 => x"FF",
		39875 => x"FF",
		39876 => x"FF",
		39877 => x"FF",
		39878 => x"FF",
		39879 => x"FF",
		39880 => x"FF",
		39881 => x"FF",
		39882 => x"FF",
		39883 => x"FF",
		39884 => x"FF",
		39885 => x"FF",
		39886 => x"FF",
		39887 => x"FF",
		39888 => x"FF",
		39889 => x"FF",
		39890 => x"FF",
		39891 => x"FF",
		39892 => x"FF",
		39893 => x"FF",
		39894 => x"FF",
		39895 => x"FF",
		39896 => x"FF",
		39897 => x"FF",
		39898 => x"FF",
		39963 => x"FF",
		39964 => x"FF",
		39965 => x"FF",
		40026 => x"FF",
		40027 => x"FF",
		40028 => x"FF",
		40089 => x"FF",
		40090 => x"FF",
		40091 => x"FF",
		40152 => x"FF",
		40153 => x"FF",
		40154 => x"FF",
		40219 => x"FF",
		40220 => x"FF",
		40221 => x"FF",
		40282 => x"FF",
		40283 => x"FF",
		40284 => x"FF",
		40345 => x"FF",
		40346 => x"FF",
		40347 => x"FF",
		40408 => x"FF",
		40409 => x"FF",
		40410 => x"FF",
		40475 => x"FF",
		40476 => x"FF",
		40477 => x"FF",
		40538 => x"FF",
		40539 => x"FF",
		40540 => x"FF",
		40601 => x"FF",
		40602 => x"FF",
		40603 => x"FF",
		40664 => x"FF",
		40665 => x"FF",
		40666 => x"FF",
		40731 => x"FF",
		40732 => x"FF",
		40733 => x"FF",
		40794 => x"FF",
		40795 => x"FF",
		40796 => x"FF",
		40857 => x"FF",
		40858 => x"FF",
		40859 => x"FF",
		40920 => x"FF",
		40921 => x"FF",
		40922 => x"FF",
		40987 => x"FF",
		40988 => x"FF",
		40989 => x"FF",
		41050 => x"FF",
		41051 => x"FF",
		41052 => x"FF",
		41113 => x"FF",
		41114 => x"FF",
		41115 => x"FF",
		41176 => x"FF",
		41177 => x"FF",
		41178 => x"FF",
		41243 => x"FF",
		41244 => x"FF",
		41245 => x"FF",
		41306 => x"FF",
		41307 => x"FF",
		41308 => x"FF",
		41369 => x"FF",
		41370 => x"FF",
		41371 => x"FF",
		41432 => x"FF",
		41433 => x"FF",
		41434 => x"FF",
		41499 => x"FF",
		41500 => x"FF",
		41501 => x"FF",
		41562 => x"FF",
		41563 => x"FF",
		41564 => x"FF",
		41625 => x"FF",
		41626 => x"FF",
		41627 => x"FF",
		41688 => x"FF",
		41689 => x"FF",
		41690 => x"FF",
		41755 => x"FF",
		41756 => x"FF",
		41757 => x"FF",
		41818 => x"FF",
		41819 => x"FF",
		41820 => x"FF",
		41881 => x"FF",
		41882 => x"FF",
		41883 => x"FF",
		41944 => x"FF",
		41945 => x"FF",
		41946 => x"FF",
		42011 => x"FF",
		42012 => x"FF",
		42013 => x"FF",
		42074 => x"FF",
		42075 => x"FF",
		42076 => x"FF",
		42137 => x"FF",
		42138 => x"FF",
		42139 => x"FF",
		42200 => x"FF",
		42201 => x"FF",
		42202 => x"FF",
		42267 => x"FF",
		42268 => x"FF",
		42269 => x"FF",
		42330 => x"FF",
		42331 => x"FF",
		42332 => x"FF",
		42393 => x"FF",
		42394 => x"FF",
		42395 => x"FF",
		42456 => x"FF",
		42457 => x"FF",
		42458 => x"FF",
		42523 => x"FF",
		42524 => x"FF",
		42525 => x"FF",
		42586 => x"FF",
		42587 => x"FF",
		42588 => x"FF",
		42649 => x"FF",
		42650 => x"FF",
		42651 => x"FF",
		42712 => x"FF",
		42713 => x"FF",
		42714 => x"FF",
		42779 => x"FF",
		42780 => x"FF",
		42781 => x"FF",
		42842 => x"FF",
		42843 => x"FF",
		42844 => x"FF",
		42905 => x"FF",
		42906 => x"FF",
		42907 => x"FF",
		42968 => x"FF",
		42969 => x"FF",
		42970 => x"FF",
		43035 => x"FF",
		43036 => x"FF",
		43037 => x"FF",
		43098 => x"FF",
		43099 => x"FF",
		43100 => x"FF",
		43161 => x"FF",
		43162 => x"FF",
		43163 => x"FF",
		43224 => x"FF",
		43225 => x"FF",
		43226 => x"FF",
		43291 => x"FF",
		43292 => x"FF",
		43293 => x"FF",
		43354 => x"FF",
		43355 => x"FF",
		43356 => x"FF",
		43417 => x"FF",
		43418 => x"FF",
		43419 => x"FF",
		43480 => x"FF",
		43481 => x"FF",
		43482 => x"FF",
		43547 => x"FF",
		43548 => x"FF",
		43549 => x"FF",
		43610 => x"FF",
		43611 => x"FF",
		43612 => x"FF",
		43673 => x"FF",
		43674 => x"FF",
		43675 => x"FF",
		43736 => x"FF",
		43737 => x"FF",
		43738 => x"FF",
		43803 => x"FF",
		43804 => x"FF",
		43805 => x"FF",
		43866 => x"FF",
		43867 => x"FF",
		43868 => x"FF",
		43929 => x"FF",
		43930 => x"FF",
		43931 => x"FF",
		43992 => x"FF",
		43993 => x"FF",
		43994 => x"FF",
		44059 => x"FF",
		44060 => x"FF",
		44061 => x"FF",
		44122 => x"FF",
		44123 => x"FF",
		44124 => x"FF",
		44185 => x"FF",
		44186 => x"FF",
		44187 => x"FF",
		44248 => x"FF",
		44249 => x"FF",
		44250 => x"FF",
		44315 => x"FF",
		44316 => x"FF",
		44317 => x"FF",
		44378 => x"FF",
		44379 => x"FF",
		44380 => x"FF",
		44441 => x"FF",
		44442 => x"FF",
		44443 => x"FF",
		44504 => x"FF",
		44505 => x"FF",
		44506 => x"FF",
		44571 => x"FF",
		44572 => x"FF",
		44573 => x"FF",
		44634 => x"FF",
		44635 => x"FF",
		44636 => x"FF",
		44697 => x"FF",
		44698 => x"FF",
		44699 => x"FF",
		44760 => x"FF",
		44761 => x"FF",
		44762 => x"FF",
		44827 => x"FF",
		44828 => x"FF",
		44829 => x"FF",
		44890 => x"FF",
		44891 => x"FF",
		44892 => x"FF",
		44953 => x"FF",
		44954 => x"FF",
		44955 => x"FF",
		45016 => x"FF",
		45017 => x"FF",
		45018 => x"FF",
		45083 => x"FF",
		45084 => x"FF",
		45085 => x"FF",
		45146 => x"FF",
		45147 => x"FF",
		45148 => x"FF",
		45209 => x"FF",
		45210 => x"FF",
		45211 => x"FF",
		45272 => x"FF",
		45273 => x"FF",
		45274 => x"FF",
		45339 => x"FF",
		45340 => x"FF",
		45341 => x"FF",
		45402 => x"FF",
		45403 => x"FF",
		45404 => x"FF",
		45465 => x"FF",
		45466 => x"FF",
		45467 => x"FF",
		45528 => x"FF",
		45529 => x"FF",
		45530 => x"FF",
		45595 => x"FF",
		45596 => x"FF",
		45597 => x"FF",
		45658 => x"FF",
		45659 => x"FF",
		45660 => x"FF",
		45721 => x"FF",
		45722 => x"FF",
		45723 => x"FF",
		45784 => x"FF",
		45785 => x"FF",
		45786 => x"FF",
		45851 => x"FF",
		45852 => x"FF",
		45853 => x"FF",
		45914 => x"FF",
		45915 => x"FF",
		45916 => x"FF",
		45977 => x"FF",
		45978 => x"FF",
		45979 => x"FF",
		46040 => x"FF",
		46041 => x"FF",
		46042 => x"FF",
		46107 => x"FF",
		46108 => x"FF",
		46109 => x"FF",
		46170 => x"FF",
		46171 => x"FF",
		46172 => x"FF",
		46233 => x"FF",
		46234 => x"FF",
		46235 => x"FF",
		46296 => x"FF",
		46297 => x"FF",
		46298 => x"FF",
		46363 => x"FF",
		46364 => x"FF",
		46365 => x"FF",
		46426 => x"FF",
		46427 => x"FF",
		46428 => x"FF",
		46489 => x"FF",
		46490 => x"FF",
		46491 => x"FF",
		46552 => x"FF",
		46553 => x"FF",
		46554 => x"FF",
		46619 => x"FF",
		46620 => x"FF",
		46621 => x"FF",
		46682 => x"FF",
		46683 => x"FF",
		46684 => x"FF",
		46745 => x"FF",
		46746 => x"FF",
		46747 => x"FF",
		46808 => x"FF",
		46809 => x"FF",
		46810 => x"FF",
		46875 => x"FF",
		46876 => x"FF",
		46877 => x"FF",
		46938 => x"FF",
		46939 => x"FF",
		46940 => x"FF",
		47001 => x"FF",
		47002 => x"FF",
		47003 => x"FF",
		47064 => x"FF",
		47065 => x"FF",
		47066 => x"FF",
		47131 => x"FF",
		47132 => x"FF",
		47133 => x"FF",
		47194 => x"FF",
		47195 => x"FF",
		47196 => x"FF",
		47257 => x"FF",
		47258 => x"FF",
		47259 => x"FF",
		47320 => x"FF",
		47321 => x"FF",
		47322 => x"FF",
		47387 => x"FF",
		47388 => x"FF",
		47389 => x"FF",
		47450 => x"FF",
		47451 => x"FF",
		47452 => x"FF",
		47513 => x"FF",
		47514 => x"FF",
		47515 => x"FF",
		47576 => x"FF",
		47577 => x"FF",
		47578 => x"FF",
		47643 => x"FF",
		47644 => x"FF",
		47645 => x"FF",
		47706 => x"FF",
		47707 => x"FF",
		47708 => x"FF",
		47769 => x"FF",
		47770 => x"FF",
		47771 => x"FF",
		47832 => x"FF",
		47833 => x"FF",
		47834 => x"FF",
		47899 => x"FF",
		47900 => x"FF",
		47901 => x"FF",
		47962 => x"FF",
		47963 => x"FF",
		47964 => x"FF",
		48025 => x"FF",
		48026 => x"FF",
		48027 => x"FF",
		48088 => x"FF",
		48089 => x"FF",
		48090 => x"FF",
		48155 => x"FF",
		48156 => x"FF",
		48157 => x"FF",
		48218 => x"FF",
		48219 => x"FF",
		48220 => x"FF",
		48281 => x"FF",
		48282 => x"FF",
		48283 => x"FF",
		48344 => x"FF",
		48345 => x"FF",
		48346 => x"FF",
		48411 => x"FF",
		48412 => x"FF",
		48413 => x"FF",
		48474 => x"FF",
		48475 => x"FF",
		48476 => x"FF",
		48537 => x"FF",
		48538 => x"FF",
		48539 => x"FF",
		48600 => x"FF",
		48601 => x"FF",
		48602 => x"FF",
		48667 => x"FF",
		48668 => x"FF",
		48669 => x"FF",
		48730 => x"FF",
		48731 => x"FF",
		48732 => x"FF",
		48793 => x"FF",
		48794 => x"FF",
		48795 => x"FF",
		48856 => x"FF",
		48857 => x"FF",
		48858 => x"FF",
		48923 => x"FF",
		48924 => x"FF",
		48925 => x"FF",
		48986 => x"FF",
		48987 => x"FF",
		48988 => x"FF",
		49049 => x"FF",
		49050 => x"FF",
		49051 => x"FF",
		49112 => x"FF",
		49113 => x"FF",
		49114 => x"FF",
		49179 => x"FF",
		49180 => x"FF",
		49181 => x"FF",
		49242 => x"FF",
		49243 => x"FF",
		49244 => x"FF",
		49305 => x"FF",
		49306 => x"FF",
		49307 => x"FF",
		49368 => x"FF",
		49369 => x"FF",
		49370 => x"FF",
		49435 => x"FF",
		49436 => x"FF",
		49437 => x"FF",
		49498 => x"FF",
		49499 => x"FF",
		49500 => x"FF",
		49561 => x"FF",
		49562 => x"FF",
		49563 => x"FF",
		49624 => x"FF",
		49625 => x"FF",
		49626 => x"FF",
		49691 => x"FF",
		49692 => x"FF",
		49693 => x"FF",
		49754 => x"FF",
		49755 => x"FF",
		49756 => x"FF",
		49817 => x"FF",
		49818 => x"FF",
		49819 => x"FF",
		49880 => x"FF",
		49881 => x"FF",
		49882 => x"FF",
		49947 => x"FF",
		49948 => x"FF",
		49949 => x"FF",
		50010 => x"FF",
		50011 => x"FF",
		50012 => x"FF",
		50073 => x"FF",
		50074 => x"FF",
		50075 => x"FF",
		50136 => x"FF",
		50137 => x"FF",
		50138 => x"FF",
		50203 => x"FF",
		50204 => x"FF",
		50205 => x"FF",
		50266 => x"FF",
		50267 => x"FF",
		50268 => x"FF",
		50329 => x"FF",
		50330 => x"FF",
		50331 => x"FF",
		50392 => x"FF",
		50393 => x"FF",
		50394 => x"FF",
		50459 => x"FF",
		50460 => x"FF",
		50461 => x"FF",
		50522 => x"FF",
		50523 => x"FF",
		50524 => x"FF",
		50585 => x"FF",
		50586 => x"FF",
		50587 => x"FF",
		50648 => x"FF",
		50649 => x"FF",
		50650 => x"FF",
		50715 => x"FF",
		50716 => x"FF",
		50717 => x"FF",
		50778 => x"FF",
		50779 => x"FF",
		50780 => x"FF",
		50841 => x"FF",
		50842 => x"FF",
		50843 => x"FF",
		50904 => x"FF",
		50905 => x"FF",
		50906 => x"FF",
		50971 => x"FF",
		50972 => x"FF",
		50973 => x"FF",
		51034 => x"FF",
		51035 => x"FF",
		51036 => x"FF",
		51097 => x"FF",
		51098 => x"FF",
		51099 => x"FF",
		51160 => x"FF",
		51161 => x"FF",
		51162 => x"FF",
		51227 => x"FF",
		51228 => x"FF",
		51229 => x"FF",
		51290 => x"FF",
		51291 => x"FF",
		51292 => x"FF",
		51353 => x"FF",
		51354 => x"FF",
		51355 => x"FF",
		51416 => x"FF",
		51417 => x"FF",
		51418 => x"FF",
		51483 => x"FF",
		51484 => x"FF",
		51485 => x"FF",
		51546 => x"FF",
		51547 => x"FF",
		51548 => x"FF",
		51609 => x"FF",
		51610 => x"FF",
		51611 => x"FF",
		51672 => x"FF",
		51673 => x"FF",
		51674 => x"FF",
		51739 => x"FF",
		51740 => x"FF",
		51741 => x"FF",
		51802 => x"FF",
		51803 => x"FF",
		51804 => x"FF",
		51865 => x"FF",
		51866 => x"FF",
		51867 => x"FF",
		51928 => x"FF",
		51929 => x"FF",
		51930 => x"FF",
		51995 => x"FF",
		51996 => x"FF",
		51997 => x"FF",
		52058 => x"FF",
		52059 => x"FF",
		52060 => x"FF",
		52121 => x"FF",
		52122 => x"FF",
		52123 => x"FF",
		52184 => x"FF",
		52185 => x"FF",
		52186 => x"FF",
		52251 => x"FF",
		52252 => x"FF",
		52253 => x"FF",
		52314 => x"FF",
		52315 => x"FF",
		52316 => x"FF",
		52377 => x"FF",
		52378 => x"FF",
		52379 => x"FF",
		52440 => x"FF",
		52441 => x"FF",
		52442 => x"FF",
		52507 => x"FF",
		52508 => x"FF",
		52509 => x"FF",
		52570 => x"FF",
		52571 => x"FF",
		52572 => x"FF",
		52633 => x"FF",
		52634 => x"FF",
		52635 => x"FF",
		52696 => x"FF",
		52697 => x"FF",
		52698 => x"FF",
		52763 => x"FF",
		52764 => x"FF",
		52765 => x"FF",
		52826 => x"FF",
		52827 => x"FF",
		52828 => x"FF",
		52889 => x"FF",
		52890 => x"FF",
		52891 => x"FF",
		52952 => x"FF",
		52953 => x"FF",
		52954 => x"FF",
		53019 => x"FF",
		53020 => x"FF",
		53021 => x"FF",
		53082 => x"FF",
		53083 => x"FF",
		53084 => x"FF",
		53145 => x"FF",
		53146 => x"FF",
		53147 => x"FF",
		53208 => x"FF",
		53209 => x"FF",
		53210 => x"FF",
		53275 => x"FF",
		53276 => x"FF",
		53277 => x"FF",
		53338 => x"FF",
		53339 => x"FF",
		53340 => x"FF",
		53401 => x"FF",
		53402 => x"FF",
		53403 => x"FF",
		53464 => x"FF",
		53465 => x"FF",
		53466 => x"FF",
		53531 => x"FF",
		53532 => x"FF",
		53533 => x"FF",
		53594 => x"FF",
		53595 => x"FF",
		53596 => x"FF",
		53657 => x"FF",
		53658 => x"FF",
		53659 => x"FF",
		53720 => x"FF",
		53721 => x"FF",
		53722 => x"FF",
		53787 => x"FF",
		53788 => x"FF",
		53789 => x"FF",
		53850 => x"FF",
		53851 => x"FF",
		53852 => x"FF",
		53913 => x"FF",
		53914 => x"FF",
		53915 => x"FF",
		53976 => x"FF",
		53977 => x"FF",
		53978 => x"FF",
		54043 => x"FF",
		54044 => x"FF",
		54045 => x"FF",
		54106 => x"FF",
		54107 => x"FF",
		54108 => x"FF",
		54169 => x"FF",
		54170 => x"FF",
		54171 => x"FF",
		54232 => x"FF",
		54233 => x"FF",
		54234 => x"FF",
		54299 => x"FF",
		54300 => x"FF",
		54301 => x"FF",
		54362 => x"FF",
		54363 => x"FF",
		54364 => x"FF",
		54425 => x"FF",
		54426 => x"FF",
		54427 => x"FF",
		54488 => x"FF",
		54489 => x"FF",
		54490 => x"FF",
		54555 => x"FF",
		54556 => x"FF",
		54557 => x"FF",
		54618 => x"FF",
		54619 => x"FF",
		54620 => x"FF",
		54681 => x"FF",
		54682 => x"FF",
		54683 => x"FF",
		54744 => x"FF",
		54745 => x"FF",
		54746 => x"FF",
		54811 => x"FF",
		54812 => x"FF",
		54813 => x"FF",
		54874 => x"FF",
		54875 => x"FF",
		54876 => x"FF",
		54937 => x"FF",
		54938 => x"FF",
		54939 => x"FF",
		55000 => x"FF",
		55001 => x"FF",
		55002 => x"FF",
		55067 => x"FF",
		55068 => x"FF",
		55069 => x"FF",
		55130 => x"FF",
		55131 => x"FF",
		55132 => x"FF",
		55193 => x"FF",
		55194 => x"FF",
		55195 => x"FF",
		55256 => x"FF",
		55257 => x"FF",
		55258 => x"FF",
		55323 => x"FF",
		55324 => x"FF",
		55325 => x"FF",
		55326 => x"FF",
		55327 => x"FF",
		55328 => x"FF",
		55329 => x"FF",
		55330 => x"FF",
		55331 => x"FF",
		55332 => x"FF",
		55333 => x"FF",
		55334 => x"FF",
		55335 => x"FF",
		55336 => x"FF",
		55337 => x"FF",
		55338 => x"FF",
		55339 => x"FF",
		55340 => x"FF",
		55341 => x"FF",
		55342 => x"FF",
		55343 => x"FF",
		55344 => x"FF",
		55345 => x"FF",
		55346 => x"FF",
		55347 => x"FF",
		55348 => x"FF",
		55349 => x"FF",
		55350 => x"FF",
		55351 => x"FF",
		55352 => x"FF",
		55353 => x"FF",
		55354 => x"FF",
		55355 => x"FF",
		55356 => x"FF",
		55357 => x"FF",
		55358 => x"FF",
		55359 => x"FF",
		55360 => x"FF",
		55361 => x"FF",
		55362 => x"FF",
		55363 => x"FF",
		55364 => x"FF",
		55365 => x"FF",
		55366 => x"FF",
		55367 => x"FF",
		55368 => x"FF",
		55369 => x"FF",
		55370 => x"FF",
		55371 => x"FF",
		55372 => x"FF",
		55373 => x"FF",
		55374 => x"FF",
		55375 => x"FF",
		55376 => x"FF",
		55377 => x"FF",
		55378 => x"FF",
		55379 => x"FF",
		55380 => x"FF",
		55381 => x"FF",
		55382 => x"FF",
		55383 => x"FF",
		55384 => x"FF",
		55385 => x"FF",
		55386 => x"FF",
		55387 => x"FF",
		55388 => x"FF",
		55389 => x"FF",
		55390 => x"FF",
		55391 => x"FF",
		55392 => x"FF",
		55393 => x"FF",
		55394 => x"FF",
		55395 => x"FF",
		55396 => x"FF",
		55397 => x"FF",
		55398 => x"FF",
		55399 => x"FF",
		55400 => x"FF",
		55401 => x"FF",
		55402 => x"FF",
		55403 => x"FF",
		55404 => x"FF",
		55405 => x"FF",
		55406 => x"FF",
		55407 => x"FF",
		55408 => x"FF",
		55409 => x"FF",
		55410 => x"FF",
		55411 => x"FF",
		55412 => x"FF",
		55413 => x"FF",
		55414 => x"FF",
		55415 => x"FF",
		55416 => x"FF",
		55417 => x"FF",
		55418 => x"FF",
		55419 => x"FF",
		55420 => x"FF",
		55421 => x"FF",
		55422 => x"FF",
		55423 => x"FF",
		55424 => x"FF",
		55425 => x"FF",
		55426 => x"FF",
		55427 => x"FF",
		55428 => x"FF",
		55429 => x"FF",
		55430 => x"FF",
		55431 => x"FF",
		55432 => x"FF",
		55433 => x"FF",
		55434 => x"FF",
		55435 => x"FF",
		55436 => x"FF",
		55437 => x"FF",
		55438 => x"FF",
		55439 => x"FF",
		55440 => x"FF",
		55441 => x"FF",
		55442 => x"FF",
		55443 => x"FF",
		55444 => x"FF",
		55445 => x"FF",
		55446 => x"FF",
		55447 => x"FF",
		55448 => x"FF",
		55449 => x"FF",
		55450 => x"FF",
		55451 => x"FF",
		55452 => x"FF",
		55453 => x"FF",
		55454 => x"FF",
		55455 => x"FF",
		55456 => x"FF",
		55457 => x"FF",
		55458 => x"FF",
		55459 => x"FF",
		55460 => x"FF",
		55461 => x"FF",
		55462 => x"FF",
		55463 => x"FF",
		55464 => x"FF",
		55465 => x"FF",
		55466 => x"FF",
		55467 => x"FF",
		55468 => x"FF",
		55469 => x"FF",
		55470 => x"FF",
		55471 => x"FF",
		55472 => x"FF",
		55473 => x"FF",
		55474 => x"FF",
		55475 => x"FF",
		55476 => x"FF",
		55477 => x"FF",
		55478 => x"FF",
		55479 => x"FF",
		55480 => x"FF",
		55481 => x"FF",
		55482 => x"FF",
		55483 => x"FF",
		55484 => x"FF",
		55485 => x"FF",
		55486 => x"FF",
		55487 => x"FF",
		55488 => x"FF",
		55489 => x"FF",
		55490 => x"FF",
		55491 => x"FF",
		55492 => x"FF",
		55493 => x"FF",
		55494 => x"FF",
		55495 => x"FF",
		55496 => x"FF",
		55497 => x"FF",
		55498 => x"FF",
		55499 => x"FF",
		55500 => x"FF",
		55501 => x"FF",
		55502 => x"FF",
		55503 => x"FF",
		55504 => x"FF",
		55505 => x"FF",
		55506 => x"FF",
		55507 => x"FF",
		55508 => x"FF",
		55509 => x"FF",
		55510 => x"FF",
		55511 => x"FF",
		55512 => x"FF",
		55513 => x"FF",
		55514 => x"FF",
		55579 => x"FF",
		55580 => x"FF",
		55581 => x"FF",
		55582 => x"FF",
		55583 => x"FF",
		55584 => x"FF",
		55585 => x"FF",
		55586 => x"FF",
		55587 => x"FF",
		55588 => x"FF",
		55589 => x"FF",
		55590 => x"FF",
		55591 => x"FF",
		55592 => x"FF",
		55593 => x"FF",
		55594 => x"FF",
		55595 => x"FF",
		55596 => x"FF",
		55597 => x"FF",
		55598 => x"FF",
		55599 => x"FF",
		55600 => x"FF",
		55601 => x"FF",
		55602 => x"FF",
		55603 => x"FF",
		55604 => x"FF",
		55605 => x"FF",
		55606 => x"FF",
		55607 => x"FF",
		55608 => x"FF",
		55609 => x"FF",
		55610 => x"FF",
		55611 => x"FF",
		55612 => x"FF",
		55613 => x"FF",
		55614 => x"FF",
		55615 => x"FF",
		55616 => x"FF",
		55617 => x"FF",
		55618 => x"FF",
		55619 => x"FF",
		55620 => x"FF",
		55621 => x"FF",
		55622 => x"FF",
		55623 => x"FF",
		55624 => x"FF",
		55625 => x"FF",
		55626 => x"FF",
		55627 => x"FF",
		55628 => x"FF",
		55629 => x"FF",
		55630 => x"FF",
		55631 => x"FF",
		55632 => x"FF",
		55633 => x"FF",
		55634 => x"FF",
		55635 => x"FF",
		55636 => x"FF",
		55637 => x"FF",
		55638 => x"FF",
		55639 => x"FF",
		55640 => x"FF",
		55641 => x"FF",
		55642 => x"FF",
		55643 => x"FF",
		55644 => x"FF",
		55645 => x"FF",
		55646 => x"FF",
		55647 => x"FF",
		55648 => x"FF",
		55649 => x"FF",
		55650 => x"FF",
		55651 => x"FF",
		55652 => x"FF",
		55653 => x"FF",
		55654 => x"FF",
		55655 => x"FF",
		55656 => x"FF",
		55657 => x"FF",
		55658 => x"FF",
		55659 => x"FF",
		55660 => x"FF",
		55661 => x"FF",
		55662 => x"FF",
		55663 => x"FF",
		55664 => x"FF",
		55665 => x"FF",
		55666 => x"FF",
		55667 => x"FF",
		55668 => x"FF",
		55669 => x"FF",
		55670 => x"FF",
		55671 => x"FF",
		55672 => x"FF",
		55673 => x"FF",
		55674 => x"FF",
		55675 => x"FF",
		55676 => x"FF",
		55677 => x"FF",
		55678 => x"FF",
		55679 => x"FF",
		55680 => x"FF",
		55681 => x"FF",
		55682 => x"FF",
		55683 => x"FF",
		55684 => x"FF",
		55685 => x"FF",
		55686 => x"FF",
		55687 => x"FF",
		55688 => x"FF",
		55689 => x"FF",
		55690 => x"FF",
		55691 => x"FF",
		55692 => x"FF",
		55693 => x"FF",
		55694 => x"FF",
		55695 => x"FF",
		55696 => x"FF",
		55697 => x"FF",
		55698 => x"FF",
		55699 => x"FF",
		55700 => x"FF",
		55701 => x"FF",
		55702 => x"FF",
		55703 => x"FF",
		55704 => x"FF",
		55705 => x"FF",
		55706 => x"FF",
		55707 => x"FF",
		55708 => x"FF",
		55709 => x"FF",
		55710 => x"FF",
		55711 => x"FF",
		55712 => x"FF",
		55713 => x"FF",
		55714 => x"FF",
		55715 => x"FF",
		55716 => x"FF",
		55717 => x"FF",
		55718 => x"FF",
		55719 => x"FF",
		55720 => x"FF",
		55721 => x"FF",
		55722 => x"FF",
		55723 => x"FF",
		55724 => x"FF",
		55725 => x"FF",
		55726 => x"FF",
		55727 => x"FF",
		55728 => x"FF",
		55729 => x"FF",
		55730 => x"FF",
		55731 => x"FF",
		55732 => x"FF",
		55733 => x"FF",
		55734 => x"FF",
		55735 => x"FF",
		55736 => x"FF",
		55737 => x"FF",
		55738 => x"FF",
		55739 => x"FF",
		55740 => x"FF",
		55741 => x"FF",
		55742 => x"FF",
		55743 => x"FF",
		55744 => x"FF",
		55745 => x"FF",
		55746 => x"FF",
		55747 => x"FF",
		55748 => x"FF",
		55749 => x"FF",
		55750 => x"FF",
		55751 => x"FF",
		55752 => x"FF",
		55753 => x"FF",
		55754 => x"FF",
		55755 => x"FF",
		55756 => x"FF",
		55757 => x"FF",
		55758 => x"FF",
		55759 => x"FF",
		55760 => x"FF",
		55761 => x"FF",
		55762 => x"FF",
		55763 => x"FF",
		55764 => x"FF",
		55765 => x"FF",
		55766 => x"FF",
		55767 => x"FF",
		55768 => x"FF",
		55769 => x"FF",
		55770 => x"FF",
		55835 => x"FF",
		55836 => x"FF",
		55837 => x"FF",
		55838 => x"FF",
		55839 => x"FF",
		55840 => x"FF",
		55841 => x"FF",
		55842 => x"FF",
		55843 => x"FF",
		55844 => x"FF",
		55845 => x"FF",
		55846 => x"FF",
		55847 => x"FF",
		55848 => x"FF",
		55849 => x"FF",
		55850 => x"FF",
		55851 => x"FF",
		55852 => x"FF",
		55853 => x"FF",
		55854 => x"FF",
		55855 => x"FF",
		55856 => x"FF",
		55857 => x"FF",
		55858 => x"FF",
		55859 => x"FF",
		55860 => x"FF",
		55861 => x"FF",
		55862 => x"FF",
		55863 => x"FF",
		55864 => x"FF",
		55865 => x"FF",
		55866 => x"FF",
		55867 => x"FF",
		55868 => x"FF",
		55869 => x"FF",
		55870 => x"FF",
		55871 => x"FF",
		55872 => x"FF",
		55873 => x"FF",
		55874 => x"FF",
		55875 => x"FF",
		55876 => x"FF",
		55877 => x"FF",
		55878 => x"FF",
		55879 => x"FF",
		55880 => x"FF",
		55881 => x"FF",
		55882 => x"FF",
		55883 => x"FF",
		55884 => x"FF",
		55885 => x"FF",
		55886 => x"FF",
		55887 => x"FF",
		55888 => x"FF",
		55889 => x"FF",
		55890 => x"FF",
		55891 => x"FF",
		55892 => x"FF",
		55893 => x"FF",
		55894 => x"FF",
		55895 => x"FF",
		55896 => x"FF",
		55897 => x"FF",
		55898 => x"FF",
		55899 => x"FF",
		55900 => x"FF",
		55901 => x"FF",
		55902 => x"FF",
		55903 => x"FF",
		55904 => x"FF",
		55905 => x"FF",
		55906 => x"FF",
		55907 => x"FF",
		55908 => x"FF",
		55909 => x"FF",
		55910 => x"FF",
		55911 => x"FF",
		55912 => x"FF",
		55913 => x"FF",
		55914 => x"FF",
		55915 => x"FF",
		55916 => x"FF",
		55917 => x"FF",
		55918 => x"FF",
		55919 => x"FF",
		55920 => x"FF",
		55921 => x"FF",
		55922 => x"FF",
		55923 => x"FF",
		55924 => x"FF",
		55925 => x"FF",
		55926 => x"FF",
		55927 => x"FF",
		55928 => x"FF",
		55929 => x"FF",
		55930 => x"FF",
		55931 => x"FF",
		55932 => x"FF",
		55933 => x"FF",
		55934 => x"FF",
		55935 => x"FF",
		55936 => x"FF",
		55937 => x"FF",
		55938 => x"FF",
		55939 => x"FF",
		55940 => x"FF",
		55941 => x"FF",
		55942 => x"FF",
		55943 => x"FF",
		55944 => x"FF",
		55945 => x"FF",
		55946 => x"FF",
		55947 => x"FF",
		55948 => x"FF",
		55949 => x"FF",
		55950 => x"FF",
		55951 => x"FF",
		55952 => x"FF",
		55953 => x"FF",
		55954 => x"FF",
		55955 => x"FF",
		55956 => x"FF",
		55957 => x"FF",
		55958 => x"FF",
		55959 => x"FF",
		55960 => x"FF",
		55961 => x"FF",
		55962 => x"FF",
		55963 => x"FF",
		55964 => x"FF",
		55965 => x"FF",
		55966 => x"FF",
		55967 => x"FF",
		55968 => x"FF",
		55969 => x"FF",
		55970 => x"FF",
		55971 => x"FF",
		55972 => x"FF",
		55973 => x"FF",
		55974 => x"FF",
		55975 => x"FF",
		55976 => x"FF",
		55977 => x"FF",
		55978 => x"FF",
		55979 => x"FF",
		55980 => x"FF",
		55981 => x"FF",
		55982 => x"FF",
		55983 => x"FF",
		55984 => x"FF",
		55985 => x"FF",
		55986 => x"FF",
		55987 => x"FF",
		55988 => x"FF",
		55989 => x"FF",
		55990 => x"FF",
		55991 => x"FF",
		55992 => x"FF",
		55993 => x"FF",
		55994 => x"FF",
		55995 => x"FF",
		55996 => x"FF",
		55997 => x"FF",
		55998 => x"FF",
		55999 => x"FF",
		56000 => x"FF",
		56001 => x"FF",
		56002 => x"FF",
		56003 => x"FF",
		56004 => x"FF",
		56005 => x"FF",
		56006 => x"FF",
		56007 => x"FF",
		56008 => x"FF",
		56009 => x"FF",
		56010 => x"FF",
		56011 => x"FF",
		56012 => x"FF",
		56013 => x"FF",
		56014 => x"FF",
		56015 => x"FF",
		56016 => x"FF",
		56017 => x"FF",
		56018 => x"FF",
		56019 => x"FF",
		56020 => x"FF",
		56021 => x"FF",
		56022 => x"FF",
		56023 => x"FF",
		56024 => x"FF",
		56025 => x"FF",
		56026 => x"FF",
