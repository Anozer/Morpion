library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity ROM_vide_sel is
	port (CLK : in std_logic;
		  EN : in std_logic;
		  ADDR : in std_logic_vector(13 downto 0);
		  DATA : out std_logic);
end ROM_vide_sel;

architecture Behavioral of ROM_vide_sel is

type zone_memoire is array ((2**14)-1 downto 0) of std_logic;
constant ROM: zone_memoire := (
		0 => '0',
		1 => '1',
		2 => '0',
		3 => '1',
		4 => '0',
		5 => '1',
		6 => '0',
		7 => '1',
		8 => '0',
		9 => '1',
		10 => '0',
		11 => '1',
		12 => '0',
		13 => '1',
		14 => '0',
		15 => '1',
		16 => '0',
		17 => '1',
		18 => '0',
		19 => '1',
		20 => '0',
		21 => '1',
		22 => '0',
		23 => '1',
		24 => '0',
		25 => '1',
		26 => '0',
		27 => '1',
		28 => '0',
		29 => '1',
		30 => '0',
		31 => '1',
		32 => '0',
		33 => '1',
		34 => '0',
		35 => '1',
		36 => '0',
		37 => '1',
		38 => '0',
		39 => '1',
		40 => '0',
		41 => '1',
		42 => '0',
		43 => '1',
		44 => '0',
		45 => '1',
		46 => '0',
		47 => '1',
		48 => '0',
		49 => '1',
		50 => '0',
		51 => '1',
		52 => '0',
		53 => '1',
		54 => '0',
		55 => '1',
		56 => '0',
		57 => '1',
		58 => '0',
		59 => '1',
		60 => '0',
		61 => '1',
		62 => '0',
		63 => '1',
		64 => '0',
		65 => '1',
		66 => '0',
		67 => '1',
		68 => '0',
		69 => '1',
		70 => '0',
		71 => '1',
		72 => '0',
		73 => '1',
		74 => '0',
		75 => '1',
		76 => '0',
		77 => '1',
		78 => '0',
		79 => '1',
		80 => '0',
		81 => '1',
		82 => '0',
		83 => '1',
		84 => '0',
		85 => '1',
		86 => '0',
		87 => '1',
		88 => '0',
		89 => '1',
		90 => '0',
		91 => '1',
		92 => '0',
		93 => '1',
		94 => '0',
		95 => '1',
		96 => '0',
		97 => '1',
		98 => '0',
		99 => '1',
		100 => '0',
		101 => '1',
		102 => '0',
		103 => '1',
		104 => '0',
		105 => '1',
		106 => '0',
		107 => '1',
		108 => '0',
		109 => '1',
		110 => '0',
		111 => '1',
		112 => '0',
		113 => '1',
		114 => '0',
		115 => '1',
		116 => '0',
		117 => '1',
		118 => '0',
		119 => '1',
		128 => '1',
		129 => '0',
		130 => '1',
		131 => '0',
		132 => '1',
		133 => '0',
		134 => '1',
		135 => '0',
		136 => '1',
		137 => '0',
		138 => '1',
		139 => '0',
		140 => '1',
		141 => '0',
		142 => '1',
		143 => '0',
		144 => '1',
		145 => '0',
		146 => '1',
		147 => '0',
		148 => '1',
		149 => '0',
		150 => '1',
		151 => '0',
		152 => '1',
		153 => '0',
		154 => '1',
		155 => '0',
		156 => '1',
		157 => '0',
		158 => '1',
		159 => '0',
		160 => '1',
		161 => '0',
		162 => '1',
		163 => '0',
		164 => '1',
		165 => '0',
		166 => '1',
		167 => '0',
		168 => '1',
		169 => '0',
		170 => '1',
		171 => '0',
		172 => '1',
		173 => '0',
		174 => '1',
		175 => '0',
		176 => '1',
		177 => '0',
		178 => '1',
		179 => '0',
		180 => '1',
		181 => '0',
		182 => '1',
		183 => '0',
		184 => '1',
		185 => '0',
		186 => '1',
		187 => '0',
		188 => '1',
		189 => '0',
		190 => '1',
		191 => '0',
		192 => '1',
		193 => '0',
		194 => '1',
		195 => '0',
		196 => '1',
		197 => '0',
		198 => '1',
		199 => '0',
		200 => '1',
		201 => '0',
		202 => '1',
		203 => '0',
		204 => '1',
		205 => '0',
		206 => '1',
		207 => '0',
		208 => '1',
		209 => '0',
		210 => '1',
		211 => '0',
		212 => '1',
		213 => '0',
		214 => '1',
		215 => '0',
		216 => '1',
		217 => '0',
		218 => '1',
		219 => '0',
		220 => '1',
		221 => '0',
		222 => '1',
		223 => '0',
		224 => '1',
		225 => '0',
		226 => '1',
		227 => '0',
		228 => '1',
		229 => '0',
		230 => '1',
		231 => '0',
		232 => '1',
		233 => '0',
		234 => '1',
		235 => '0',
		236 => '1',
		237 => '0',
		238 => '1',
		239 => '0',
		240 => '1',
		241 => '0',
		242 => '1',
		243 => '0',
		244 => '1',
		245 => '0',
		246 => '1',
		247 => '0',
		256 => '0',
		257 => '1',
		258 => '0',
		259 => '1',
		260 => '0',
		261 => '1',
		262 => '0',
		263 => '1',
		264 => '0',
		265 => '1',
		266 => '0',
		267 => '1',
		268 => '0',
		269 => '1',
		270 => '0',
		271 => '1',
		272 => '0',
		273 => '1',
		274 => '0',
		275 => '1',
		276 => '0',
		277 => '1',
		278 => '0',
		279 => '1',
		280 => '0',
		281 => '1',
		282 => '0',
		283 => '1',
		284 => '0',
		285 => '1',
		286 => '0',
		287 => '1',
		288 => '0',
		289 => '1',
		290 => '0',
		291 => '1',
		292 => '0',
		293 => '1',
		294 => '0',
		295 => '1',
		296 => '0',
		297 => '1',
		298 => '0',
		299 => '1',
		300 => '0',
		301 => '1',
		302 => '0',
		303 => '1',
		304 => '0',
		305 => '1',
		306 => '0',
		307 => '1',
		308 => '0',
		309 => '1',
		310 => '0',
		311 => '1',
		312 => '0',
		313 => '1',
		314 => '0',
		315 => '1',
		316 => '0',
		317 => '1',
		318 => '0',
		319 => '1',
		320 => '0',
		321 => '1',
		322 => '0',
		323 => '1',
		324 => '0',
		325 => '1',
		326 => '0',
		327 => '1',
		328 => '0',
		329 => '1',
		330 => '0',
		331 => '1',
		332 => '0',
		333 => '1',
		334 => '0',
		335 => '1',
		336 => '0',
		337 => '1',
		338 => '0',
		339 => '1',
		340 => '0',
		341 => '1',
		342 => '0',
		343 => '1',
		344 => '0',
		345 => '1',
		346 => '0',
		347 => '1',
		348 => '0',
		349 => '1',
		350 => '0',
		351 => '1',
		352 => '0',
		353 => '1',
		354 => '0',
		355 => '1',
		356 => '0',
		357 => '1',
		358 => '0',
		359 => '1',
		360 => '0',
		361 => '1',
		362 => '0',
		363 => '1',
		364 => '0',
		365 => '1',
		366 => '0',
		367 => '1',
		368 => '0',
		369 => '1',
		370 => '0',
		371 => '1',
		372 => '0',
		373 => '1',
		374 => '0',
		375 => '1',
		384 => '1',
		385 => '0',
		386 => '1',
		387 => '0',
		388 => '1',
		389 => '0',
		390 => '1',
		391 => '0',
		392 => '1',
		393 => '0',
		394 => '1',
		395 => '0',
		396 => '1',
		397 => '0',
		398 => '1',
		399 => '0',
		400 => '1',
		401 => '0',
		402 => '1',
		403 => '0',
		404 => '1',
		405 => '0',
		406 => '1',
		407 => '0',
		408 => '1',
		409 => '0',
		410 => '1',
		411 => '0',
		412 => '1',
		413 => '0',
		414 => '1',
		415 => '0',
		416 => '1',
		417 => '0',
		418 => '1',
		419 => '0',
		420 => '1',
		421 => '0',
		422 => '1',
		423 => '0',
		424 => '1',
		425 => '0',
		426 => '1',
		427 => '0',
		428 => '1',
		429 => '0',
		430 => '1',
		431 => '0',
		432 => '1',
		433 => '0',
		434 => '1',
		435 => '0',
		436 => '1',
		437 => '0',
		438 => '1',
		439 => '0',
		440 => '1',
		441 => '0',
		442 => '1',
		443 => '0',
		444 => '1',
		445 => '0',
		446 => '1',
		447 => '0',
		448 => '1',
		449 => '0',
		450 => '1',
		451 => '0',
		452 => '1',
		453 => '0',
		454 => '1',
		455 => '0',
		456 => '1',
		457 => '0',
		458 => '1',
		459 => '0',
		460 => '1',
		461 => '0',
		462 => '1',
		463 => '0',
		464 => '1',
		465 => '0',
		466 => '1',
		467 => '0',
		468 => '1',
		469 => '0',
		470 => '1',
		471 => '0',
		472 => '1',
		473 => '0',
		474 => '1',
		475 => '0',
		476 => '1',
		477 => '0',
		478 => '1',
		479 => '0',
		480 => '1',
		481 => '0',
		482 => '1',
		483 => '0',
		484 => '1',
		485 => '0',
		486 => '1',
		487 => '0',
		488 => '1',
		489 => '0',
		490 => '1',
		491 => '0',
		492 => '1',
		493 => '0',
		494 => '1',
		495 => '0',
		496 => '1',
		497 => '0',
		498 => '1',
		499 => '0',
		500 => '1',
		501 => '0',
		502 => '1',
		503 => '0',
		512 => '0',
		513 => '1',
		514 => '0',
		515 => '1',
		516 => '0',
		517 => '1',
		518 => '0',
		519 => '1',
		520 => '0',
		521 => '1',
		522 => '0',
		523 => '1',
		524 => '0',
		525 => '1',
		526 => '0',
		527 => '1',
		528 => '0',
		529 => '1',
		530 => '0',
		531 => '1',
		532 => '0',
		533 => '1',
		534 => '0',
		535 => '1',
		536 => '0',
		537 => '1',
		538 => '0',
		539 => '1',
		540 => '0',
		541 => '1',
		542 => '0',
		543 => '1',
		544 => '0',
		545 => '1',
		546 => '0',
		547 => '1',
		548 => '0',
		549 => '1',
		550 => '0',
		551 => '1',
		552 => '0',
		553 => '1',
		554 => '0',
		555 => '1',
		556 => '0',
		557 => '1',
		558 => '0',
		559 => '1',
		560 => '0',
		561 => '1',
		562 => '0',
		563 => '1',
		564 => '0',
		565 => '1',
		566 => '0',
		567 => '1',
		568 => '0',
		569 => '1',
		570 => '0',
		571 => '1',
		572 => '0',
		573 => '1',
		574 => '0',
		575 => '1',
		576 => '0',
		577 => '1',
		578 => '0',
		579 => '1',
		580 => '0',
		581 => '1',
		582 => '0',
		583 => '1',
		584 => '0',
		585 => '1',
		586 => '0',
		587 => '1',
		588 => '0',
		589 => '1',
		590 => '0',
		591 => '1',
		592 => '0',
		593 => '1',
		594 => '0',
		595 => '1',
		596 => '0',
		597 => '1',
		598 => '0',
		599 => '1',
		600 => '0',
		601 => '1',
		602 => '0',
		603 => '1',
		604 => '0',
		605 => '1',
		606 => '0',
		607 => '1',
		608 => '0',
		609 => '1',
		610 => '0',
		611 => '1',
		612 => '0',
		613 => '1',
		614 => '0',
		615 => '1',
		616 => '0',
		617 => '1',
		618 => '0',
		619 => '1',
		620 => '0',
		621 => '1',
		622 => '0',
		623 => '1',
		624 => '0',
		625 => '1',
		626 => '0',
		627 => '1',
		628 => '0',
		629 => '1',
		630 => '0',
		631 => '1',
		640 => '1',
		641 => '0',
		642 => '1',
		643 => '0',
		644 => '1',
		645 => '0',
		646 => '1',
		647 => '0',
		648 => '1',
		649 => '0',
		650 => '1',
		651 => '0',
		652 => '1',
		653 => '0',
		654 => '1',
		655 => '0',
		656 => '1',
		657 => '0',
		658 => '1',
		659 => '0',
		660 => '1',
		661 => '0',
		662 => '1',
		663 => '0',
		664 => '1',
		665 => '0',
		666 => '1',
		667 => '0',
		668 => '1',
		669 => '0',
		670 => '1',
		671 => '0',
		672 => '1',
		673 => '0',
		674 => '1',
		675 => '0',
		676 => '1',
		677 => '0',
		678 => '1',
		679 => '0',
		680 => '1',
		681 => '0',
		682 => '1',
		683 => '0',
		684 => '1',
		685 => '0',
		686 => '1',
		687 => '0',
		688 => '1',
		689 => '0',
		690 => '1',
		691 => '0',
		692 => '1',
		693 => '0',
		694 => '1',
		695 => '0',
		696 => '1',
		697 => '0',
		698 => '1',
		699 => '0',
		700 => '1',
		701 => '0',
		702 => '1',
		703 => '0',
		704 => '1',
		705 => '0',
		706 => '1',
		707 => '0',
		708 => '1',
		709 => '0',
		710 => '1',
		711 => '0',
		712 => '1',
		713 => '0',
		714 => '1',
		715 => '0',
		716 => '1',
		717 => '0',
		718 => '1',
		719 => '0',
		720 => '1',
		721 => '0',
		722 => '1',
		723 => '0',
		724 => '1',
		725 => '0',
		726 => '1',
		727 => '0',
		728 => '1',
		729 => '0',
		730 => '1',
		731 => '0',
		732 => '1',
		733 => '0',
		734 => '1',
		735 => '0',
		736 => '1',
		737 => '0',
		738 => '1',
		739 => '0',
		740 => '1',
		741 => '0',
		742 => '1',
		743 => '0',
		744 => '1',
		745 => '0',
		746 => '1',
		747 => '0',
		748 => '1',
		749 => '0',
		750 => '1',
		751 => '0',
		752 => '1',
		753 => '0',
		754 => '1',
		755 => '0',
		756 => '1',
		757 => '0',
		758 => '1',
		759 => '0',
		768 => '0',
		769 => '1',
		770 => '0',
		771 => '1',
		772 => '0',
		773 => '1',
		774 => '0',
		775 => '1',
		776 => '0',
		777 => '1',
		778 => '0',
		779 => '1',
		780 => '0',
		781 => '1',
		782 => '0',
		783 => '1',
		784 => '0',
		785 => '1',
		786 => '0',
		787 => '1',
		788 => '0',
		789 => '1',
		790 => '0',
		791 => '1',
		792 => '0',
		793 => '1',
		794 => '0',
		795 => '1',
		796 => '0',
		797 => '1',
		798 => '0',
		799 => '1',
		800 => '0',
		801 => '1',
		802 => '0',
		803 => '1',
		804 => '0',
		805 => '1',
		806 => '0',
		807 => '1',
		808 => '0',
		809 => '1',
		810 => '0',
		811 => '1',
		812 => '0',
		813 => '1',
		814 => '0',
		815 => '1',
		816 => '0',
		817 => '1',
		818 => '0',
		819 => '1',
		820 => '0',
		821 => '1',
		822 => '0',
		823 => '1',
		824 => '0',
		825 => '1',
		826 => '0',
		827 => '1',
		828 => '0',
		829 => '1',
		830 => '0',
		831 => '1',
		832 => '0',
		833 => '1',
		834 => '0',
		835 => '1',
		836 => '0',
		837 => '1',
		838 => '0',
		839 => '1',
		840 => '0',
		841 => '1',
		842 => '0',
		843 => '1',
		844 => '0',
		845 => '1',
		846 => '0',
		847 => '1',
		848 => '0',
		849 => '1',
		850 => '0',
		851 => '1',
		852 => '0',
		853 => '1',
		854 => '0',
		855 => '1',
		856 => '0',
		857 => '1',
		858 => '0',
		859 => '1',
		860 => '0',
		861 => '1',
		862 => '0',
		863 => '1',
		864 => '0',
		865 => '1',
		866 => '0',
		867 => '1',
		868 => '0',
		869 => '1',
		870 => '0',
		871 => '1',
		872 => '0',
		873 => '1',
		874 => '0',
		875 => '1',
		876 => '0',
		877 => '1',
		878 => '0',
		879 => '1',
		880 => '0',
		881 => '1',
		882 => '0',
		883 => '1',
		884 => '0',
		885 => '1',
		886 => '0',
		887 => '1',
		896 => '1',
		897 => '0',
		898 => '1',
		899 => '0',
		900 => '1',
		901 => '0',
		902 => '1',
		903 => '0',
		904 => '1',
		905 => '0',
		906 => '1',
		907 => '0',
		908 => '1',
		909 => '0',
		910 => '1',
		911 => '0',
		912 => '1',
		913 => '0',
		914 => '1',
		915 => '0',
		916 => '1',
		917 => '0',
		918 => '1',
		919 => '0',
		920 => '1',
		921 => '0',
		922 => '1',
		923 => '0',
		924 => '1',
		925 => '0',
		926 => '1',
		927 => '0',
		928 => '1',
		929 => '0',
		930 => '1',
		931 => '0',
		932 => '1',
		933 => '0',
		934 => '1',
		935 => '0',
		936 => '1',
		937 => '0',
		938 => '1',
		939 => '0',
		940 => '1',
		941 => '0',
		942 => '1',
		943 => '0',
		944 => '1',
		945 => '0',
		946 => '1',
		947 => '0',
		948 => '1',
		949 => '0',
		950 => '1',
		951 => '0',
		952 => '1',
		953 => '0',
		954 => '1',
		955 => '0',
		956 => '1',
		957 => '0',
		958 => '1',
		959 => '0',
		960 => '1',
		961 => '0',
		962 => '1',
		963 => '0',
		964 => '1',
		965 => '0',
		966 => '1',
		967 => '0',
		968 => '1',
		969 => '0',
		970 => '1',
		971 => '0',
		972 => '1',
		973 => '0',
		974 => '1',
		975 => '0',
		976 => '1',
		977 => '0',
		978 => '1',
		979 => '0',
		980 => '1',
		981 => '0',
		982 => '1',
		983 => '0',
		984 => '1',
		985 => '0',
		986 => '1',
		987 => '0',
		988 => '1',
		989 => '0',
		990 => '1',
		991 => '0',
		992 => '1',
		993 => '0',
		994 => '1',
		995 => '0',
		996 => '1',
		997 => '0',
		998 => '1',
		999 => '0',
		1000 => '1',
		1001 => '0',
		1002 => '1',
		1003 => '0',
		1004 => '1',
		1005 => '0',
		1006 => '1',
		1007 => '0',
		1008 => '1',
		1009 => '0',
		1010 => '1',
		1011 => '0',
		1012 => '1',
		1013 => '0',
		1014 => '1',
		1015 => '0',
		1024 => '0',
		1025 => '1',
		1026 => '0',
		1027 => '1',
		1028 => '0',
		1029 => '1',
		1030 => '0',
		1031 => '1',
		1032 => '0',
		1033 => '1',
		1034 => '0',
		1035 => '1',
		1036 => '0',
		1037 => '1',
		1038 => '0',
		1039 => '1',
		1040 => '0',
		1041 => '1',
		1042 => '0',
		1043 => '1',
		1044 => '0',
		1045 => '1',
		1046 => '0',
		1047 => '1',
		1048 => '0',
		1049 => '1',
		1050 => '0',
		1051 => '1',
		1052 => '0',
		1053 => '1',
		1054 => '0',
		1055 => '1',
		1056 => '0',
		1057 => '1',
		1058 => '0',
		1059 => '1',
		1060 => '0',
		1061 => '1',
		1062 => '0',
		1063 => '1',
		1064 => '0',
		1065 => '1',
		1066 => '0',
		1067 => '1',
		1068 => '0',
		1069 => '1',
		1070 => '0',
		1071 => '1',
		1072 => '0',
		1073 => '1',
		1074 => '0',
		1075 => '1',
		1076 => '0',
		1077 => '1',
		1078 => '0',
		1079 => '1',
		1080 => '0',
		1081 => '1',
		1082 => '0',
		1083 => '1',
		1084 => '0',
		1085 => '1',
		1086 => '0',
		1087 => '1',
		1088 => '0',
		1089 => '1',
		1090 => '0',
		1091 => '1',
		1092 => '0',
		1093 => '1',
		1094 => '0',
		1095 => '1',
		1096 => '0',
		1097 => '1',
		1098 => '0',
		1099 => '1',
		1100 => '0',
		1101 => '1',
		1102 => '0',
		1103 => '1',
		1104 => '0',
		1105 => '1',
		1106 => '0',
		1107 => '1',
		1108 => '0',
		1109 => '1',
		1110 => '0',
		1111 => '1',
		1112 => '0',
		1113 => '1',
		1114 => '0',
		1115 => '1',
		1116 => '0',
		1117 => '1',
		1118 => '0',
		1119 => '1',
		1120 => '0',
		1121 => '1',
		1122 => '0',
		1123 => '1',
		1124 => '0',
		1125 => '1',
		1126 => '0',
		1127 => '1',
		1128 => '0',
		1129 => '1',
		1130 => '0',
		1131 => '1',
		1132 => '0',
		1133 => '1',
		1134 => '0',
		1135 => '1',
		1136 => '0',
		1137 => '1',
		1138 => '0',
		1139 => '1',
		1140 => '0',
		1141 => '1',
		1142 => '0',
		1143 => '1',
		1152 => '1',
		1153 => '0',
		1154 => '1',
		1155 => '0',
		1156 => '1',
		1157 => '0',
		1158 => '1',
		1159 => '0',
		1160 => '1',
		1161 => '0',
		1162 => '1',
		1163 => '0',
		1164 => '1',
		1165 => '0',
		1166 => '1',
		1167 => '0',
		1168 => '1',
		1169 => '0',
		1170 => '1',
		1171 => '0',
		1172 => '1',
		1173 => '0',
		1174 => '1',
		1175 => '0',
		1176 => '1',
		1177 => '0',
		1178 => '1',
		1179 => '0',
		1180 => '1',
		1181 => '0',
		1182 => '1',
		1183 => '0',
		1184 => '1',
		1185 => '0',
		1186 => '1',
		1187 => '0',
		1188 => '1',
		1189 => '0',
		1190 => '1',
		1191 => '0',
		1192 => '1',
		1193 => '0',
		1194 => '1',
		1195 => '0',
		1196 => '1',
		1197 => '0',
		1198 => '1',
		1199 => '0',
		1200 => '1',
		1201 => '0',
		1202 => '1',
		1203 => '0',
		1204 => '1',
		1205 => '0',
		1206 => '1',
		1207 => '0',
		1208 => '1',
		1209 => '0',
		1210 => '1',
		1211 => '0',
		1212 => '1',
		1213 => '0',
		1214 => '1',
		1215 => '0',
		1216 => '1',
		1217 => '0',
		1218 => '1',
		1219 => '0',
		1220 => '1',
		1221 => '0',
		1222 => '1',
		1223 => '0',
		1224 => '1',
		1225 => '0',
		1226 => '1',
		1227 => '0',
		1228 => '1',
		1229 => '0',
		1230 => '1',
		1231 => '0',
		1232 => '1',
		1233 => '0',
		1234 => '1',
		1235 => '0',
		1236 => '1',
		1237 => '0',
		1238 => '1',
		1239 => '0',
		1240 => '1',
		1241 => '0',
		1242 => '1',
		1243 => '0',
		1244 => '1',
		1245 => '0',
		1246 => '1',
		1247 => '0',
		1248 => '1',
		1249 => '0',
		1250 => '1',
		1251 => '0',
		1252 => '1',
		1253 => '0',
		1254 => '1',
		1255 => '0',
		1256 => '1',
		1257 => '0',
		1258 => '1',
		1259 => '0',
		1260 => '1',
		1261 => '0',
		1262 => '1',
		1263 => '0',
		1264 => '1',
		1265 => '0',
		1266 => '1',
		1267 => '0',
		1268 => '1',
		1269 => '0',
		1270 => '1',
		1271 => '0',
		1280 => '0',
		1281 => '1',
		1282 => '0',
		1283 => '1',
		1284 => '0',
		1285 => '1',
		1286 => '0',
		1287 => '1',
		1288 => '0',
		1289 => '1',
		1290 => '0',
		1291 => '1',
		1292 => '0',
		1293 => '1',
		1294 => '0',
		1295 => '1',
		1296 => '0',
		1297 => '1',
		1298 => '0',
		1299 => '1',
		1300 => '0',
		1301 => '1',
		1302 => '0',
		1303 => '1',
		1304 => '0',
		1305 => '1',
		1306 => '0',
		1307 => '1',
		1308 => '0',
		1309 => '1',
		1310 => '0',
		1311 => '1',
		1312 => '0',
		1313 => '1',
		1314 => '0',
		1315 => '1',
		1316 => '0',
		1317 => '1',
		1318 => '0',
		1319 => '1',
		1320 => '0',
		1321 => '1',
		1322 => '0',
		1323 => '1',
		1324 => '0',
		1325 => '1',
		1326 => '0',
		1327 => '1',
		1328 => '0',
		1329 => '1',
		1330 => '0',
		1331 => '1',
		1332 => '0',
		1333 => '1',
		1334 => '0',
		1335 => '1',
		1336 => '0',
		1337 => '1',
		1338 => '0',
		1339 => '1',
		1340 => '0',
		1341 => '1',
		1342 => '0',
		1343 => '1',
		1344 => '0',
		1345 => '1',
		1346 => '0',
		1347 => '1',
		1348 => '0',
		1349 => '1',
		1350 => '0',
		1351 => '1',
		1352 => '0',
		1353 => '1',
		1354 => '0',
		1355 => '1',
		1356 => '0',
		1357 => '1',
		1358 => '0',
		1359 => '1',
		1360 => '0',
		1361 => '1',
		1362 => '0',
		1363 => '1',
		1364 => '0',
		1365 => '1',
		1366 => '0',
		1367 => '1',
		1368 => '0',
		1369 => '1',
		1370 => '0',
		1371 => '1',
		1372 => '0',
		1373 => '1',
		1374 => '0',
		1375 => '1',
		1376 => '0',
		1377 => '1',
		1378 => '0',
		1379 => '1',
		1380 => '0',
		1381 => '1',
		1382 => '0',
		1383 => '1',
		1384 => '0',
		1385 => '1',
		1386 => '0',
		1387 => '1',
		1388 => '0',
		1389 => '1',
		1390 => '0',
		1391 => '1',
		1392 => '0',
		1393 => '1',
		1394 => '0',
		1395 => '1',
		1396 => '0',
		1397 => '1',
		1398 => '0',
		1399 => '1',
		1408 => '1',
		1409 => '0',
		1410 => '1',
		1411 => '0',
		1412 => '1',
		1413 => '0',
		1414 => '1',
		1415 => '0',
		1416 => '1',
		1417 => '0',
		1418 => '1',
		1419 => '0',
		1420 => '1',
		1421 => '0',
		1422 => '1',
		1423 => '0',
		1424 => '1',
		1425 => '0',
		1426 => '1',
		1427 => '0',
		1428 => '1',
		1429 => '0',
		1430 => '1',
		1431 => '0',
		1432 => '1',
		1433 => '0',
		1434 => '1',
		1435 => '0',
		1436 => '1',
		1437 => '0',
		1438 => '1',
		1439 => '0',
		1440 => '1',
		1441 => '0',
		1442 => '1',
		1443 => '0',
		1444 => '1',
		1445 => '0',
		1446 => '1',
		1447 => '0',
		1448 => '1',
		1449 => '0',
		1450 => '1',
		1451 => '0',
		1452 => '1',
		1453 => '0',
		1454 => '1',
		1455 => '0',
		1456 => '1',
		1457 => '0',
		1458 => '1',
		1459 => '0',
		1460 => '1',
		1461 => '0',
		1462 => '1',
		1463 => '0',
		1464 => '1',
		1465 => '0',
		1466 => '1',
		1467 => '0',
		1468 => '1',
		1469 => '0',
		1470 => '1',
		1471 => '0',
		1472 => '1',
		1473 => '0',
		1474 => '1',
		1475 => '0',
		1476 => '1',
		1477 => '0',
		1478 => '1',
		1479 => '0',
		1480 => '1',
		1481 => '0',
		1482 => '1',
		1483 => '0',
		1484 => '1',
		1485 => '0',
		1486 => '1',
		1487 => '0',
		1488 => '1',
		1489 => '0',
		1490 => '1',
		1491 => '0',
		1492 => '1',
		1493 => '0',
		1494 => '1',
		1495 => '0',
		1496 => '1',
		1497 => '0',
		1498 => '1',
		1499 => '0',
		1500 => '1',
		1501 => '0',
		1502 => '1',
		1503 => '0',
		1504 => '1',
		1505 => '0',
		1506 => '1',
		1507 => '0',
		1508 => '1',
		1509 => '0',
		1510 => '1',
		1511 => '0',
		1512 => '1',
		1513 => '0',
		1514 => '1',
		1515 => '0',
		1516 => '1',
		1517 => '0',
		1518 => '1',
		1519 => '0',
		1520 => '1',
		1521 => '0',
		1522 => '1',
		1523 => '0',
		1524 => '1',
		1525 => '0',
		1526 => '1',
		1527 => '0',
		1536 => '0',
		1537 => '1',
		1538 => '0',
		1539 => '1',
		1540 => '0',
		1541 => '1',
		1542 => '0',
		1543 => '1',
		1544 => '0',
		1545 => '1',
		1546 => '0',
		1547 => '1',
		1548 => '0',
		1549 => '1',
		1550 => '0',
		1551 => '1',
		1552 => '0',
		1553 => '1',
		1554 => '0',
		1555 => '1',
		1556 => '0',
		1557 => '1',
		1558 => '0',
		1559 => '1',
		1560 => '0',
		1561 => '1',
		1562 => '0',
		1563 => '1',
		1564 => '0',
		1565 => '1',
		1566 => '0',
		1567 => '1',
		1568 => '0',
		1569 => '1',
		1570 => '0',
		1571 => '1',
		1572 => '0',
		1573 => '1',
		1574 => '0',
		1575 => '1',
		1576 => '0',
		1577 => '1',
		1578 => '0',
		1579 => '1',
		1580 => '0',
		1581 => '1',
		1582 => '0',
		1583 => '1',
		1584 => '0',
		1585 => '1',
		1586 => '0',
		1587 => '1',
		1588 => '0',
		1589 => '1',
		1590 => '0',
		1591 => '1',
		1592 => '0',
		1593 => '1',
		1594 => '0',
		1595 => '1',
		1596 => '0',
		1597 => '1',
		1598 => '0',
		1599 => '1',
		1600 => '0',
		1601 => '1',
		1602 => '0',
		1603 => '1',
		1604 => '0',
		1605 => '1',
		1606 => '0',
		1607 => '1',
		1608 => '0',
		1609 => '1',
		1610 => '0',
		1611 => '1',
		1612 => '0',
		1613 => '1',
		1614 => '0',
		1615 => '1',
		1616 => '0',
		1617 => '1',
		1618 => '0',
		1619 => '1',
		1620 => '0',
		1621 => '1',
		1622 => '0',
		1623 => '1',
		1624 => '0',
		1625 => '1',
		1626 => '0',
		1627 => '1',
		1628 => '0',
		1629 => '1',
		1630 => '0',
		1631 => '1',
		1632 => '0',
		1633 => '1',
		1634 => '0',
		1635 => '1',
		1636 => '0',
		1637 => '1',
		1638 => '0',
		1639 => '1',
		1640 => '0',
		1641 => '1',
		1642 => '0',
		1643 => '1',
		1644 => '0',
		1645 => '1',
		1646 => '0',
		1647 => '1',
		1648 => '0',
		1649 => '1',
		1650 => '0',
		1651 => '1',
		1652 => '0',
		1653 => '1',
		1654 => '0',
		1655 => '1',
		1664 => '1',
		1665 => '0',
		1666 => '1',
		1667 => '0',
		1668 => '1',
		1669 => '0',
		1670 => '1',
		1671 => '0',
		1672 => '1',
		1673 => '0',
		1674 => '1',
		1675 => '0',
		1676 => '1',
		1677 => '0',
		1678 => '1',
		1679 => '0',
		1680 => '1',
		1681 => '0',
		1682 => '1',
		1683 => '0',
		1684 => '1',
		1685 => '0',
		1686 => '1',
		1687 => '0',
		1688 => '1',
		1689 => '0',
		1690 => '1',
		1691 => '0',
		1692 => '1',
		1693 => '0',
		1694 => '1',
		1695 => '0',
		1696 => '1',
		1697 => '0',
		1698 => '1',
		1699 => '0',
		1700 => '1',
		1701 => '0',
		1702 => '1',
		1703 => '0',
		1704 => '1',
		1705 => '0',
		1706 => '1',
		1707 => '0',
		1708 => '1',
		1709 => '0',
		1710 => '1',
		1711 => '0',
		1712 => '1',
		1713 => '0',
		1714 => '1',
		1715 => '0',
		1716 => '1',
		1717 => '0',
		1718 => '1',
		1719 => '0',
		1720 => '1',
		1721 => '0',
		1722 => '1',
		1723 => '0',
		1724 => '1',
		1725 => '0',
		1726 => '1',
		1727 => '0',
		1728 => '1',
		1729 => '0',
		1730 => '1',
		1731 => '0',
		1732 => '1',
		1733 => '0',
		1734 => '1',
		1735 => '0',
		1736 => '1',
		1737 => '0',
		1738 => '1',
		1739 => '0',
		1740 => '1',
		1741 => '0',
		1742 => '1',
		1743 => '0',
		1744 => '1',
		1745 => '0',
		1746 => '1',
		1747 => '0',
		1748 => '1',
		1749 => '0',
		1750 => '1',
		1751 => '0',
		1752 => '1',
		1753 => '0',
		1754 => '1',
		1755 => '0',
		1756 => '1',
		1757 => '0',
		1758 => '1',
		1759 => '0',
		1760 => '1',
		1761 => '0',
		1762 => '1',
		1763 => '0',
		1764 => '1',
		1765 => '0',
		1766 => '1',
		1767 => '0',
		1768 => '1',
		1769 => '0',
		1770 => '1',
		1771 => '0',
		1772 => '1',
		1773 => '0',
		1774 => '1',
		1775 => '0',
		1776 => '1',
		1777 => '0',
		1778 => '1',
		1779 => '0',
		1780 => '1',
		1781 => '0',
		1782 => '1',
		1783 => '0',
		1792 => '0',
		1793 => '1',
		1794 => '0',
		1795 => '1',
		1796 => '0',
		1797 => '1',
		1798 => '0',
		1799 => '1',
		1800 => '0',
		1801 => '1',
		1802 => '0',
		1803 => '1',
		1804 => '0',
		1805 => '1',
		1806 => '0',
		1807 => '1',
		1808 => '0',
		1809 => '1',
		1810 => '0',
		1811 => '1',
		1812 => '0',
		1813 => '1',
		1814 => '0',
		1815 => '1',
		1816 => '0',
		1817 => '1',
		1818 => '0',
		1819 => '1',
		1820 => '0',
		1821 => '1',
		1822 => '0',
		1823 => '1',
		1824 => '0',
		1825 => '1',
		1826 => '0',
		1827 => '1',
		1828 => '0',
		1829 => '1',
		1830 => '0',
		1831 => '1',
		1832 => '0',
		1833 => '1',
		1834 => '0',
		1835 => '1',
		1836 => '0',
		1837 => '1',
		1838 => '0',
		1839 => '1',
		1840 => '0',
		1841 => '1',
		1842 => '0',
		1843 => '1',
		1844 => '0',
		1845 => '1',
		1846 => '0',
		1847 => '1',
		1848 => '0',
		1849 => '1',
		1850 => '0',
		1851 => '1',
		1852 => '0',
		1853 => '1',
		1854 => '0',
		1855 => '1',
		1856 => '0',
		1857 => '1',
		1858 => '0',
		1859 => '1',
		1860 => '0',
		1861 => '1',
		1862 => '0',
		1863 => '1',
		1864 => '0',
		1865 => '1',
		1866 => '0',
		1867 => '1',
		1868 => '0',
		1869 => '1',
		1870 => '0',
		1871 => '1',
		1872 => '0',
		1873 => '1',
		1874 => '0',
		1875 => '1',
		1876 => '0',
		1877 => '1',
		1878 => '0',
		1879 => '1',
		1880 => '0',
		1881 => '1',
		1882 => '0',
		1883 => '1',
		1884 => '0',
		1885 => '1',
		1886 => '0',
		1887 => '1',
		1888 => '0',
		1889 => '1',
		1890 => '0',
		1891 => '1',
		1892 => '0',
		1893 => '1',
		1894 => '0',
		1895 => '1',
		1896 => '0',
		1897 => '1',
		1898 => '0',
		1899 => '1',
		1900 => '0',
		1901 => '1',
		1902 => '0',
		1903 => '1',
		1904 => '0',
		1905 => '1',
		1906 => '0',
		1907 => '1',
		1908 => '0',
		1909 => '1',
		1910 => '0',
		1911 => '1',
		1920 => '1',
		1921 => '0',
		1922 => '1',
		1923 => '0',
		1924 => '1',
		1925 => '0',
		1926 => '1',
		1927 => '0',
		1928 => '1',
		1929 => '0',
		1930 => '1',
		1931 => '0',
		1932 => '1',
		1933 => '0',
		1934 => '1',
		1935 => '0',
		1936 => '1',
		1937 => '0',
		1938 => '1',
		1939 => '0',
		1940 => '1',
		1941 => '0',
		1942 => '1',
		1943 => '0',
		1944 => '1',
		1945 => '0',
		1946 => '1',
		1947 => '0',
		1948 => '1',
		1949 => '0',
		1950 => '1',
		1951 => '0',
		1952 => '1',
		1953 => '0',
		1954 => '1',
		1955 => '0',
		1956 => '1',
		1957 => '0',
		1958 => '1',
		1959 => '0',
		1960 => '1',
		1961 => '0',
		1962 => '1',
		1963 => '0',
		1964 => '1',
		1965 => '0',
		1966 => '1',
		1967 => '0',
		1968 => '1',
		1969 => '0',
		1970 => '1',
		1971 => '0',
		1972 => '1',
		1973 => '0',
		1974 => '1',
		1975 => '0',
		1976 => '1',
		1977 => '0',
		1978 => '1',
		1979 => '0',
		1980 => '1',
		1981 => '0',
		1982 => '1',
		1983 => '0',
		1984 => '1',
		1985 => '0',
		1986 => '1',
		1987 => '0',
		1988 => '1',
		1989 => '0',
		1990 => '1',
		1991 => '0',
		1992 => '1',
		1993 => '0',
		1994 => '1',
		1995 => '0',
		1996 => '1',
		1997 => '0',
		1998 => '1',
		1999 => '0',
		2000 => '1',
		2001 => '0',
		2002 => '1',
		2003 => '0',
		2004 => '1',
		2005 => '0',
		2006 => '1',
		2007 => '0',
		2008 => '1',
		2009 => '0',
		2010 => '1',
		2011 => '0',
		2012 => '1',
		2013 => '0',
		2014 => '1',
		2015 => '0',
		2016 => '1',
		2017 => '0',
		2018 => '1',
		2019 => '0',
		2020 => '1',
		2021 => '0',
		2022 => '1',
		2023 => '0',
		2024 => '1',
		2025 => '0',
		2026 => '1',
		2027 => '0',
		2028 => '1',
		2029 => '0',
		2030 => '1',
		2031 => '0',
		2032 => '1',
		2033 => '0',
		2034 => '1',
		2035 => '0',
		2036 => '1',
		2037 => '0',
		2038 => '1',
		2039 => '0',
		2048 => '0',
		2049 => '1',
		2050 => '0',
		2051 => '1',
		2052 => '0',
		2053 => '1',
		2054 => '0',
		2055 => '1',
		2056 => '0',
		2057 => '1',
		2058 => '0',
		2059 => '1',
		2060 => '0',
		2061 => '1',
		2062 => '0',
		2063 => '1',
		2064 => '0',
		2065 => '1',
		2066 => '0',
		2067 => '1',
		2068 => '0',
		2069 => '1',
		2070 => '0',
		2071 => '1',
		2072 => '0',
		2073 => '1',
		2074 => '0',
		2075 => '1',
		2076 => '0',
		2077 => '1',
		2078 => '0',
		2079 => '1',
		2080 => '0',
		2081 => '1',
		2082 => '0',
		2083 => '1',
		2084 => '0',
		2085 => '1',
		2086 => '0',
		2087 => '1',
		2088 => '0',
		2089 => '1',
		2090 => '0',
		2091 => '1',
		2092 => '0',
		2093 => '1',
		2094 => '0',
		2095 => '1',
		2096 => '0',
		2097 => '1',
		2098 => '0',
		2099 => '1',
		2100 => '0',
		2101 => '1',
		2102 => '0',
		2103 => '1',
		2104 => '0',
		2105 => '1',
		2106 => '0',
		2107 => '1',
		2108 => '0',
		2109 => '1',
		2110 => '0',
		2111 => '1',
		2112 => '0',
		2113 => '1',
		2114 => '0',
		2115 => '1',
		2116 => '0',
		2117 => '1',
		2118 => '0',
		2119 => '1',
		2120 => '0',
		2121 => '1',
		2122 => '0',
		2123 => '1',
		2124 => '0',
		2125 => '1',
		2126 => '0',
		2127 => '1',
		2128 => '0',
		2129 => '1',
		2130 => '0',
		2131 => '1',
		2132 => '0',
		2133 => '1',
		2134 => '0',
		2135 => '1',
		2136 => '0',
		2137 => '1',
		2138 => '0',
		2139 => '1',
		2140 => '0',
		2141 => '1',
		2142 => '0',
		2143 => '1',
		2144 => '0',
		2145 => '1',
		2146 => '0',
		2147 => '1',
		2148 => '0',
		2149 => '1',
		2150 => '0',
		2151 => '1',
		2152 => '0',
		2153 => '1',
		2154 => '0',
		2155 => '1',
		2156 => '0',
		2157 => '1',
		2158 => '0',
		2159 => '1',
		2160 => '0',
		2161 => '1',
		2162 => '0',
		2163 => '1',
		2164 => '0',
		2165 => '1',
		2166 => '0',
		2167 => '1',
		2176 => '1',
		2177 => '0',
		2178 => '1',
		2179 => '0',
		2180 => '1',
		2181 => '0',
		2182 => '1',
		2183 => '0',
		2184 => '1',
		2185 => '0',
		2186 => '1',
		2187 => '0',
		2188 => '1',
		2189 => '0',
		2190 => '1',
		2191 => '0',
		2192 => '1',
		2193 => '0',
		2194 => '1',
		2195 => '0',
		2196 => '1',
		2197 => '0',
		2198 => '1',
		2199 => '0',
		2200 => '1',
		2201 => '0',
		2202 => '1',
		2203 => '0',
		2204 => '1',
		2205 => '0',
		2206 => '1',
		2207 => '0',
		2208 => '1',
		2209 => '0',
		2210 => '1',
		2211 => '0',
		2212 => '1',
		2213 => '0',
		2214 => '1',
		2215 => '0',
		2216 => '1',
		2217 => '0',
		2218 => '1',
		2219 => '0',
		2220 => '1',
		2221 => '0',
		2222 => '1',
		2223 => '0',
		2224 => '1',
		2225 => '0',
		2226 => '1',
		2227 => '0',
		2228 => '1',
		2229 => '0',
		2230 => '1',
		2231 => '0',
		2232 => '1',
		2233 => '0',
		2234 => '1',
		2235 => '0',
		2236 => '1',
		2237 => '0',
		2238 => '1',
		2239 => '0',
		2240 => '1',
		2241 => '0',
		2242 => '1',
		2243 => '0',
		2244 => '1',
		2245 => '0',
		2246 => '1',
		2247 => '0',
		2248 => '1',
		2249 => '0',
		2250 => '1',
		2251 => '0',
		2252 => '1',
		2253 => '0',
		2254 => '1',
		2255 => '0',
		2256 => '1',
		2257 => '0',
		2258 => '1',
		2259 => '0',
		2260 => '1',
		2261 => '0',
		2262 => '1',
		2263 => '0',
		2264 => '1',
		2265 => '0',
		2266 => '1',
		2267 => '0',
		2268 => '1',
		2269 => '0',
		2270 => '1',
		2271 => '0',
		2272 => '1',
		2273 => '0',
		2274 => '1',
		2275 => '0',
		2276 => '1',
		2277 => '0',
		2278 => '1',
		2279 => '0',
		2280 => '1',
		2281 => '0',
		2282 => '1',
		2283 => '0',
		2284 => '1',
		2285 => '0',
		2286 => '1',
		2287 => '0',
		2288 => '1',
		2289 => '0',
		2290 => '1',
		2291 => '0',
		2292 => '1',
		2293 => '0',
		2294 => '1',
		2295 => '0',
		2304 => '0',
		2305 => '1',
		2306 => '0',
		2307 => '1',
		2308 => '0',
		2309 => '1',
		2310 => '0',
		2311 => '1',
		2312 => '0',
		2313 => '1',
		2314 => '0',
		2315 => '1',
		2316 => '0',
		2317 => '1',
		2318 => '0',
		2319 => '1',
		2320 => '0',
		2321 => '1',
		2322 => '0',
		2323 => '1',
		2324 => '0',
		2325 => '1',
		2326 => '0',
		2327 => '1',
		2328 => '0',
		2329 => '1',
		2330 => '0',
		2331 => '1',
		2332 => '0',
		2333 => '1',
		2334 => '0',
		2335 => '1',
		2336 => '0',
		2337 => '1',
		2338 => '0',
		2339 => '1',
		2340 => '0',
		2341 => '1',
		2342 => '0',
		2343 => '1',
		2344 => '0',
		2345 => '1',
		2346 => '0',
		2347 => '1',
		2348 => '0',
		2349 => '1',
		2350 => '0',
		2351 => '1',
		2352 => '0',
		2353 => '1',
		2354 => '0',
		2355 => '1',
		2356 => '0',
		2357 => '1',
		2358 => '0',
		2359 => '1',
		2360 => '0',
		2361 => '1',
		2362 => '0',
		2363 => '1',
		2364 => '0',
		2365 => '1',
		2366 => '0',
		2367 => '1',
		2368 => '0',
		2369 => '1',
		2370 => '0',
		2371 => '1',
		2372 => '0',
		2373 => '1',
		2374 => '0',
		2375 => '1',
		2376 => '0',
		2377 => '1',
		2378 => '0',
		2379 => '1',
		2380 => '0',
		2381 => '1',
		2382 => '0',
		2383 => '1',
		2384 => '0',
		2385 => '1',
		2386 => '0',
		2387 => '1',
		2388 => '0',
		2389 => '1',
		2390 => '0',
		2391 => '1',
		2392 => '0',
		2393 => '1',
		2394 => '0',
		2395 => '1',
		2396 => '0',
		2397 => '1',
		2398 => '0',
		2399 => '1',
		2400 => '0',
		2401 => '1',
		2402 => '0',
		2403 => '1',
		2404 => '0',
		2405 => '1',
		2406 => '0',
		2407 => '1',
		2408 => '0',
		2409 => '1',
		2410 => '0',
		2411 => '1',
		2412 => '0',
		2413 => '1',
		2414 => '0',
		2415 => '1',
		2416 => '0',
		2417 => '1',
		2418 => '0',
		2419 => '1',
		2420 => '0',
		2421 => '1',
		2422 => '0',
		2423 => '1',
		2432 => '1',
		2433 => '0',
		2434 => '1',
		2435 => '0',
		2436 => '1',
		2437 => '0',
		2438 => '1',
		2439 => '0',
		2440 => '1',
		2441 => '0',
		2442 => '1',
		2443 => '0',
		2444 => '1',
		2445 => '0',
		2446 => '1',
		2447 => '0',
		2448 => '1',
		2449 => '0',
		2450 => '1',
		2451 => '0',
		2452 => '1',
		2453 => '0',
		2454 => '1',
		2455 => '0',
		2456 => '1',
		2457 => '0',
		2458 => '1',
		2459 => '0',
		2460 => '1',
		2461 => '0',
		2462 => '1',
		2463 => '0',
		2464 => '1',
		2465 => '0',
		2466 => '1',
		2467 => '0',
		2468 => '1',
		2469 => '0',
		2470 => '1',
		2471 => '0',
		2472 => '1',
		2473 => '0',
		2474 => '1',
		2475 => '0',
		2476 => '1',
		2477 => '0',
		2478 => '1',
		2479 => '0',
		2480 => '1',
		2481 => '0',
		2482 => '1',
		2483 => '0',
		2484 => '1',
		2485 => '0',
		2486 => '1',
		2487 => '0',
		2488 => '1',
		2489 => '0',
		2490 => '1',
		2491 => '0',
		2492 => '1',
		2493 => '0',
		2494 => '1',
		2495 => '0',
		2496 => '1',
		2497 => '0',
		2498 => '1',
		2499 => '0',
		2500 => '1',
		2501 => '0',
		2502 => '1',
		2503 => '0',
		2504 => '1',
		2505 => '0',
		2506 => '1',
		2507 => '0',
		2508 => '1',
		2509 => '0',
		2510 => '1',
		2511 => '0',
		2512 => '1',
		2513 => '0',
		2514 => '1',
		2515 => '0',
		2516 => '1',
		2517 => '0',
		2518 => '1',
		2519 => '0',
		2520 => '1',
		2521 => '0',
		2522 => '1',
		2523 => '0',
		2524 => '1',
		2525 => '0',
		2526 => '1',
		2527 => '0',
		2528 => '1',
		2529 => '0',
		2530 => '1',
		2531 => '0',
		2532 => '1',
		2533 => '0',
		2534 => '1',
		2535 => '0',
		2536 => '1',
		2537 => '0',
		2538 => '1',
		2539 => '0',
		2540 => '1',
		2541 => '0',
		2542 => '1',
		2543 => '0',
		2544 => '1',
		2545 => '0',
		2546 => '1',
		2547 => '0',
		2548 => '1',
		2549 => '0',
		2550 => '1',
		2551 => '0',
		2560 => '0',
		2561 => '1',
		2562 => '0',
		2563 => '1',
		2564 => '0',
		2565 => '1',
		2566 => '0',
		2567 => '1',
		2568 => '0',
		2569 => '1',
		2570 => '0',
		2571 => '1',
		2572 => '0',
		2573 => '1',
		2574 => '0',
		2575 => '1',
		2576 => '0',
		2577 => '1',
		2578 => '0',
		2579 => '1',
		2580 => '0',
		2581 => '1',
		2582 => '0',
		2583 => '1',
		2584 => '0',
		2585 => '1',
		2586 => '0',
		2587 => '1',
		2588 => '0',
		2589 => '1',
		2590 => '0',
		2591 => '1',
		2592 => '0',
		2593 => '1',
		2594 => '0',
		2595 => '1',
		2596 => '0',
		2597 => '1',
		2598 => '0',
		2599 => '1',
		2600 => '0',
		2601 => '1',
		2602 => '0',
		2603 => '1',
		2604 => '0',
		2605 => '1',
		2606 => '0',
		2607 => '1',
		2608 => '0',
		2609 => '1',
		2610 => '0',
		2611 => '1',
		2612 => '0',
		2613 => '1',
		2614 => '0',
		2615 => '1',
		2616 => '0',
		2617 => '1',
		2618 => '0',
		2619 => '1',
		2620 => '0',
		2621 => '1',
		2622 => '0',
		2623 => '1',
		2624 => '0',
		2625 => '1',
		2626 => '0',
		2627 => '1',
		2628 => '0',
		2629 => '1',
		2630 => '0',
		2631 => '1',
		2632 => '0',
		2633 => '1',
		2634 => '0',
		2635 => '1',
		2636 => '0',
		2637 => '1',
		2638 => '0',
		2639 => '1',
		2640 => '0',
		2641 => '1',
		2642 => '0',
		2643 => '1',
		2644 => '0',
		2645 => '1',
		2646 => '0',
		2647 => '1',
		2648 => '0',
		2649 => '1',
		2650 => '0',
		2651 => '1',
		2652 => '0',
		2653 => '1',
		2654 => '0',
		2655 => '1',
		2656 => '0',
		2657 => '1',
		2658 => '0',
		2659 => '1',
		2660 => '0',
		2661 => '1',
		2662 => '0',
		2663 => '1',
		2664 => '0',
		2665 => '1',
		2666 => '0',
		2667 => '1',
		2668 => '0',
		2669 => '1',
		2670 => '0',
		2671 => '1',
		2672 => '0',
		2673 => '1',
		2674 => '0',
		2675 => '1',
		2676 => '0',
		2677 => '1',
		2678 => '0',
		2679 => '1',
		2688 => '1',
		2689 => '0',
		2690 => '1',
		2691 => '0',
		2692 => '1',
		2693 => '0',
		2694 => '1',
		2695 => '0',
		2696 => '1',
		2697 => '0',
		2698 => '1',
		2699 => '0',
		2700 => '1',
		2701 => '0',
		2702 => '1',
		2703 => '0',
		2704 => '1',
		2705 => '0',
		2706 => '1',
		2707 => '0',
		2708 => '1',
		2709 => '0',
		2710 => '1',
		2711 => '0',
		2712 => '1',
		2713 => '0',
		2714 => '1',
		2715 => '0',
		2716 => '1',
		2717 => '0',
		2718 => '1',
		2719 => '0',
		2720 => '1',
		2721 => '0',
		2722 => '1',
		2723 => '0',
		2724 => '1',
		2725 => '0',
		2726 => '1',
		2727 => '0',
		2728 => '1',
		2729 => '0',
		2730 => '1',
		2731 => '0',
		2732 => '1',
		2733 => '0',
		2734 => '1',
		2735 => '0',
		2736 => '1',
		2737 => '0',
		2738 => '1',
		2739 => '0',
		2740 => '1',
		2741 => '0',
		2742 => '1',
		2743 => '0',
		2744 => '1',
		2745 => '0',
		2746 => '1',
		2747 => '0',
		2748 => '1',
		2749 => '0',
		2750 => '1',
		2751 => '0',
		2752 => '1',
		2753 => '0',
		2754 => '1',
		2755 => '0',
		2756 => '1',
		2757 => '0',
		2758 => '1',
		2759 => '0',
		2760 => '1',
		2761 => '0',
		2762 => '1',
		2763 => '0',
		2764 => '1',
		2765 => '0',
		2766 => '1',
		2767 => '0',
		2768 => '1',
		2769 => '0',
		2770 => '1',
		2771 => '0',
		2772 => '1',
		2773 => '0',
		2774 => '1',
		2775 => '0',
		2776 => '1',
		2777 => '0',
		2778 => '1',
		2779 => '0',
		2780 => '1',
		2781 => '0',
		2782 => '1',
		2783 => '0',
		2784 => '1',
		2785 => '0',
		2786 => '1',
		2787 => '0',
		2788 => '1',
		2789 => '0',
		2790 => '1',
		2791 => '0',
		2792 => '1',
		2793 => '0',
		2794 => '1',
		2795 => '0',
		2796 => '1',
		2797 => '0',
		2798 => '1',
		2799 => '0',
		2800 => '1',
		2801 => '0',
		2802 => '1',
		2803 => '0',
		2804 => '1',
		2805 => '0',
		2806 => '1',
		2807 => '0',
		2816 => '0',
		2817 => '1',
		2818 => '0',
		2819 => '1',
		2820 => '0',
		2821 => '1',
		2822 => '0',
		2823 => '1',
		2824 => '0',
		2825 => '1',
		2826 => '0',
		2827 => '1',
		2828 => '0',
		2829 => '1',
		2830 => '0',
		2831 => '1',
		2832 => '0',
		2833 => '1',
		2834 => '0',
		2835 => '1',
		2836 => '0',
		2837 => '1',
		2838 => '0',
		2839 => '1',
		2840 => '0',
		2841 => '1',
		2842 => '0',
		2843 => '1',
		2844 => '0',
		2845 => '1',
		2846 => '0',
		2847 => '1',
		2848 => '0',
		2849 => '1',
		2850 => '0',
		2851 => '1',
		2852 => '0',
		2853 => '1',
		2854 => '0',
		2855 => '1',
		2856 => '0',
		2857 => '1',
		2858 => '0',
		2859 => '1',
		2860 => '0',
		2861 => '1',
		2862 => '0',
		2863 => '1',
		2864 => '0',
		2865 => '1',
		2866 => '0',
		2867 => '1',
		2868 => '0',
		2869 => '1',
		2870 => '0',
		2871 => '1',
		2872 => '0',
		2873 => '1',
		2874 => '0',
		2875 => '1',
		2876 => '0',
		2877 => '1',
		2878 => '0',
		2879 => '1',
		2880 => '0',
		2881 => '1',
		2882 => '0',
		2883 => '1',
		2884 => '0',
		2885 => '1',
		2886 => '0',
		2887 => '1',
		2888 => '0',
		2889 => '1',
		2890 => '0',
		2891 => '1',
		2892 => '0',
		2893 => '1',
		2894 => '0',
		2895 => '1',
		2896 => '0',
		2897 => '1',
		2898 => '0',
		2899 => '1',
		2900 => '0',
		2901 => '1',
		2902 => '0',
		2903 => '1',
		2904 => '0',
		2905 => '1',
		2906 => '0',
		2907 => '1',
		2908 => '0',
		2909 => '1',
		2910 => '0',
		2911 => '1',
		2912 => '0',
		2913 => '1',
		2914 => '0',
		2915 => '1',
		2916 => '0',
		2917 => '1',
		2918 => '0',
		2919 => '1',
		2920 => '0',
		2921 => '1',
		2922 => '0',
		2923 => '1',
		2924 => '0',
		2925 => '1',
		2926 => '0',
		2927 => '1',
		2928 => '0',
		2929 => '1',
		2930 => '0',
		2931 => '1',
		2932 => '0',
		2933 => '1',
		2934 => '0',
		2935 => '1',
		2944 => '1',
		2945 => '0',
		2946 => '1',
		2947 => '0',
		2948 => '1',
		2949 => '0',
		2950 => '1',
		2951 => '0',
		2952 => '1',
		2953 => '0',
		2954 => '1',
		2955 => '0',
		2956 => '1',
		2957 => '0',
		2958 => '1',
		2959 => '0',
		2960 => '1',
		2961 => '0',
		2962 => '1',
		2963 => '0',
		2964 => '1',
		2965 => '0',
		2966 => '1',
		2967 => '0',
		2968 => '1',
		2969 => '0',
		2970 => '1',
		2971 => '0',
		2972 => '1',
		2973 => '0',
		2974 => '1',
		2975 => '0',
		2976 => '1',
		2977 => '0',
		2978 => '1',
		2979 => '0',
		2980 => '1',
		2981 => '0',
		2982 => '1',
		2983 => '0',
		2984 => '1',
		2985 => '0',
		2986 => '1',
		2987 => '0',
		2988 => '1',
		2989 => '0',
		2990 => '1',
		2991 => '0',
		2992 => '1',
		2993 => '0',
		2994 => '1',
		2995 => '0',
		2996 => '1',
		2997 => '0',
		2998 => '1',
		2999 => '0',
		3000 => '1',
		3001 => '0',
		3002 => '1',
		3003 => '0',
		3004 => '1',
		3005 => '0',
		3006 => '1',
		3007 => '0',
		3008 => '1',
		3009 => '0',
		3010 => '1',
		3011 => '0',
		3012 => '1',
		3013 => '0',
		3014 => '1',
		3015 => '0',
		3016 => '1',
		3017 => '0',
		3018 => '1',
		3019 => '0',
		3020 => '1',
		3021 => '0',
		3022 => '1',
		3023 => '0',
		3024 => '1',
		3025 => '0',
		3026 => '1',
		3027 => '0',
		3028 => '1',
		3029 => '0',
		3030 => '1',
		3031 => '0',
		3032 => '1',
		3033 => '0',
		3034 => '1',
		3035 => '0',
		3036 => '1',
		3037 => '0',
		3038 => '1',
		3039 => '0',
		3040 => '1',
		3041 => '0',
		3042 => '1',
		3043 => '0',
		3044 => '1',
		3045 => '0',
		3046 => '1',
		3047 => '0',
		3048 => '1',
		3049 => '0',
		3050 => '1',
		3051 => '0',
		3052 => '1',
		3053 => '0',
		3054 => '1',
		3055 => '0',
		3056 => '1',
		3057 => '0',
		3058 => '1',
		3059 => '0',
		3060 => '1',
		3061 => '0',
		3062 => '1',
		3063 => '0',
		3072 => '0',
		3073 => '1',
		3074 => '0',
		3075 => '1',
		3076 => '0',
		3077 => '1',
		3078 => '0',
		3079 => '1',
		3080 => '0',
		3081 => '1',
		3082 => '0',
		3083 => '1',
		3084 => '0',
		3085 => '1',
		3086 => '0',
		3087 => '1',
		3088 => '0',
		3089 => '1',
		3090 => '0',
		3091 => '1',
		3092 => '0',
		3093 => '1',
		3094 => '0',
		3095 => '1',
		3096 => '0',
		3097 => '1',
		3098 => '0',
		3099 => '1',
		3100 => '0',
		3101 => '1',
		3102 => '0',
		3103 => '1',
		3104 => '0',
		3105 => '1',
		3106 => '0',
		3107 => '1',
		3108 => '0',
		3109 => '1',
		3110 => '0',
		3111 => '1',
		3112 => '0',
		3113 => '1',
		3114 => '0',
		3115 => '1',
		3116 => '0',
		3117 => '1',
		3118 => '0',
		3119 => '1',
		3120 => '0',
		3121 => '1',
		3122 => '0',
		3123 => '1',
		3124 => '0',
		3125 => '1',
		3126 => '0',
		3127 => '1',
		3128 => '0',
		3129 => '1',
		3130 => '0',
		3131 => '1',
		3132 => '0',
		3133 => '1',
		3134 => '0',
		3135 => '1',
		3136 => '0',
		3137 => '1',
		3138 => '0',
		3139 => '1',
		3140 => '0',
		3141 => '1',
		3142 => '0',
		3143 => '1',
		3144 => '0',
		3145 => '1',
		3146 => '0',
		3147 => '1',
		3148 => '0',
		3149 => '1',
		3150 => '0',
		3151 => '1',
		3152 => '0',
		3153 => '1',
		3154 => '0',
		3155 => '1',
		3156 => '0',
		3157 => '1',
		3158 => '0',
		3159 => '1',
		3160 => '0',
		3161 => '1',
		3162 => '0',
		3163 => '1',
		3164 => '0',
		3165 => '1',
		3166 => '0',
		3167 => '1',
		3168 => '0',
		3169 => '1',
		3170 => '0',
		3171 => '1',
		3172 => '0',
		3173 => '1',
		3174 => '0',
		3175 => '1',
		3176 => '0',
		3177 => '1',
		3178 => '0',
		3179 => '1',
		3180 => '0',
		3181 => '1',
		3182 => '0',
		3183 => '1',
		3184 => '0',
		3185 => '1',
		3186 => '0',
		3187 => '1',
		3188 => '0',
		3189 => '1',
		3190 => '0',
		3191 => '1',
		3200 => '1',
		3201 => '0',
		3202 => '1',
		3203 => '0',
		3204 => '1',
		3205 => '0',
		3206 => '1',
		3207 => '0',
		3208 => '1',
		3209 => '0',
		3210 => '1',
		3211 => '0',
		3212 => '1',
		3213 => '0',
		3214 => '1',
		3215 => '0',
		3216 => '1',
		3217 => '0',
		3218 => '1',
		3219 => '0',
		3220 => '1',
		3221 => '0',
		3222 => '1',
		3223 => '0',
		3224 => '1',
		3225 => '0',
		3226 => '1',
		3227 => '0',
		3228 => '1',
		3229 => '0',
		3230 => '1',
		3231 => '0',
		3232 => '1',
		3233 => '0',
		3234 => '1',
		3235 => '0',
		3236 => '1',
		3237 => '0',
		3238 => '1',
		3239 => '0',
		3240 => '1',
		3241 => '0',
		3242 => '1',
		3243 => '0',
		3244 => '1',
		3245 => '0',
		3246 => '1',
		3247 => '0',
		3248 => '1',
		3249 => '0',
		3250 => '1',
		3251 => '0',
		3252 => '1',
		3253 => '0',
		3254 => '1',
		3255 => '0',
		3256 => '1',
		3257 => '0',
		3258 => '1',
		3259 => '0',
		3260 => '1',
		3261 => '0',
		3262 => '1',
		3263 => '0',
		3264 => '1',
		3265 => '0',
		3266 => '1',
		3267 => '0',
		3268 => '1',
		3269 => '0',
		3270 => '1',
		3271 => '0',
		3272 => '1',
		3273 => '0',
		3274 => '1',
		3275 => '0',
		3276 => '1',
		3277 => '0',
		3278 => '1',
		3279 => '0',
		3280 => '1',
		3281 => '0',
		3282 => '1',
		3283 => '0',
		3284 => '1',
		3285 => '0',
		3286 => '1',
		3287 => '0',
		3288 => '1',
		3289 => '0',
		3290 => '1',
		3291 => '0',
		3292 => '1',
		3293 => '0',
		3294 => '1',
		3295 => '0',
		3296 => '1',
		3297 => '0',
		3298 => '1',
		3299 => '0',
		3300 => '1',
		3301 => '0',
		3302 => '1',
		3303 => '0',
		3304 => '1',
		3305 => '0',
		3306 => '1',
		3307 => '0',
		3308 => '1',
		3309 => '0',
		3310 => '1',
		3311 => '0',
		3312 => '1',
		3313 => '0',
		3314 => '1',
		3315 => '0',
		3316 => '1',
		3317 => '0',
		3318 => '1',
		3319 => '0',
		3328 => '0',
		3329 => '1',
		3330 => '0',
		3331 => '1',
		3332 => '0',
		3333 => '1',
		3334 => '0',
		3335 => '1',
		3336 => '0',
		3337 => '1',
		3338 => '0',
		3339 => '1',
		3340 => '0',
		3341 => '1',
		3342 => '0',
		3343 => '1',
		3344 => '0',
		3345 => '1',
		3346 => '0',
		3347 => '1',
		3348 => '0',
		3349 => '1',
		3350 => '0',
		3351 => '1',
		3352 => '0',
		3353 => '1',
		3354 => '0',
		3355 => '1',
		3356 => '0',
		3357 => '1',
		3358 => '0',
		3359 => '1',
		3360 => '0',
		3361 => '1',
		3362 => '0',
		3363 => '1',
		3364 => '0',
		3365 => '1',
		3366 => '0',
		3367 => '1',
		3368 => '0',
		3369 => '1',
		3370 => '0',
		3371 => '1',
		3372 => '0',
		3373 => '1',
		3374 => '0',
		3375 => '1',
		3376 => '0',
		3377 => '1',
		3378 => '0',
		3379 => '1',
		3380 => '0',
		3381 => '1',
		3382 => '0',
		3383 => '1',
		3384 => '0',
		3385 => '1',
		3386 => '0',
		3387 => '1',
		3388 => '0',
		3389 => '1',
		3390 => '0',
		3391 => '1',
		3392 => '0',
		3393 => '1',
		3394 => '0',
		3395 => '1',
		3396 => '0',
		3397 => '1',
		3398 => '0',
		3399 => '1',
		3400 => '0',
		3401 => '1',
		3402 => '0',
		3403 => '1',
		3404 => '0',
		3405 => '1',
		3406 => '0',
		3407 => '1',
		3408 => '0',
		3409 => '1',
		3410 => '0',
		3411 => '1',
		3412 => '0',
		3413 => '1',
		3414 => '0',
		3415 => '1',
		3416 => '0',
		3417 => '1',
		3418 => '0',
		3419 => '1',
		3420 => '0',
		3421 => '1',
		3422 => '0',
		3423 => '1',
		3424 => '0',
		3425 => '1',
		3426 => '0',
		3427 => '1',
		3428 => '0',
		3429 => '1',
		3430 => '0',
		3431 => '1',
		3432 => '0',
		3433 => '1',
		3434 => '0',
		3435 => '1',
		3436 => '0',
		3437 => '1',
		3438 => '0',
		3439 => '1',
		3440 => '0',
		3441 => '1',
		3442 => '0',
		3443 => '1',
		3444 => '0',
		3445 => '1',
		3446 => '0',
		3447 => '1',
		3456 => '1',
		3457 => '0',
		3458 => '1',
		3459 => '0',
		3460 => '1',
		3461 => '0',
		3462 => '1',
		3463 => '0',
		3464 => '1',
		3465 => '0',
		3466 => '1',
		3467 => '0',
		3468 => '1',
		3469 => '0',
		3470 => '1',
		3471 => '0',
		3472 => '1',
		3473 => '0',
		3474 => '1',
		3475 => '0',
		3476 => '1',
		3477 => '0',
		3478 => '1',
		3479 => '0',
		3480 => '1',
		3481 => '0',
		3482 => '1',
		3483 => '0',
		3484 => '1',
		3485 => '0',
		3486 => '1',
		3487 => '0',
		3488 => '1',
		3489 => '0',
		3490 => '1',
		3491 => '0',
		3492 => '1',
		3493 => '0',
		3494 => '1',
		3495 => '0',
		3496 => '1',
		3497 => '0',
		3498 => '1',
		3499 => '0',
		3500 => '1',
		3501 => '0',
		3502 => '1',
		3503 => '0',
		3504 => '1',
		3505 => '0',
		3506 => '1',
		3507 => '0',
		3508 => '1',
		3509 => '0',
		3510 => '1',
		3511 => '0',
		3512 => '1',
		3513 => '0',
		3514 => '1',
		3515 => '0',
		3516 => '1',
		3517 => '0',
		3518 => '1',
		3519 => '0',
		3520 => '1',
		3521 => '0',
		3522 => '1',
		3523 => '0',
		3524 => '1',
		3525 => '0',
		3526 => '1',
		3527 => '0',
		3528 => '1',
		3529 => '0',
		3530 => '1',
		3531 => '0',
		3532 => '1',
		3533 => '0',
		3534 => '1',
		3535 => '0',
		3536 => '1',
		3537 => '0',
		3538 => '1',
		3539 => '0',
		3540 => '1',
		3541 => '0',
		3542 => '1',
		3543 => '0',
		3544 => '1',
		3545 => '0',
		3546 => '1',
		3547 => '0',
		3548 => '1',
		3549 => '0',
		3550 => '1',
		3551 => '0',
		3552 => '1',
		3553 => '0',
		3554 => '1',
		3555 => '0',
		3556 => '1',
		3557 => '0',
		3558 => '1',
		3559 => '0',
		3560 => '1',
		3561 => '0',
		3562 => '1',
		3563 => '0',
		3564 => '1',
		3565 => '0',
		3566 => '1',
		3567 => '0',
		3568 => '1',
		3569 => '0',
		3570 => '1',
		3571 => '0',
		3572 => '1',
		3573 => '0',
		3574 => '1',
		3575 => '0',
		3584 => '0',
		3585 => '1',
		3586 => '0',
		3587 => '1',
		3588 => '0',
		3589 => '1',
		3590 => '0',
		3591 => '1',
		3592 => '0',
		3593 => '1',
		3594 => '0',
		3595 => '1',
		3596 => '0',
		3597 => '1',
		3598 => '0',
		3599 => '1',
		3600 => '0',
		3601 => '1',
		3602 => '0',
		3603 => '1',
		3604 => '0',
		3605 => '1',
		3606 => '0',
		3607 => '1',
		3608 => '0',
		3609 => '1',
		3610 => '0',
		3611 => '1',
		3612 => '0',
		3613 => '1',
		3614 => '0',
		3615 => '1',
		3616 => '0',
		3617 => '1',
		3618 => '0',
		3619 => '1',
		3620 => '0',
		3621 => '1',
		3622 => '0',
		3623 => '1',
		3624 => '0',
		3625 => '1',
		3626 => '0',
		3627 => '1',
		3628 => '0',
		3629 => '1',
		3630 => '0',
		3631 => '1',
		3632 => '0',
		3633 => '1',
		3634 => '0',
		3635 => '1',
		3636 => '0',
		3637 => '1',
		3638 => '0',
		3639 => '1',
		3640 => '0',
		3641 => '1',
		3642 => '0',
		3643 => '1',
		3644 => '0',
		3645 => '1',
		3646 => '0',
		3647 => '1',
		3648 => '0',
		3649 => '1',
		3650 => '0',
		3651 => '1',
		3652 => '0',
		3653 => '1',
		3654 => '0',
		3655 => '1',
		3656 => '0',
		3657 => '1',
		3658 => '0',
		3659 => '1',
		3660 => '0',
		3661 => '1',
		3662 => '0',
		3663 => '1',
		3664 => '0',
		3665 => '1',
		3666 => '0',
		3667 => '1',
		3668 => '0',
		3669 => '1',
		3670 => '0',
		3671 => '1',
		3672 => '0',
		3673 => '1',
		3674 => '0',
		3675 => '1',
		3676 => '0',
		3677 => '1',
		3678 => '0',
		3679 => '1',
		3680 => '0',
		3681 => '1',
		3682 => '0',
		3683 => '1',
		3684 => '0',
		3685 => '1',
		3686 => '0',
		3687 => '1',
		3688 => '0',
		3689 => '1',
		3690 => '0',
		3691 => '1',
		3692 => '0',
		3693 => '1',
		3694 => '0',
		3695 => '1',
		3696 => '0',
		3697 => '1',
		3698 => '0',
		3699 => '1',
		3700 => '0',
		3701 => '1',
		3702 => '0',
		3703 => '1',
		3712 => '1',
		3713 => '0',
		3714 => '1',
		3715 => '0',
		3716 => '1',
		3717 => '0',
		3718 => '1',
		3719 => '0',
		3720 => '1',
		3721 => '0',
		3722 => '1',
		3723 => '0',
		3724 => '1',
		3725 => '0',
		3726 => '1',
		3727 => '0',
		3728 => '1',
		3729 => '0',
		3730 => '1',
		3731 => '0',
		3732 => '1',
		3733 => '0',
		3734 => '1',
		3735 => '0',
		3736 => '1',
		3737 => '0',
		3738 => '1',
		3739 => '0',
		3740 => '1',
		3741 => '0',
		3742 => '1',
		3743 => '0',
		3744 => '1',
		3745 => '0',
		3746 => '1',
		3747 => '0',
		3748 => '1',
		3749 => '0',
		3750 => '1',
		3751 => '0',
		3752 => '1',
		3753 => '0',
		3754 => '1',
		3755 => '0',
		3756 => '1',
		3757 => '0',
		3758 => '1',
		3759 => '0',
		3760 => '1',
		3761 => '0',
		3762 => '1',
		3763 => '0',
		3764 => '1',
		3765 => '0',
		3766 => '1',
		3767 => '0',
		3768 => '1',
		3769 => '0',
		3770 => '1',
		3771 => '0',
		3772 => '1',
		3773 => '0',
		3774 => '1',
		3775 => '0',
		3776 => '1',
		3777 => '0',
		3778 => '1',
		3779 => '0',
		3780 => '1',
		3781 => '0',
		3782 => '1',
		3783 => '0',
		3784 => '1',
		3785 => '0',
		3786 => '1',
		3787 => '0',
		3788 => '1',
		3789 => '0',
		3790 => '1',
		3791 => '0',
		3792 => '1',
		3793 => '0',
		3794 => '1',
		3795 => '0',
		3796 => '1',
		3797 => '0',
		3798 => '1',
		3799 => '0',
		3800 => '1',
		3801 => '0',
		3802 => '1',
		3803 => '0',
		3804 => '1',
		3805 => '0',
		3806 => '1',
		3807 => '0',
		3808 => '1',
		3809 => '0',
		3810 => '1',
		3811 => '0',
		3812 => '1',
		3813 => '0',
		3814 => '1',
		3815 => '0',
		3816 => '1',
		3817 => '0',
		3818 => '1',
		3819 => '0',
		3820 => '1',
		3821 => '0',
		3822 => '1',
		3823 => '0',
		3824 => '1',
		3825 => '0',
		3826 => '1',
		3827 => '0',
		3828 => '1',
		3829 => '0',
		3830 => '1',
		3831 => '0',
		3840 => '0',
		3841 => '1',
		3842 => '0',
		3843 => '1',
		3844 => '0',
		3845 => '1',
		3846 => '0',
		3847 => '1',
		3848 => '0',
		3849 => '1',
		3850 => '0',
		3851 => '1',
		3852 => '0',
		3853 => '1',
		3854 => '0',
		3855 => '1',
		3856 => '0',
		3857 => '1',
		3858 => '0',
		3859 => '1',
		3860 => '0',
		3861 => '1',
		3862 => '0',
		3863 => '1',
		3864 => '0',
		3865 => '1',
		3866 => '0',
		3867 => '1',
		3868 => '0',
		3869 => '1',
		3870 => '0',
		3871 => '1',
		3872 => '0',
		3873 => '1',
		3874 => '0',
		3875 => '1',
		3876 => '0',
		3877 => '1',
		3878 => '0',
		3879 => '1',
		3880 => '0',
		3881 => '1',
		3882 => '0',
		3883 => '1',
		3884 => '0',
		3885 => '1',
		3886 => '0',
		3887 => '1',
		3888 => '0',
		3889 => '1',
		3890 => '0',
		3891 => '1',
		3892 => '0',
		3893 => '1',
		3894 => '0',
		3895 => '1',
		3896 => '0',
		3897 => '1',
		3898 => '0',
		3899 => '1',
		3900 => '0',
		3901 => '1',
		3902 => '0',
		3903 => '1',
		3904 => '0',
		3905 => '1',
		3906 => '0',
		3907 => '1',
		3908 => '0',
		3909 => '1',
		3910 => '0',
		3911 => '1',
		3912 => '0',
		3913 => '1',
		3914 => '0',
		3915 => '1',
		3916 => '0',
		3917 => '1',
		3918 => '0',
		3919 => '1',
		3920 => '0',
		3921 => '1',
		3922 => '0',
		3923 => '1',
		3924 => '0',
		3925 => '1',
		3926 => '0',
		3927 => '1',
		3928 => '0',
		3929 => '1',
		3930 => '0',
		3931 => '1',
		3932 => '0',
		3933 => '1',
		3934 => '0',
		3935 => '1',
		3936 => '0',
		3937 => '1',
		3938 => '0',
		3939 => '1',
		3940 => '0',
		3941 => '1',
		3942 => '0',
		3943 => '1',
		3944 => '0',
		3945 => '1',
		3946 => '0',
		3947 => '1',
		3948 => '0',
		3949 => '1',
		3950 => '0',
		3951 => '1',
		3952 => '0',
		3953 => '1',
		3954 => '0',
		3955 => '1',
		3956 => '0',
		3957 => '1',
		3958 => '0',
		3959 => '1',
		3968 => '1',
		3969 => '0',
		3970 => '1',
		3971 => '0',
		3972 => '1',
		3973 => '0',
		3974 => '1',
		3975 => '0',
		3976 => '1',
		3977 => '0',
		3978 => '1',
		3979 => '0',
		3980 => '1',
		3981 => '0',
		3982 => '1',
		3983 => '0',
		3984 => '1',
		3985 => '0',
		3986 => '1',
		3987 => '0',
		3988 => '1',
		3989 => '0',
		3990 => '1',
		3991 => '0',
		3992 => '1',
		3993 => '0',
		3994 => '1',
		3995 => '0',
		3996 => '1',
		3997 => '0',
		3998 => '1',
		3999 => '0',
		4000 => '1',
		4001 => '0',
		4002 => '1',
		4003 => '0',
		4004 => '1',
		4005 => '0',
		4006 => '1',
		4007 => '0',
		4008 => '1',
		4009 => '0',
		4010 => '1',
		4011 => '0',
		4012 => '1',
		4013 => '0',
		4014 => '1',
		4015 => '0',
		4016 => '1',
		4017 => '0',
		4018 => '1',
		4019 => '0',
		4020 => '1',
		4021 => '0',
		4022 => '1',
		4023 => '0',
		4024 => '1',
		4025 => '0',
		4026 => '1',
		4027 => '0',
		4028 => '1',
		4029 => '0',
		4030 => '1',
		4031 => '0',
		4032 => '1',
		4033 => '0',
		4034 => '1',
		4035 => '0',
		4036 => '1',
		4037 => '0',
		4038 => '1',
		4039 => '0',
		4040 => '1',
		4041 => '0',
		4042 => '1',
		4043 => '0',
		4044 => '1',
		4045 => '0',
		4046 => '1',
		4047 => '0',
		4048 => '1',
		4049 => '0',
		4050 => '1',
		4051 => '0',
		4052 => '1',
		4053 => '0',
		4054 => '1',
		4055 => '0',
		4056 => '1',
		4057 => '0',
		4058 => '1',
		4059 => '0',
		4060 => '1',
		4061 => '0',
		4062 => '1',
		4063 => '0',
		4064 => '1',
		4065 => '0',
		4066 => '1',
		4067 => '0',
		4068 => '1',
		4069 => '0',
		4070 => '1',
		4071 => '0',
		4072 => '1',
		4073 => '0',
		4074 => '1',
		4075 => '0',
		4076 => '1',
		4077 => '0',
		4078 => '1',
		4079 => '0',
		4080 => '1',
		4081 => '0',
		4082 => '1',
		4083 => '0',
		4084 => '1',
		4085 => '0',
		4086 => '1',
		4087 => '0',
		4096 => '0',
		4097 => '1',
		4098 => '0',
		4099 => '1',
		4100 => '0',
		4101 => '1',
		4102 => '0',
		4103 => '1',
		4104 => '0',
		4105 => '1',
		4106 => '0',
		4107 => '1',
		4108 => '0',
		4109 => '1',
		4110 => '0',
		4111 => '1',
		4112 => '0',
		4113 => '1',
		4114 => '0',
		4115 => '1',
		4116 => '0',
		4117 => '1',
		4118 => '0',
		4119 => '1',
		4120 => '0',
		4121 => '1',
		4122 => '0',
		4123 => '1',
		4124 => '0',
		4125 => '1',
		4126 => '0',
		4127 => '1',
		4128 => '0',
		4129 => '1',
		4130 => '0',
		4131 => '1',
		4132 => '0',
		4133 => '1',
		4134 => '0',
		4135 => '1',
		4136 => '0',
		4137 => '1',
		4138 => '0',
		4139 => '1',
		4140 => '0',
		4141 => '1',
		4142 => '0',
		4143 => '1',
		4144 => '0',
		4145 => '1',
		4146 => '0',
		4147 => '1',
		4148 => '0',
		4149 => '1',
		4150 => '0',
		4151 => '1',
		4152 => '0',
		4153 => '1',
		4154 => '0',
		4155 => '1',
		4156 => '0',
		4157 => '1',
		4158 => '0',
		4159 => '1',
		4160 => '0',
		4161 => '1',
		4162 => '0',
		4163 => '1',
		4164 => '0',
		4165 => '1',
		4166 => '0',
		4167 => '1',
		4168 => '0',
		4169 => '1',
		4170 => '0',
		4171 => '1',
		4172 => '0',
		4173 => '1',
		4174 => '0',
		4175 => '1',
		4176 => '0',
		4177 => '1',
		4178 => '0',
		4179 => '1',
		4180 => '0',
		4181 => '1',
		4182 => '0',
		4183 => '1',
		4184 => '0',
		4185 => '1',
		4186 => '0',
		4187 => '1',
		4188 => '0',
		4189 => '1',
		4190 => '0',
		4191 => '1',
		4192 => '0',
		4193 => '1',
		4194 => '0',
		4195 => '1',
		4196 => '0',
		4197 => '1',
		4198 => '0',
		4199 => '1',
		4200 => '0',
		4201 => '1',
		4202 => '0',
		4203 => '1',
		4204 => '0',
		4205 => '1',
		4206 => '0',
		4207 => '1',
		4208 => '0',
		4209 => '1',
		4210 => '0',
		4211 => '1',
		4212 => '0',
		4213 => '1',
		4214 => '0',
		4215 => '1',
		4224 => '1',
		4225 => '0',
		4226 => '1',
		4227 => '0',
		4228 => '1',
		4229 => '0',
		4230 => '1',
		4231 => '0',
		4232 => '1',
		4233 => '0',
		4234 => '1',
		4235 => '0',
		4236 => '1',
		4237 => '0',
		4238 => '1',
		4239 => '0',
		4240 => '1',
		4241 => '0',
		4242 => '1',
		4243 => '0',
		4244 => '1',
		4245 => '0',
		4246 => '1',
		4247 => '0',
		4248 => '1',
		4249 => '0',
		4250 => '1',
		4251 => '0',
		4252 => '1',
		4253 => '0',
		4254 => '1',
		4255 => '0',
		4256 => '1',
		4257 => '0',
		4258 => '1',
		4259 => '0',
		4260 => '1',
		4261 => '0',
		4262 => '1',
		4263 => '0',
		4264 => '1',
		4265 => '0',
		4266 => '1',
		4267 => '0',
		4268 => '1',
		4269 => '0',
		4270 => '1',
		4271 => '0',
		4272 => '1',
		4273 => '0',
		4274 => '1',
		4275 => '0',
		4276 => '1',
		4277 => '0',
		4278 => '1',
		4279 => '0',
		4280 => '1',
		4281 => '0',
		4282 => '1',
		4283 => '0',
		4284 => '1',
		4285 => '0',
		4286 => '1',
		4287 => '0',
		4288 => '1',
		4289 => '0',
		4290 => '1',
		4291 => '0',
		4292 => '1',
		4293 => '0',
		4294 => '1',
		4295 => '0',
		4296 => '1',
		4297 => '0',
		4298 => '1',
		4299 => '0',
		4300 => '1',
		4301 => '0',
		4302 => '1',
		4303 => '0',
		4304 => '1',
		4305 => '0',
		4306 => '1',
		4307 => '0',
		4308 => '1',
		4309 => '0',
		4310 => '1',
		4311 => '0',
		4312 => '1',
		4313 => '0',
		4314 => '1',
		4315 => '0',
		4316 => '1',
		4317 => '0',
		4318 => '1',
		4319 => '0',
		4320 => '1',
		4321 => '0',
		4322 => '1',
		4323 => '0',
		4324 => '1',
		4325 => '0',
		4326 => '1',
		4327 => '0',
		4328 => '1',
		4329 => '0',
		4330 => '1',
		4331 => '0',
		4332 => '1',
		4333 => '0',
		4334 => '1',
		4335 => '0',
		4336 => '1',
		4337 => '0',
		4338 => '1',
		4339 => '0',
		4340 => '1',
		4341 => '0',
		4342 => '1',
		4343 => '0',
		4352 => '0',
		4353 => '1',
		4354 => '0',
		4355 => '1',
		4356 => '0',
		4357 => '1',
		4358 => '0',
		4359 => '1',
		4360 => '0',
		4361 => '1',
		4362 => '0',
		4363 => '1',
		4364 => '0',
		4365 => '1',
		4366 => '0',
		4367 => '1',
		4368 => '0',
		4369 => '1',
		4370 => '0',
		4371 => '1',
		4372 => '0',
		4373 => '1',
		4374 => '0',
		4375 => '1',
		4376 => '0',
		4377 => '1',
		4378 => '0',
		4379 => '1',
		4380 => '0',
		4381 => '1',
		4382 => '0',
		4383 => '1',
		4384 => '0',
		4385 => '1',
		4386 => '0',
		4387 => '1',
		4388 => '0',
		4389 => '1',
		4390 => '0',
		4391 => '1',
		4392 => '0',
		4393 => '1',
		4394 => '0',
		4395 => '1',
		4396 => '0',
		4397 => '1',
		4398 => '0',
		4399 => '1',
		4400 => '0',
		4401 => '1',
		4402 => '0',
		4403 => '1',
		4404 => '0',
		4405 => '1',
		4406 => '0',
		4407 => '1',
		4408 => '0',
		4409 => '1',
		4410 => '0',
		4411 => '1',
		4412 => '0',
		4413 => '1',
		4414 => '0',
		4415 => '1',
		4416 => '0',
		4417 => '1',
		4418 => '0',
		4419 => '1',
		4420 => '0',
		4421 => '1',
		4422 => '0',
		4423 => '1',
		4424 => '0',
		4425 => '1',
		4426 => '0',
		4427 => '1',
		4428 => '0',
		4429 => '1',
		4430 => '0',
		4431 => '1',
		4432 => '0',
		4433 => '1',
		4434 => '0',
		4435 => '1',
		4436 => '0',
		4437 => '1',
		4438 => '0',
		4439 => '1',
		4440 => '0',
		4441 => '1',
		4442 => '0',
		4443 => '1',
		4444 => '0',
		4445 => '1',
		4446 => '0',
		4447 => '1',
		4448 => '0',
		4449 => '1',
		4450 => '0',
		4451 => '1',
		4452 => '0',
		4453 => '1',
		4454 => '0',
		4455 => '1',
		4456 => '0',
		4457 => '1',
		4458 => '0',
		4459 => '1',
		4460 => '0',
		4461 => '1',
		4462 => '0',
		4463 => '1',
		4464 => '0',
		4465 => '1',
		4466 => '0',
		4467 => '1',
		4468 => '0',
		4469 => '1',
		4470 => '0',
		4471 => '1',
		4480 => '1',
		4481 => '0',
		4482 => '1',
		4483 => '0',
		4484 => '1',
		4485 => '0',
		4486 => '1',
		4487 => '0',
		4488 => '1',
		4489 => '0',
		4490 => '1',
		4491 => '0',
		4492 => '1',
		4493 => '0',
		4494 => '1',
		4495 => '0',
		4496 => '1',
		4497 => '0',
		4498 => '1',
		4499 => '0',
		4500 => '1',
		4501 => '0',
		4502 => '1',
		4503 => '0',
		4504 => '1',
		4505 => '0',
		4506 => '1',
		4507 => '0',
		4508 => '1',
		4509 => '0',
		4510 => '1',
		4511 => '0',
		4512 => '1',
		4513 => '0',
		4514 => '1',
		4515 => '0',
		4516 => '1',
		4517 => '0',
		4518 => '1',
		4519 => '0',
		4520 => '1',
		4521 => '0',
		4522 => '1',
		4523 => '0',
		4524 => '1',
		4525 => '0',
		4526 => '1',
		4527 => '0',
		4528 => '1',
		4529 => '0',
		4530 => '1',
		4531 => '0',
		4532 => '1',
		4533 => '0',
		4534 => '1',
		4535 => '0',
		4536 => '1',
		4537 => '0',
		4538 => '1',
		4539 => '0',
		4540 => '1',
		4541 => '0',
		4542 => '1',
		4543 => '0',
		4544 => '1',
		4545 => '0',
		4546 => '1',
		4547 => '0',
		4548 => '1',
		4549 => '0',
		4550 => '1',
		4551 => '0',
		4552 => '1',
		4553 => '0',
		4554 => '1',
		4555 => '0',
		4556 => '1',
		4557 => '0',
		4558 => '1',
		4559 => '0',
		4560 => '1',
		4561 => '0',
		4562 => '1',
		4563 => '0',
		4564 => '1',
		4565 => '0',
		4566 => '1',
		4567 => '0',
		4568 => '1',
		4569 => '0',
		4570 => '1',
		4571 => '0',
		4572 => '1',
		4573 => '0',
		4574 => '1',
		4575 => '0',
		4576 => '1',
		4577 => '0',
		4578 => '1',
		4579 => '0',
		4580 => '1',
		4581 => '0',
		4582 => '1',
		4583 => '0',
		4584 => '1',
		4585 => '0',
		4586 => '1',
		4587 => '0',
		4588 => '1',
		4589 => '0',
		4590 => '1',
		4591 => '0',
		4592 => '1',
		4593 => '0',
		4594 => '1',
		4595 => '0',
		4596 => '1',
		4597 => '0',
		4598 => '1',
		4599 => '0',
		4608 => '0',
		4609 => '1',
		4610 => '0',
		4611 => '1',
		4612 => '0',
		4613 => '1',
		4614 => '0',
		4615 => '1',
		4616 => '0',
		4617 => '1',
		4618 => '0',
		4619 => '1',
		4620 => '0',
		4621 => '1',
		4622 => '0',
		4623 => '1',
		4624 => '0',
		4625 => '1',
		4626 => '0',
		4627 => '1',
		4628 => '0',
		4629 => '1',
		4630 => '0',
		4631 => '1',
		4632 => '0',
		4633 => '1',
		4634 => '0',
		4635 => '1',
		4636 => '0',
		4637 => '1',
		4638 => '0',
		4639 => '1',
		4640 => '0',
		4641 => '1',
		4642 => '0',
		4643 => '1',
		4644 => '0',
		4645 => '1',
		4646 => '0',
		4647 => '1',
		4648 => '0',
		4649 => '1',
		4650 => '0',
		4651 => '1',
		4652 => '0',
		4653 => '1',
		4654 => '0',
		4655 => '1',
		4656 => '0',
		4657 => '1',
		4658 => '0',
		4659 => '1',
		4660 => '0',
		4661 => '1',
		4662 => '0',
		4663 => '1',
		4664 => '0',
		4665 => '1',
		4666 => '0',
		4667 => '1',
		4668 => '0',
		4669 => '1',
		4670 => '0',
		4671 => '1',
		4672 => '0',
		4673 => '1',
		4674 => '0',
		4675 => '1',
		4676 => '0',
		4677 => '1',
		4678 => '0',
		4679 => '1',
		4680 => '0',
		4681 => '1',
		4682 => '0',
		4683 => '1',
		4684 => '0',
		4685 => '1',
		4686 => '0',
		4687 => '1',
		4688 => '0',
		4689 => '1',
		4690 => '0',
		4691 => '1',
		4692 => '0',
		4693 => '1',
		4694 => '0',
		4695 => '1',
		4696 => '0',
		4697 => '1',
		4698 => '0',
		4699 => '1',
		4700 => '0',
		4701 => '1',
		4702 => '0',
		4703 => '1',
		4704 => '0',
		4705 => '1',
		4706 => '0',
		4707 => '1',
		4708 => '0',
		4709 => '1',
		4710 => '0',
		4711 => '1',
		4712 => '0',
		4713 => '1',
		4714 => '0',
		4715 => '1',
		4716 => '0',
		4717 => '1',
		4718 => '0',
		4719 => '1',
		4720 => '0',
		4721 => '1',
		4722 => '0',
		4723 => '1',
		4724 => '0',
		4725 => '1',
		4726 => '0',
		4727 => '1',
		4736 => '1',
		4737 => '0',
		4738 => '1',
		4739 => '0',
		4740 => '1',
		4741 => '0',
		4742 => '1',
		4743 => '0',
		4744 => '1',
		4745 => '0',
		4746 => '1',
		4747 => '0',
		4748 => '1',
		4749 => '0',
		4750 => '1',
		4751 => '0',
		4752 => '1',
		4753 => '0',
		4754 => '1',
		4755 => '0',
		4756 => '1',
		4757 => '0',
		4758 => '1',
		4759 => '0',
		4760 => '1',
		4761 => '0',
		4762 => '1',
		4763 => '0',
		4764 => '1',
		4765 => '0',
		4766 => '1',
		4767 => '0',
		4768 => '1',
		4769 => '0',
		4770 => '1',
		4771 => '0',
		4772 => '1',
		4773 => '0',
		4774 => '1',
		4775 => '0',
		4776 => '1',
		4777 => '0',
		4778 => '1',
		4779 => '0',
		4780 => '1',
		4781 => '0',
		4782 => '1',
		4783 => '0',
		4784 => '1',
		4785 => '0',
		4786 => '1',
		4787 => '0',
		4788 => '1',
		4789 => '0',
		4790 => '1',
		4791 => '0',
		4792 => '1',
		4793 => '0',
		4794 => '1',
		4795 => '0',
		4796 => '1',
		4797 => '0',
		4798 => '1',
		4799 => '0',
		4800 => '1',
		4801 => '0',
		4802 => '1',
		4803 => '0',
		4804 => '1',
		4805 => '0',
		4806 => '1',
		4807 => '0',
		4808 => '1',
		4809 => '0',
		4810 => '1',
		4811 => '0',
		4812 => '1',
		4813 => '0',
		4814 => '1',
		4815 => '0',
		4816 => '1',
		4817 => '0',
		4818 => '1',
		4819 => '0',
		4820 => '1',
		4821 => '0',
		4822 => '1',
		4823 => '0',
		4824 => '1',
		4825 => '0',
		4826 => '1',
		4827 => '0',
		4828 => '1',
		4829 => '0',
		4830 => '1',
		4831 => '0',
		4832 => '1',
		4833 => '0',
		4834 => '1',
		4835 => '0',
		4836 => '1',
		4837 => '0',
		4838 => '1',
		4839 => '0',
		4840 => '1',
		4841 => '0',
		4842 => '1',
		4843 => '0',
		4844 => '1',
		4845 => '0',
		4846 => '1',
		4847 => '0',
		4848 => '1',
		4849 => '0',
		4850 => '1',
		4851 => '0',
		4852 => '1',
		4853 => '0',
		4854 => '1',
		4855 => '0',
		4864 => '0',
		4865 => '1',
		4866 => '0',
		4867 => '1',
		4868 => '0',
		4869 => '1',
		4870 => '0',
		4871 => '1',
		4872 => '0',
		4873 => '1',
		4874 => '0',
		4875 => '1',
		4876 => '0',
		4877 => '1',
		4878 => '0',
		4879 => '1',
		4880 => '0',
		4881 => '1',
		4882 => '0',
		4883 => '1',
		4884 => '0',
		4885 => '1',
		4886 => '0',
		4887 => '1',
		4888 => '0',
		4889 => '1',
		4890 => '0',
		4891 => '1',
		4892 => '0',
		4893 => '1',
		4894 => '0',
		4895 => '1',
		4896 => '0',
		4897 => '1',
		4898 => '0',
		4899 => '1',
		4900 => '0',
		4901 => '1',
		4902 => '0',
		4903 => '1',
		4904 => '0',
		4905 => '1',
		4906 => '0',
		4907 => '1',
		4908 => '0',
		4909 => '1',
		4910 => '0',
		4911 => '1',
		4912 => '0',
		4913 => '1',
		4914 => '0',
		4915 => '1',
		4916 => '0',
		4917 => '1',
		4918 => '0',
		4919 => '1',
		4920 => '0',
		4921 => '1',
		4922 => '0',
		4923 => '1',
		4924 => '0',
		4925 => '1',
		4926 => '0',
		4927 => '1',
		4928 => '0',
		4929 => '1',
		4930 => '0',
		4931 => '1',
		4932 => '0',
		4933 => '1',
		4934 => '0',
		4935 => '1',
		4936 => '0',
		4937 => '1',
		4938 => '0',
		4939 => '1',
		4940 => '0',
		4941 => '1',
		4942 => '0',
		4943 => '1',
		4944 => '0',
		4945 => '1',
		4946 => '0',
		4947 => '1',
		4948 => '0',
		4949 => '1',
		4950 => '0',
		4951 => '1',
		4952 => '0',
		4953 => '1',
		4954 => '0',
		4955 => '1',
		4956 => '0',
		4957 => '1',
		4958 => '0',
		4959 => '1',
		4960 => '0',
		4961 => '1',
		4962 => '0',
		4963 => '1',
		4964 => '0',
		4965 => '1',
		4966 => '0',
		4967 => '1',
		4968 => '0',
		4969 => '1',
		4970 => '0',
		4971 => '1',
		4972 => '0',
		4973 => '1',
		4974 => '0',
		4975 => '1',
		4976 => '0',
		4977 => '1',
		4978 => '0',
		4979 => '1',
		4980 => '0',
		4981 => '1',
		4982 => '0',
		4983 => '1',
		4992 => '1',
		4993 => '0',
		4994 => '1',
		4995 => '0',
		4996 => '1',
		4997 => '0',
		4998 => '1',
		4999 => '0',
		5000 => '1',
		5001 => '0',
		5002 => '1',
		5003 => '0',
		5004 => '1',
		5005 => '0',
		5006 => '1',
		5007 => '0',
		5008 => '1',
		5009 => '0',
		5010 => '1',
		5011 => '0',
		5012 => '1',
		5013 => '0',
		5014 => '1',
		5015 => '0',
		5016 => '1',
		5017 => '0',
		5018 => '1',
		5019 => '0',
		5020 => '1',
		5021 => '0',
		5022 => '1',
		5023 => '0',
		5024 => '1',
		5025 => '0',
		5026 => '1',
		5027 => '0',
		5028 => '1',
		5029 => '0',
		5030 => '1',
		5031 => '0',
		5032 => '1',
		5033 => '0',
		5034 => '1',
		5035 => '0',
		5036 => '1',
		5037 => '0',
		5038 => '1',
		5039 => '0',
		5040 => '1',
		5041 => '0',
		5042 => '1',
		5043 => '0',
		5044 => '1',
		5045 => '0',
		5046 => '1',
		5047 => '0',
		5048 => '1',
		5049 => '0',
		5050 => '1',
		5051 => '0',
		5052 => '1',
		5053 => '0',
		5054 => '1',
		5055 => '0',
		5056 => '1',
		5057 => '0',
		5058 => '1',
		5059 => '0',
		5060 => '1',
		5061 => '0',
		5062 => '1',
		5063 => '0',
		5064 => '1',
		5065 => '0',
		5066 => '1',
		5067 => '0',
		5068 => '1',
		5069 => '0',
		5070 => '1',
		5071 => '0',
		5072 => '1',
		5073 => '0',
		5074 => '1',
		5075 => '0',
		5076 => '1',
		5077 => '0',
		5078 => '1',
		5079 => '0',
		5080 => '1',
		5081 => '0',
		5082 => '1',
		5083 => '0',
		5084 => '1',
		5085 => '0',
		5086 => '1',
		5087 => '0',
		5088 => '1',
		5089 => '0',
		5090 => '1',
		5091 => '0',
		5092 => '1',
		5093 => '0',
		5094 => '1',
		5095 => '0',
		5096 => '1',
		5097 => '0',
		5098 => '1',
		5099 => '0',
		5100 => '1',
		5101 => '0',
		5102 => '1',
		5103 => '0',
		5104 => '1',
		5105 => '0',
		5106 => '1',
		5107 => '0',
		5108 => '1',
		5109 => '0',
		5110 => '1',
		5111 => '0',
		5120 => '0',
		5121 => '1',
		5122 => '0',
		5123 => '1',
		5124 => '0',
		5125 => '1',
		5126 => '0',
		5127 => '1',
		5128 => '0',
		5129 => '1',
		5130 => '0',
		5131 => '1',
		5132 => '0',
		5133 => '1',
		5134 => '0',
		5135 => '1',
		5136 => '0',
		5137 => '1',
		5138 => '0',
		5139 => '1',
		5140 => '0',
		5141 => '1',
		5142 => '0',
		5143 => '1',
		5144 => '0',
		5145 => '1',
		5146 => '0',
		5147 => '1',
		5148 => '0',
		5149 => '1',
		5150 => '0',
		5151 => '1',
		5152 => '0',
		5153 => '1',
		5154 => '0',
		5155 => '1',
		5156 => '0',
		5157 => '1',
		5158 => '0',
		5159 => '1',
		5160 => '0',
		5161 => '1',
		5162 => '0',
		5163 => '1',
		5164 => '0',
		5165 => '1',
		5166 => '0',
		5167 => '1',
		5168 => '0',
		5169 => '1',
		5170 => '0',
		5171 => '1',
		5172 => '0',
		5173 => '1',
		5174 => '0',
		5175 => '1',
		5176 => '0',
		5177 => '1',
		5178 => '0',
		5179 => '1',
		5180 => '0',
		5181 => '1',
		5182 => '0',
		5183 => '1',
		5184 => '0',
		5185 => '1',
		5186 => '0',
		5187 => '1',
		5188 => '0',
		5189 => '1',
		5190 => '0',
		5191 => '1',
		5192 => '0',
		5193 => '1',
		5194 => '0',
		5195 => '1',
		5196 => '0',
		5197 => '1',
		5198 => '0',
		5199 => '1',
		5200 => '0',
		5201 => '1',
		5202 => '0',
		5203 => '1',
		5204 => '0',
		5205 => '1',
		5206 => '0',
		5207 => '1',
		5208 => '0',
		5209 => '1',
		5210 => '0',
		5211 => '1',
		5212 => '0',
		5213 => '1',
		5214 => '0',
		5215 => '1',
		5216 => '0',
		5217 => '1',
		5218 => '0',
		5219 => '1',
		5220 => '0',
		5221 => '1',
		5222 => '0',
		5223 => '1',
		5224 => '0',
		5225 => '1',
		5226 => '0',
		5227 => '1',
		5228 => '0',
		5229 => '1',
		5230 => '0',
		5231 => '1',
		5232 => '0',
		5233 => '1',
		5234 => '0',
		5235 => '1',
		5236 => '0',
		5237 => '1',
		5238 => '0',
		5239 => '1',
		5248 => '1',
		5249 => '0',
		5250 => '1',
		5251 => '0',
		5252 => '1',
		5253 => '0',
		5254 => '1',
		5255 => '0',
		5256 => '1',
		5257 => '0',
		5258 => '1',
		5259 => '0',
		5260 => '1',
		5261 => '0',
		5262 => '1',
		5263 => '0',
		5264 => '1',
		5265 => '0',
		5266 => '1',
		5267 => '0',
		5268 => '1',
		5269 => '0',
		5270 => '1',
		5271 => '0',
		5272 => '1',
		5273 => '0',
		5274 => '1',
		5275 => '0',
		5276 => '1',
		5277 => '0',
		5278 => '1',
		5279 => '0',
		5280 => '1',
		5281 => '0',
		5282 => '1',
		5283 => '0',
		5284 => '1',
		5285 => '0',
		5286 => '1',
		5287 => '0',
		5288 => '1',
		5289 => '0',
		5290 => '1',
		5291 => '0',
		5292 => '1',
		5293 => '0',
		5294 => '1',
		5295 => '0',
		5296 => '1',
		5297 => '0',
		5298 => '1',
		5299 => '0',
		5300 => '1',
		5301 => '0',
		5302 => '1',
		5303 => '0',
		5304 => '1',
		5305 => '0',
		5306 => '1',
		5307 => '0',
		5308 => '1',
		5309 => '0',
		5310 => '1',
		5311 => '0',
		5312 => '1',
		5313 => '0',
		5314 => '1',
		5315 => '0',
		5316 => '1',
		5317 => '0',
		5318 => '1',
		5319 => '0',
		5320 => '1',
		5321 => '0',
		5322 => '1',
		5323 => '0',
		5324 => '1',
		5325 => '0',
		5326 => '1',
		5327 => '0',
		5328 => '1',
		5329 => '0',
		5330 => '1',
		5331 => '0',
		5332 => '1',
		5333 => '0',
		5334 => '1',
		5335 => '0',
		5336 => '1',
		5337 => '0',
		5338 => '1',
		5339 => '0',
		5340 => '1',
		5341 => '0',
		5342 => '1',
		5343 => '0',
		5344 => '1',
		5345 => '0',
		5346 => '1',
		5347 => '0',
		5348 => '1',
		5349 => '0',
		5350 => '1',
		5351 => '0',
		5352 => '1',
		5353 => '0',
		5354 => '1',
		5355 => '0',
		5356 => '1',
		5357 => '0',
		5358 => '1',
		5359 => '0',
		5360 => '1',
		5361 => '0',
		5362 => '1',
		5363 => '0',
		5364 => '1',
		5365 => '0',
		5366 => '1',
		5367 => '0',
		5376 => '0',
		5377 => '1',
		5378 => '0',
		5379 => '1',
		5380 => '0',
		5381 => '1',
		5382 => '0',
		5383 => '1',
		5384 => '0',
		5385 => '1',
		5386 => '0',
		5387 => '1',
		5388 => '0',
		5389 => '1',
		5390 => '0',
		5391 => '1',
		5392 => '0',
		5393 => '1',
		5394 => '0',
		5395 => '1',
		5396 => '0',
		5397 => '1',
		5398 => '0',
		5399 => '1',
		5400 => '0',
		5401 => '1',
		5402 => '0',
		5403 => '1',
		5404 => '0',
		5405 => '1',
		5406 => '0',
		5407 => '1',
		5408 => '0',
		5409 => '1',
		5410 => '0',
		5411 => '1',
		5412 => '0',
		5413 => '1',
		5414 => '0',
		5415 => '1',
		5416 => '0',
		5417 => '1',
		5418 => '0',
		5419 => '1',
		5420 => '0',
		5421 => '1',
		5422 => '0',
		5423 => '1',
		5424 => '0',
		5425 => '1',
		5426 => '0',
		5427 => '1',
		5428 => '0',
		5429 => '1',
		5430 => '0',
		5431 => '1',
		5432 => '0',
		5433 => '1',
		5434 => '0',
		5435 => '1',
		5436 => '0',
		5437 => '1',
		5438 => '0',
		5439 => '1',
		5440 => '0',
		5441 => '1',
		5442 => '0',
		5443 => '1',
		5444 => '0',
		5445 => '1',
		5446 => '0',
		5447 => '1',
		5448 => '0',
		5449 => '1',
		5450 => '0',
		5451 => '1',
		5452 => '0',
		5453 => '1',
		5454 => '0',
		5455 => '1',
		5456 => '0',
		5457 => '1',
		5458 => '0',
		5459 => '1',
		5460 => '0',
		5461 => '1',
		5462 => '0',
		5463 => '1',
		5464 => '0',
		5465 => '1',
		5466 => '0',
		5467 => '1',
		5468 => '0',
		5469 => '1',
		5470 => '0',
		5471 => '1',
		5472 => '0',
		5473 => '1',
		5474 => '0',
		5475 => '1',
		5476 => '0',
		5477 => '1',
		5478 => '0',
		5479 => '1',
		5480 => '0',
		5481 => '1',
		5482 => '0',
		5483 => '1',
		5484 => '0',
		5485 => '1',
		5486 => '0',
		5487 => '1',
		5488 => '0',
		5489 => '1',
		5490 => '0',
		5491 => '1',
		5492 => '0',
		5493 => '1',
		5494 => '0',
		5495 => '1',
		5504 => '1',
		5505 => '0',
		5506 => '1',
		5507 => '0',
		5508 => '1',
		5509 => '0',
		5510 => '1',
		5511 => '0',
		5512 => '1',
		5513 => '0',
		5514 => '1',
		5515 => '0',
		5516 => '1',
		5517 => '0',
		5518 => '1',
		5519 => '0',
		5520 => '1',
		5521 => '0',
		5522 => '1',
		5523 => '0',
		5524 => '1',
		5525 => '0',
		5526 => '1',
		5527 => '0',
		5528 => '1',
		5529 => '0',
		5530 => '1',
		5531 => '0',
		5532 => '1',
		5533 => '0',
		5534 => '1',
		5535 => '0',
		5536 => '1',
		5537 => '0',
		5538 => '1',
		5539 => '0',
		5540 => '1',
		5541 => '0',
		5542 => '1',
		5543 => '0',
		5544 => '1',
		5545 => '0',
		5546 => '1',
		5547 => '0',
		5548 => '1',
		5549 => '0',
		5550 => '1',
		5551 => '0',
		5552 => '1',
		5553 => '0',
		5554 => '1',
		5555 => '0',
		5556 => '1',
		5557 => '0',
		5558 => '1',
		5559 => '0',
		5560 => '1',
		5561 => '0',
		5562 => '1',
		5563 => '0',
		5564 => '1',
		5565 => '0',
		5566 => '1',
		5567 => '0',
		5568 => '1',
		5569 => '0',
		5570 => '1',
		5571 => '0',
		5572 => '1',
		5573 => '0',
		5574 => '1',
		5575 => '0',
		5576 => '1',
		5577 => '0',
		5578 => '1',
		5579 => '0',
		5580 => '1',
		5581 => '0',
		5582 => '1',
		5583 => '0',
		5584 => '1',
		5585 => '0',
		5586 => '1',
		5587 => '0',
		5588 => '1',
		5589 => '0',
		5590 => '1',
		5591 => '0',
		5592 => '1',
		5593 => '0',
		5594 => '1',
		5595 => '0',
		5596 => '1',
		5597 => '0',
		5598 => '1',
		5599 => '0',
		5600 => '1',
		5601 => '0',
		5602 => '1',
		5603 => '0',
		5604 => '1',
		5605 => '0',
		5606 => '1',
		5607 => '0',
		5608 => '1',
		5609 => '0',
		5610 => '1',
		5611 => '0',
		5612 => '1',
		5613 => '0',
		5614 => '1',
		5615 => '0',
		5616 => '1',
		5617 => '0',
		5618 => '1',
		5619 => '0',
		5620 => '1',
		5621 => '0',
		5622 => '1',
		5623 => '0',
		5632 => '0',
		5633 => '1',
		5634 => '0',
		5635 => '1',
		5636 => '0',
		5637 => '1',
		5638 => '0',
		5639 => '1',
		5640 => '0',
		5641 => '1',
		5642 => '0',
		5643 => '1',
		5644 => '0',
		5645 => '1',
		5646 => '0',
		5647 => '1',
		5648 => '0',
		5649 => '1',
		5650 => '0',
		5651 => '1',
		5652 => '0',
		5653 => '1',
		5654 => '0',
		5655 => '1',
		5656 => '0',
		5657 => '1',
		5658 => '0',
		5659 => '1',
		5660 => '0',
		5661 => '1',
		5662 => '0',
		5663 => '1',
		5664 => '0',
		5665 => '1',
		5666 => '0',
		5667 => '1',
		5668 => '0',
		5669 => '1',
		5670 => '0',
		5671 => '1',
		5672 => '0',
		5673 => '1',
		5674 => '0',
		5675 => '1',
		5676 => '0',
		5677 => '1',
		5678 => '0',
		5679 => '1',
		5680 => '0',
		5681 => '1',
		5682 => '0',
		5683 => '1',
		5684 => '0',
		5685 => '1',
		5686 => '0',
		5687 => '1',
		5688 => '0',
		5689 => '1',
		5690 => '0',
		5691 => '1',
		5692 => '0',
		5693 => '1',
		5694 => '0',
		5695 => '1',
		5696 => '0',
		5697 => '1',
		5698 => '0',
		5699 => '1',
		5700 => '0',
		5701 => '1',
		5702 => '0',
		5703 => '1',
		5704 => '0',
		5705 => '1',
		5706 => '0',
		5707 => '1',
		5708 => '0',
		5709 => '1',
		5710 => '0',
		5711 => '1',
		5712 => '0',
		5713 => '1',
		5714 => '0',
		5715 => '1',
		5716 => '0',
		5717 => '1',
		5718 => '0',
		5719 => '1',
		5720 => '0',
		5721 => '1',
		5722 => '0',
		5723 => '1',
		5724 => '0',
		5725 => '1',
		5726 => '0',
		5727 => '1',
		5728 => '0',
		5729 => '1',
		5730 => '0',
		5731 => '1',
		5732 => '0',
		5733 => '1',
		5734 => '0',
		5735 => '1',
		5736 => '0',
		5737 => '1',
		5738 => '0',
		5739 => '1',
		5740 => '0',
		5741 => '1',
		5742 => '0',
		5743 => '1',
		5744 => '0',
		5745 => '1',
		5746 => '0',
		5747 => '1',
		5748 => '0',
		5749 => '1',
		5750 => '0',
		5751 => '1',
		5760 => '1',
		5761 => '0',
		5762 => '1',
		5763 => '0',
		5764 => '1',
		5765 => '0',
		5766 => '1',
		5767 => '0',
		5768 => '1',
		5769 => '0',
		5770 => '1',
		5771 => '0',
		5772 => '1',
		5773 => '0',
		5774 => '1',
		5775 => '0',
		5776 => '1',
		5777 => '0',
		5778 => '1',
		5779 => '0',
		5780 => '1',
		5781 => '0',
		5782 => '1',
		5783 => '0',
		5784 => '1',
		5785 => '0',
		5786 => '1',
		5787 => '0',
		5788 => '1',
		5789 => '0',
		5790 => '1',
		5791 => '0',
		5792 => '1',
		5793 => '0',
		5794 => '1',
		5795 => '0',
		5796 => '1',
		5797 => '0',
		5798 => '1',
		5799 => '0',
		5800 => '1',
		5801 => '0',
		5802 => '1',
		5803 => '0',
		5804 => '1',
		5805 => '0',
		5806 => '1',
		5807 => '0',
		5808 => '1',
		5809 => '0',
		5810 => '1',
		5811 => '0',
		5812 => '1',
		5813 => '0',
		5814 => '1',
		5815 => '0',
		5816 => '1',
		5817 => '0',
		5818 => '1',
		5819 => '0',
		5820 => '1',
		5821 => '0',
		5822 => '1',
		5823 => '0',
		5824 => '1',
		5825 => '0',
		5826 => '1',
		5827 => '0',
		5828 => '1',
		5829 => '0',
		5830 => '1',
		5831 => '0',
		5832 => '1',
		5833 => '0',
		5834 => '1',
		5835 => '0',
		5836 => '1',
		5837 => '0',
		5838 => '1',
		5839 => '0',
		5840 => '1',
		5841 => '0',
		5842 => '1',
		5843 => '0',
		5844 => '1',
		5845 => '0',
		5846 => '1',
		5847 => '0',
		5848 => '1',
		5849 => '0',
		5850 => '1',
		5851 => '0',
		5852 => '1',
		5853 => '0',
		5854 => '1',
		5855 => '0',
		5856 => '1',
		5857 => '0',
		5858 => '1',
		5859 => '0',
		5860 => '1',
		5861 => '0',
		5862 => '1',
		5863 => '0',
		5864 => '1',
		5865 => '0',
		5866 => '1',
		5867 => '0',
		5868 => '1',
		5869 => '0',
		5870 => '1',
		5871 => '0',
		5872 => '1',
		5873 => '0',
		5874 => '1',
		5875 => '0',
		5876 => '1',
		5877 => '0',
		5878 => '1',
		5879 => '0',
		5888 => '0',
		5889 => '1',
		5890 => '0',
		5891 => '1',
		5892 => '0',
		5893 => '1',
		5894 => '0',
		5895 => '1',
		5896 => '0',
		5897 => '1',
		5898 => '0',
		5899 => '1',
		5900 => '0',
		5901 => '1',
		5902 => '0',
		5903 => '1',
		5904 => '0',
		5905 => '1',
		5906 => '0',
		5907 => '1',
		5908 => '0',
		5909 => '1',
		5910 => '0',
		5911 => '1',
		5912 => '0',
		5913 => '1',
		5914 => '0',
		5915 => '1',
		5916 => '0',
		5917 => '1',
		5918 => '0',
		5919 => '1',
		5920 => '0',
		5921 => '1',
		5922 => '0',
		5923 => '1',
		5924 => '0',
		5925 => '1',
		5926 => '0',
		5927 => '1',
		5928 => '0',
		5929 => '1',
		5930 => '0',
		5931 => '1',
		5932 => '0',
		5933 => '1',
		5934 => '0',
		5935 => '1',
		5936 => '0',
		5937 => '1',
		5938 => '0',
		5939 => '1',
		5940 => '0',
		5941 => '1',
		5942 => '0',
		5943 => '1',
		5944 => '0',
		5945 => '1',
		5946 => '0',
		5947 => '1',
		5948 => '0',
		5949 => '1',
		5950 => '0',
		5951 => '1',
		5952 => '0',
		5953 => '1',
		5954 => '0',
		5955 => '1',
		5956 => '0',
		5957 => '1',
		5958 => '0',
		5959 => '1',
		5960 => '0',
		5961 => '1',
		5962 => '0',
		5963 => '1',
		5964 => '0',
		5965 => '1',
		5966 => '0',
		5967 => '1',
		5968 => '0',
		5969 => '1',
		5970 => '0',
		5971 => '1',
		5972 => '0',
		5973 => '1',
		5974 => '0',
		5975 => '1',
		5976 => '0',
		5977 => '1',
		5978 => '0',
		5979 => '1',
		5980 => '0',
		5981 => '1',
		5982 => '0',
		5983 => '1',
		5984 => '0',
		5985 => '1',
		5986 => '0',
		5987 => '1',
		5988 => '0',
		5989 => '1',
		5990 => '0',
		5991 => '1',
		5992 => '0',
		5993 => '1',
		5994 => '0',
		5995 => '1',
		5996 => '0',
		5997 => '1',
		5998 => '0',
		5999 => '1',
		6000 => '0',
		6001 => '1',
		6002 => '0',
		6003 => '1',
		6004 => '0',
		6005 => '1',
		6006 => '0',
		6007 => '1',
		6016 => '1',
		6017 => '0',
		6018 => '1',
		6019 => '0',
		6020 => '1',
		6021 => '0',
		6022 => '1',
		6023 => '0',
		6024 => '1',
		6025 => '0',
		6026 => '1',
		6027 => '0',
		6028 => '1',
		6029 => '0',
		6030 => '1',
		6031 => '0',
		6032 => '1',
		6033 => '0',
		6034 => '1',
		6035 => '0',
		6036 => '1',
		6037 => '0',
		6038 => '1',
		6039 => '0',
		6040 => '1',
		6041 => '0',
		6042 => '1',
		6043 => '0',
		6044 => '1',
		6045 => '0',
		6046 => '1',
		6047 => '0',
		6048 => '1',
		6049 => '0',
		6050 => '1',
		6051 => '0',
		6052 => '1',
		6053 => '0',
		6054 => '1',
		6055 => '0',
		6056 => '1',
		6057 => '0',
		6058 => '1',
		6059 => '0',
		6060 => '1',
		6061 => '0',
		6062 => '1',
		6063 => '0',
		6064 => '1',
		6065 => '0',
		6066 => '1',
		6067 => '0',
		6068 => '1',
		6069 => '0',
		6070 => '1',
		6071 => '0',
		6072 => '1',
		6073 => '0',
		6074 => '1',
		6075 => '0',
		6076 => '1',
		6077 => '0',
		6078 => '1',
		6079 => '0',
		6080 => '1',
		6081 => '0',
		6082 => '1',
		6083 => '0',
		6084 => '1',
		6085 => '0',
		6086 => '1',
		6087 => '0',
		6088 => '1',
		6089 => '0',
		6090 => '1',
		6091 => '0',
		6092 => '1',
		6093 => '0',
		6094 => '1',
		6095 => '0',
		6096 => '1',
		6097 => '0',
		6098 => '1',
		6099 => '0',
		6100 => '1',
		6101 => '0',
		6102 => '1',
		6103 => '0',
		6104 => '1',
		6105 => '0',
		6106 => '1',
		6107 => '0',
		6108 => '1',
		6109 => '0',
		6110 => '1',
		6111 => '0',
		6112 => '1',
		6113 => '0',
		6114 => '1',
		6115 => '0',
		6116 => '1',
		6117 => '0',
		6118 => '1',
		6119 => '0',
		6120 => '1',
		6121 => '0',
		6122 => '1',
		6123 => '0',
		6124 => '1',
		6125 => '0',
		6126 => '1',
		6127 => '0',
		6128 => '1',
		6129 => '0',
		6130 => '1',
		6131 => '0',
		6132 => '1',
		6133 => '0',
		6134 => '1',
		6135 => '0',
		6144 => '0',
		6145 => '1',
		6146 => '0',
		6147 => '1',
		6148 => '0',
		6149 => '1',
		6150 => '0',
		6151 => '1',
		6152 => '0',
		6153 => '1',
		6154 => '0',
		6155 => '1',
		6156 => '0',
		6157 => '1',
		6158 => '0',
		6159 => '1',
		6160 => '0',
		6161 => '1',
		6162 => '0',
		6163 => '1',
		6164 => '0',
		6165 => '1',
		6166 => '0',
		6167 => '1',
		6168 => '0',
		6169 => '1',
		6170 => '0',
		6171 => '1',
		6172 => '0',
		6173 => '1',
		6174 => '0',
		6175 => '1',
		6176 => '0',
		6177 => '1',
		6178 => '0',
		6179 => '1',
		6180 => '0',
		6181 => '1',
		6182 => '0',
		6183 => '1',
		6184 => '0',
		6185 => '1',
		6186 => '0',
		6187 => '1',
		6188 => '0',
		6189 => '1',
		6190 => '0',
		6191 => '1',
		6192 => '0',
		6193 => '1',
		6194 => '0',
		6195 => '1',
		6196 => '0',
		6197 => '1',
		6198 => '0',
		6199 => '1',
		6200 => '0',
		6201 => '1',
		6202 => '0',
		6203 => '1',
		6204 => '0',
		6205 => '1',
		6206 => '0',
		6207 => '1',
		6208 => '0',
		6209 => '1',
		6210 => '0',
		6211 => '1',
		6212 => '0',
		6213 => '1',
		6214 => '0',
		6215 => '1',
		6216 => '0',
		6217 => '1',
		6218 => '0',
		6219 => '1',
		6220 => '0',
		6221 => '1',
		6222 => '0',
		6223 => '1',
		6224 => '0',
		6225 => '1',
		6226 => '0',
		6227 => '1',
		6228 => '0',
		6229 => '1',
		6230 => '0',
		6231 => '1',
		6232 => '0',
		6233 => '1',
		6234 => '0',
		6235 => '1',
		6236 => '0',
		6237 => '1',
		6238 => '0',
		6239 => '1',
		6240 => '0',
		6241 => '1',
		6242 => '0',
		6243 => '1',
		6244 => '0',
		6245 => '1',
		6246 => '0',
		6247 => '1',
		6248 => '0',
		6249 => '1',
		6250 => '0',
		6251 => '1',
		6252 => '0',
		6253 => '1',
		6254 => '0',
		6255 => '1',
		6256 => '0',
		6257 => '1',
		6258 => '0',
		6259 => '1',
		6260 => '0',
		6261 => '1',
		6262 => '0',
		6263 => '1',
		6272 => '1',
		6273 => '0',
		6274 => '1',
		6275 => '0',
		6276 => '1',
		6277 => '0',
		6278 => '1',
		6279 => '0',
		6280 => '1',
		6281 => '0',
		6282 => '1',
		6283 => '0',
		6284 => '1',
		6285 => '0',
		6286 => '1',
		6287 => '0',
		6288 => '1',
		6289 => '0',
		6290 => '1',
		6291 => '0',
		6292 => '1',
		6293 => '0',
		6294 => '1',
		6295 => '0',
		6296 => '1',
		6297 => '0',
		6298 => '1',
		6299 => '0',
		6300 => '1',
		6301 => '0',
		6302 => '1',
		6303 => '0',
		6304 => '1',
		6305 => '0',
		6306 => '1',
		6307 => '0',
		6308 => '1',
		6309 => '0',
		6310 => '1',
		6311 => '0',
		6312 => '1',
		6313 => '0',
		6314 => '1',
		6315 => '0',
		6316 => '1',
		6317 => '0',
		6318 => '1',
		6319 => '0',
		6320 => '1',
		6321 => '0',
		6322 => '1',
		6323 => '0',
		6324 => '1',
		6325 => '0',
		6326 => '1',
		6327 => '0',
		6328 => '1',
		6329 => '0',
		6330 => '1',
		6331 => '0',
		6332 => '1',
		6333 => '0',
		6334 => '1',
		6335 => '0',
		6336 => '1',
		6337 => '0',
		6338 => '1',
		6339 => '0',
		6340 => '1',
		6341 => '0',
		6342 => '1',
		6343 => '0',
		6344 => '1',
		6345 => '0',
		6346 => '1',
		6347 => '0',
		6348 => '1',
		6349 => '0',
		6350 => '1',
		6351 => '0',
		6352 => '1',
		6353 => '0',
		6354 => '1',
		6355 => '0',
		6356 => '1',
		6357 => '0',
		6358 => '1',
		6359 => '0',
		6360 => '1',
		6361 => '0',
		6362 => '1',
		6363 => '0',
		6364 => '1',
		6365 => '0',
		6366 => '1',
		6367 => '0',
		6368 => '1',
		6369 => '0',
		6370 => '1',
		6371 => '0',
		6372 => '1',
		6373 => '0',
		6374 => '1',
		6375 => '0',
		6376 => '1',
		6377 => '0',
		6378 => '1',
		6379 => '0',
		6380 => '1',
		6381 => '0',
		6382 => '1',
		6383 => '0',
		6384 => '1',
		6385 => '0',
		6386 => '1',
		6387 => '0',
		6388 => '1',
		6389 => '0',
		6390 => '1',
		6391 => '0',
		6400 => '0',
		6401 => '1',
		6402 => '0',
		6403 => '1',
		6404 => '0',
		6405 => '1',
		6406 => '0',
		6407 => '1',
		6408 => '0',
		6409 => '1',
		6410 => '0',
		6411 => '1',
		6412 => '0',
		6413 => '1',
		6414 => '0',
		6415 => '1',
		6416 => '0',
		6417 => '1',
		6418 => '0',
		6419 => '1',
		6420 => '0',
		6421 => '1',
		6422 => '0',
		6423 => '1',
		6424 => '0',
		6425 => '1',
		6426 => '0',
		6427 => '1',
		6428 => '0',
		6429 => '1',
		6430 => '0',
		6431 => '1',
		6432 => '0',
		6433 => '1',
		6434 => '0',
		6435 => '1',
		6436 => '0',
		6437 => '1',
		6438 => '0',
		6439 => '1',
		6440 => '0',
		6441 => '1',
		6442 => '0',
		6443 => '1',
		6444 => '0',
		6445 => '1',
		6446 => '0',
		6447 => '1',
		6448 => '0',
		6449 => '1',
		6450 => '0',
		6451 => '1',
		6452 => '0',
		6453 => '1',
		6454 => '0',
		6455 => '1',
		6456 => '0',
		6457 => '1',
		6458 => '0',
		6459 => '1',
		6460 => '0',
		6461 => '1',
		6462 => '0',
		6463 => '1',
		6464 => '0',
		6465 => '1',
		6466 => '0',
		6467 => '1',
		6468 => '0',
		6469 => '1',
		6470 => '0',
		6471 => '1',
		6472 => '0',
		6473 => '1',
		6474 => '0',
		6475 => '1',
		6476 => '0',
		6477 => '1',
		6478 => '0',
		6479 => '1',
		6480 => '0',
		6481 => '1',
		6482 => '0',
		6483 => '1',
		6484 => '0',
		6485 => '1',
		6486 => '0',
		6487 => '1',
		6488 => '0',
		6489 => '1',
		6490 => '0',
		6491 => '1',
		6492 => '0',
		6493 => '1',
		6494 => '0',
		6495 => '1',
		6496 => '0',
		6497 => '1',
		6498 => '0',
		6499 => '1',
		6500 => '0',
		6501 => '1',
		6502 => '0',
		6503 => '1',
		6504 => '0',
		6505 => '1',
		6506 => '0',
		6507 => '1',
		6508 => '0',
		6509 => '1',
		6510 => '0',
		6511 => '1',
		6512 => '0',
		6513 => '1',
		6514 => '0',
		6515 => '1',
		6516 => '0',
		6517 => '1',
		6518 => '0',
		6519 => '1',
		6528 => '1',
		6529 => '0',
		6530 => '1',
		6531 => '0',
		6532 => '1',
		6533 => '0',
		6534 => '1',
		6535 => '0',
		6536 => '1',
		6537 => '0',
		6538 => '1',
		6539 => '0',
		6540 => '1',
		6541 => '0',
		6542 => '1',
		6543 => '0',
		6544 => '1',
		6545 => '0',
		6546 => '1',
		6547 => '0',
		6548 => '1',
		6549 => '0',
		6550 => '1',
		6551 => '0',
		6552 => '1',
		6553 => '0',
		6554 => '1',
		6555 => '0',
		6556 => '1',
		6557 => '0',
		6558 => '1',
		6559 => '0',
		6560 => '1',
		6561 => '0',
		6562 => '1',
		6563 => '0',
		6564 => '1',
		6565 => '0',
		6566 => '1',
		6567 => '0',
		6568 => '1',
		6569 => '0',
		6570 => '1',
		6571 => '0',
		6572 => '1',
		6573 => '0',
		6574 => '1',
		6575 => '0',
		6576 => '1',
		6577 => '0',
		6578 => '1',
		6579 => '0',
		6580 => '1',
		6581 => '0',
		6582 => '1',
		6583 => '0',
		6584 => '1',
		6585 => '0',
		6586 => '1',
		6587 => '0',
		6588 => '1',
		6589 => '0',
		6590 => '1',
		6591 => '0',
		6592 => '1',
		6593 => '0',
		6594 => '1',
		6595 => '0',
		6596 => '1',
		6597 => '0',
		6598 => '1',
		6599 => '0',
		6600 => '1',
		6601 => '0',
		6602 => '1',
		6603 => '0',
		6604 => '1',
		6605 => '0',
		6606 => '1',
		6607 => '0',
		6608 => '1',
		6609 => '0',
		6610 => '1',
		6611 => '0',
		6612 => '1',
		6613 => '0',
		6614 => '1',
		6615 => '0',
		6616 => '1',
		6617 => '0',
		6618 => '1',
		6619 => '0',
		6620 => '1',
		6621 => '0',
		6622 => '1',
		6623 => '0',
		6624 => '1',
		6625 => '0',
		6626 => '1',
		6627 => '0',
		6628 => '1',
		6629 => '0',
		6630 => '1',
		6631 => '0',
		6632 => '1',
		6633 => '0',
		6634 => '1',
		6635 => '0',
		6636 => '1',
		6637 => '0',
		6638 => '1',
		6639 => '0',
		6640 => '1',
		6641 => '0',
		6642 => '1',
		6643 => '0',
		6644 => '1',
		6645 => '0',
		6646 => '1',
		6647 => '0',
		6656 => '0',
		6657 => '1',
		6658 => '0',
		6659 => '1',
		6660 => '0',
		6661 => '1',
		6662 => '0',
		6663 => '1',
		6664 => '0',
		6665 => '1',
		6666 => '0',
		6667 => '1',
		6668 => '0',
		6669 => '1',
		6670 => '0',
		6671 => '1',
		6672 => '0',
		6673 => '1',
		6674 => '0',
		6675 => '1',
		6676 => '0',
		6677 => '1',
		6678 => '0',
		6679 => '1',
		6680 => '0',
		6681 => '1',
		6682 => '0',
		6683 => '1',
		6684 => '0',
		6685 => '1',
		6686 => '0',
		6687 => '1',
		6688 => '0',
		6689 => '1',
		6690 => '0',
		6691 => '1',
		6692 => '0',
		6693 => '1',
		6694 => '0',
		6695 => '1',
		6696 => '0',
		6697 => '1',
		6698 => '0',
		6699 => '1',
		6700 => '0',
		6701 => '1',
		6702 => '0',
		6703 => '1',
		6704 => '0',
		6705 => '1',
		6706 => '0',
		6707 => '1',
		6708 => '0',
		6709 => '1',
		6710 => '0',
		6711 => '1',
		6712 => '0',
		6713 => '1',
		6714 => '0',
		6715 => '1',
		6716 => '0',
		6717 => '1',
		6718 => '0',
		6719 => '1',
		6720 => '0',
		6721 => '1',
		6722 => '0',
		6723 => '1',
		6724 => '0',
		6725 => '1',
		6726 => '0',
		6727 => '1',
		6728 => '0',
		6729 => '1',
		6730 => '0',
		6731 => '1',
		6732 => '0',
		6733 => '1',
		6734 => '0',
		6735 => '1',
		6736 => '0',
		6737 => '1',
		6738 => '0',
		6739 => '1',
		6740 => '0',
		6741 => '1',
		6742 => '0',
		6743 => '1',
		6744 => '0',
		6745 => '1',
		6746 => '0',
		6747 => '1',
		6748 => '0',
		6749 => '1',
		6750 => '0',
		6751 => '1',
		6752 => '0',
		6753 => '1',
		6754 => '0',
		6755 => '1',
		6756 => '0',
		6757 => '1',
		6758 => '0',
		6759 => '1',
		6760 => '0',
		6761 => '1',
		6762 => '0',
		6763 => '1',
		6764 => '0',
		6765 => '1',
		6766 => '0',
		6767 => '1',
		6768 => '0',
		6769 => '1',
		6770 => '0',
		6771 => '1',
		6772 => '0',
		6773 => '1',
		6774 => '0',
		6775 => '1',
		6784 => '1',
		6785 => '0',
		6786 => '1',
		6787 => '0',
		6788 => '1',
		6789 => '0',
		6790 => '1',
		6791 => '0',
		6792 => '1',
		6793 => '0',
		6794 => '1',
		6795 => '0',
		6796 => '1',
		6797 => '0',
		6798 => '1',
		6799 => '0',
		6800 => '1',
		6801 => '0',
		6802 => '1',
		6803 => '0',
		6804 => '1',
		6805 => '0',
		6806 => '1',
		6807 => '0',
		6808 => '1',
		6809 => '0',
		6810 => '1',
		6811 => '0',
		6812 => '1',
		6813 => '0',
		6814 => '1',
		6815 => '0',
		6816 => '1',
		6817 => '0',
		6818 => '1',
		6819 => '0',
		6820 => '1',
		6821 => '0',
		6822 => '1',
		6823 => '0',
		6824 => '1',
		6825 => '0',
		6826 => '1',
		6827 => '0',
		6828 => '1',
		6829 => '0',
		6830 => '1',
		6831 => '0',
		6832 => '1',
		6833 => '0',
		6834 => '1',
		6835 => '0',
		6836 => '1',
		6837 => '0',
		6838 => '1',
		6839 => '0',
		6840 => '1',
		6841 => '0',
		6842 => '1',
		6843 => '0',
		6844 => '1',
		6845 => '0',
		6846 => '1',
		6847 => '0',
		6848 => '1',
		6849 => '0',
		6850 => '1',
		6851 => '0',
		6852 => '1',
		6853 => '0',
		6854 => '1',
		6855 => '0',
		6856 => '1',
		6857 => '0',
		6858 => '1',
		6859 => '0',
		6860 => '1',
		6861 => '0',
		6862 => '1',
		6863 => '0',
		6864 => '1',
		6865 => '0',
		6866 => '1',
		6867 => '0',
		6868 => '1',
		6869 => '0',
		6870 => '1',
		6871 => '0',
		6872 => '1',
		6873 => '0',
		6874 => '1',
		6875 => '0',
		6876 => '1',
		6877 => '0',
		6878 => '1',
		6879 => '0',
		6880 => '1',
		6881 => '0',
		6882 => '1',
		6883 => '0',
		6884 => '1',
		6885 => '0',
		6886 => '1',
		6887 => '0',
		6888 => '1',
		6889 => '0',
		6890 => '1',
		6891 => '0',
		6892 => '1',
		6893 => '0',
		6894 => '1',
		6895 => '0',
		6896 => '1',
		6897 => '0',
		6898 => '1',
		6899 => '0',
		6900 => '1',
		6901 => '0',
		6902 => '1',
		6903 => '0',
		6912 => '0',
		6913 => '1',
		6914 => '0',
		6915 => '1',
		6916 => '0',
		6917 => '1',
		6918 => '0',
		6919 => '1',
		6920 => '0',
		6921 => '1',
		6922 => '0',
		6923 => '1',
		6924 => '0',
		6925 => '1',
		6926 => '0',
		6927 => '1',
		6928 => '0',
		6929 => '1',
		6930 => '0',
		6931 => '1',
		6932 => '0',
		6933 => '1',
		6934 => '0',
		6935 => '1',
		6936 => '0',
		6937 => '1',
		6938 => '0',
		6939 => '1',
		6940 => '0',
		6941 => '1',
		6942 => '0',
		6943 => '1',
		6944 => '0',
		6945 => '1',
		6946 => '0',
		6947 => '1',
		6948 => '0',
		6949 => '1',
		6950 => '0',
		6951 => '1',
		6952 => '0',
		6953 => '1',
		6954 => '0',
		6955 => '1',
		6956 => '0',
		6957 => '1',
		6958 => '0',
		6959 => '1',
		6960 => '0',
		6961 => '1',
		6962 => '0',
		6963 => '1',
		6964 => '0',
		6965 => '1',
		6966 => '0',
		6967 => '1',
		6968 => '0',
		6969 => '1',
		6970 => '0',
		6971 => '1',
		6972 => '0',
		6973 => '1',
		6974 => '0',
		6975 => '1',
		6976 => '0',
		6977 => '1',
		6978 => '0',
		6979 => '1',
		6980 => '0',
		6981 => '1',
		6982 => '0',
		6983 => '1',
		6984 => '0',
		6985 => '1',
		6986 => '0',
		6987 => '1',
		6988 => '0',
		6989 => '1',
		6990 => '0',
		6991 => '1',
		6992 => '0',
		6993 => '1',
		6994 => '0',
		6995 => '1',
		6996 => '0',
		6997 => '1',
		6998 => '0',
		6999 => '1',
		7000 => '0',
		7001 => '1',
		7002 => '0',
		7003 => '1',
		7004 => '0',
		7005 => '1',
		7006 => '0',
		7007 => '1',
		7008 => '0',
		7009 => '1',
		7010 => '0',
		7011 => '1',
		7012 => '0',
		7013 => '1',
		7014 => '0',
		7015 => '1',
		7016 => '0',
		7017 => '1',
		7018 => '0',
		7019 => '1',
		7020 => '0',
		7021 => '1',
		7022 => '0',
		7023 => '1',
		7024 => '0',
		7025 => '1',
		7026 => '0',
		7027 => '1',
		7028 => '0',
		7029 => '1',
		7030 => '0',
		7031 => '1',
		7040 => '1',
		7041 => '0',
		7042 => '1',
		7043 => '0',
		7044 => '1',
		7045 => '0',
		7046 => '1',
		7047 => '0',
		7048 => '1',
		7049 => '0',
		7050 => '1',
		7051 => '0',
		7052 => '1',
		7053 => '0',
		7054 => '1',
		7055 => '0',
		7056 => '1',
		7057 => '0',
		7058 => '1',
		7059 => '0',
		7060 => '1',
		7061 => '0',
		7062 => '1',
		7063 => '0',
		7064 => '1',
		7065 => '0',
		7066 => '1',
		7067 => '0',
		7068 => '1',
		7069 => '0',
		7070 => '1',
		7071 => '0',
		7072 => '1',
		7073 => '0',
		7074 => '1',
		7075 => '0',
		7076 => '1',
		7077 => '0',
		7078 => '1',
		7079 => '0',
		7080 => '1',
		7081 => '0',
		7082 => '1',
		7083 => '0',
		7084 => '1',
		7085 => '0',
		7086 => '1',
		7087 => '0',
		7088 => '1',
		7089 => '0',
		7090 => '1',
		7091 => '0',
		7092 => '1',
		7093 => '0',
		7094 => '1',
		7095 => '0',
		7096 => '1',
		7097 => '0',
		7098 => '1',
		7099 => '0',
		7100 => '1',
		7101 => '0',
		7102 => '1',
		7103 => '0',
		7104 => '1',
		7105 => '0',
		7106 => '1',
		7107 => '0',
		7108 => '1',
		7109 => '0',
		7110 => '1',
		7111 => '0',
		7112 => '1',
		7113 => '0',
		7114 => '1',
		7115 => '0',
		7116 => '1',
		7117 => '0',
		7118 => '1',
		7119 => '0',
		7120 => '1',
		7121 => '0',
		7122 => '1',
		7123 => '0',
		7124 => '1',
		7125 => '0',
		7126 => '1',
		7127 => '0',
		7128 => '1',
		7129 => '0',
		7130 => '1',
		7131 => '0',
		7132 => '1',
		7133 => '0',
		7134 => '1',
		7135 => '0',
		7136 => '1',
		7137 => '0',
		7138 => '1',
		7139 => '0',
		7140 => '1',
		7141 => '0',
		7142 => '1',
		7143 => '0',
		7144 => '1',
		7145 => '0',
		7146 => '1',
		7147 => '0',
		7148 => '1',
		7149 => '0',
		7150 => '1',
		7151 => '0',
		7152 => '1',
		7153 => '0',
		7154 => '1',
		7155 => '0',
		7156 => '1',
		7157 => '0',
		7158 => '1',
		7159 => '0',
		7168 => '0',
		7169 => '1',
		7170 => '0',
		7171 => '1',
		7172 => '0',
		7173 => '1',
		7174 => '0',
		7175 => '1',
		7176 => '0',
		7177 => '1',
		7178 => '0',
		7179 => '1',
		7180 => '0',
		7181 => '1',
		7182 => '0',
		7183 => '1',
		7184 => '0',
		7185 => '1',
		7186 => '0',
		7187 => '1',
		7188 => '0',
		7189 => '1',
		7190 => '0',
		7191 => '1',
		7192 => '0',
		7193 => '1',
		7194 => '0',
		7195 => '1',
		7196 => '0',
		7197 => '1',
		7198 => '0',
		7199 => '1',
		7200 => '0',
		7201 => '1',
		7202 => '0',
		7203 => '1',
		7204 => '0',
		7205 => '1',
		7206 => '0',
		7207 => '1',
		7208 => '0',
		7209 => '1',
		7210 => '0',
		7211 => '1',
		7212 => '0',
		7213 => '1',
		7214 => '0',
		7215 => '1',
		7216 => '0',
		7217 => '1',
		7218 => '0',
		7219 => '1',
		7220 => '0',
		7221 => '1',
		7222 => '0',
		7223 => '1',
		7224 => '0',
		7225 => '1',
		7226 => '0',
		7227 => '1',
		7228 => '0',
		7229 => '1',
		7230 => '0',
		7231 => '1',
		7232 => '0',
		7233 => '1',
		7234 => '0',
		7235 => '1',
		7236 => '0',
		7237 => '1',
		7238 => '0',
		7239 => '1',
		7240 => '0',
		7241 => '1',
		7242 => '0',
		7243 => '1',
		7244 => '0',
		7245 => '1',
		7246 => '0',
		7247 => '1',
		7248 => '0',
		7249 => '1',
		7250 => '0',
		7251 => '1',
		7252 => '0',
		7253 => '1',
		7254 => '0',
		7255 => '1',
		7256 => '0',
		7257 => '1',
		7258 => '0',
		7259 => '1',
		7260 => '0',
		7261 => '1',
		7262 => '0',
		7263 => '1',
		7264 => '0',
		7265 => '1',
		7266 => '0',
		7267 => '1',
		7268 => '0',
		7269 => '1',
		7270 => '0',
		7271 => '1',
		7272 => '0',
		7273 => '1',
		7274 => '0',
		7275 => '1',
		7276 => '0',
		7277 => '1',
		7278 => '0',
		7279 => '1',
		7280 => '0',
		7281 => '1',
		7282 => '0',
		7283 => '1',
		7284 => '0',
		7285 => '1',
		7286 => '0',
		7287 => '1',
		7296 => '1',
		7297 => '0',
		7298 => '1',
		7299 => '0',
		7300 => '1',
		7301 => '0',
		7302 => '1',
		7303 => '0',
		7304 => '1',
		7305 => '0',
		7306 => '1',
		7307 => '0',
		7308 => '1',
		7309 => '0',
		7310 => '1',
		7311 => '0',
		7312 => '1',
		7313 => '0',
		7314 => '1',
		7315 => '0',
		7316 => '1',
		7317 => '0',
		7318 => '1',
		7319 => '0',
		7320 => '1',
		7321 => '0',
		7322 => '1',
		7323 => '0',
		7324 => '1',
		7325 => '0',
		7326 => '1',
		7327 => '0',
		7328 => '1',
		7329 => '0',
		7330 => '1',
		7331 => '0',
		7332 => '1',
		7333 => '0',
		7334 => '1',
		7335 => '0',
		7336 => '1',
		7337 => '0',
		7338 => '1',
		7339 => '0',
		7340 => '1',
		7341 => '0',
		7342 => '1',
		7343 => '0',
		7344 => '1',
		7345 => '0',
		7346 => '1',
		7347 => '0',
		7348 => '1',
		7349 => '0',
		7350 => '1',
		7351 => '0',
		7352 => '1',
		7353 => '0',
		7354 => '1',
		7355 => '0',
		7356 => '1',
		7357 => '0',
		7358 => '1',
		7359 => '0',
		7360 => '1',
		7361 => '0',
		7362 => '1',
		7363 => '0',
		7364 => '1',
		7365 => '0',
		7366 => '1',
		7367 => '0',
		7368 => '1',
		7369 => '0',
		7370 => '1',
		7371 => '0',
		7372 => '1',
		7373 => '0',
		7374 => '1',
		7375 => '0',
		7376 => '1',
		7377 => '0',
		7378 => '1',
		7379 => '0',
		7380 => '1',
		7381 => '0',
		7382 => '1',
		7383 => '0',
		7384 => '1',
		7385 => '0',
		7386 => '1',
		7387 => '0',
		7388 => '1',
		7389 => '0',
		7390 => '1',
		7391 => '0',
		7392 => '1',
		7393 => '0',
		7394 => '1',
		7395 => '0',
		7396 => '1',
		7397 => '0',
		7398 => '1',
		7399 => '0',
		7400 => '1',
		7401 => '0',
		7402 => '1',
		7403 => '0',
		7404 => '1',
		7405 => '0',
		7406 => '1',
		7407 => '0',
		7408 => '1',
		7409 => '0',
		7410 => '1',
		7411 => '0',
		7412 => '1',
		7413 => '0',
		7414 => '1',
		7415 => '0',
		7424 => '0',
		7425 => '1',
		7426 => '0',
		7427 => '1',
		7428 => '0',
		7429 => '1',
		7430 => '0',
		7431 => '1',
		7432 => '0',
		7433 => '1',
		7434 => '0',
		7435 => '1',
		7436 => '0',
		7437 => '1',
		7438 => '0',
		7439 => '1',
		7440 => '0',
		7441 => '1',
		7442 => '0',
		7443 => '1',
		7444 => '0',
		7445 => '1',
		7446 => '0',
		7447 => '1',
		7448 => '0',
		7449 => '1',
		7450 => '0',
		7451 => '1',
		7452 => '0',
		7453 => '1',
		7454 => '0',
		7455 => '1',
		7456 => '0',
		7457 => '1',
		7458 => '0',
		7459 => '1',
		7460 => '0',
		7461 => '1',
		7462 => '0',
		7463 => '1',
		7464 => '0',
		7465 => '1',
		7466 => '0',
		7467 => '1',
		7468 => '0',
		7469 => '1',
		7470 => '0',
		7471 => '1',
		7472 => '0',
		7473 => '1',
		7474 => '0',
		7475 => '1',
		7476 => '0',
		7477 => '1',
		7478 => '0',
		7479 => '1',
		7480 => '0',
		7481 => '1',
		7482 => '0',
		7483 => '1',
		7484 => '0',
		7485 => '1',
		7486 => '0',
		7487 => '1',
		7488 => '0',
		7489 => '1',
		7490 => '0',
		7491 => '1',
		7492 => '0',
		7493 => '1',
		7494 => '0',
		7495 => '1',
		7496 => '0',
		7497 => '1',
		7498 => '0',
		7499 => '1',
		7500 => '0',
		7501 => '1',
		7502 => '0',
		7503 => '1',
		7504 => '0',
		7505 => '1',
		7506 => '0',
		7507 => '1',
		7508 => '0',
		7509 => '1',
		7510 => '0',
		7511 => '1',
		7512 => '0',
		7513 => '1',
		7514 => '0',
		7515 => '1',
		7516 => '0',
		7517 => '1',
		7518 => '0',
		7519 => '1',
		7520 => '0',
		7521 => '1',
		7522 => '0',
		7523 => '1',
		7524 => '0',
		7525 => '1',
		7526 => '0',
		7527 => '1',
		7528 => '0',
		7529 => '1',
		7530 => '0',
		7531 => '1',
		7532 => '0',
		7533 => '1',
		7534 => '0',
		7535 => '1',
		7536 => '0',
		7537 => '1',
		7538 => '0',
		7539 => '1',
		7540 => '0',
		7541 => '1',
		7542 => '0',
		7543 => '1',
		7552 => '1',
		7553 => '0',
		7554 => '1',
		7555 => '0',
		7556 => '1',
		7557 => '0',
		7558 => '1',
		7559 => '0',
		7560 => '1',
		7561 => '0',
		7562 => '1',
		7563 => '0',
		7564 => '1',
		7565 => '0',
		7566 => '1',
		7567 => '0',
		7568 => '1',
		7569 => '0',
		7570 => '1',
		7571 => '0',
		7572 => '1',
		7573 => '0',
		7574 => '1',
		7575 => '0',
		7576 => '1',
		7577 => '0',
		7578 => '1',
		7579 => '0',
		7580 => '1',
		7581 => '0',
		7582 => '1',
		7583 => '0',
		7584 => '1',
		7585 => '0',
		7586 => '1',
		7587 => '0',
		7588 => '1',
		7589 => '0',
		7590 => '1',
		7591 => '0',
		7592 => '1',
		7593 => '0',
		7594 => '1',
		7595 => '0',
		7596 => '1',
		7597 => '0',
		7598 => '1',
		7599 => '0',
		7600 => '1',
		7601 => '0',
		7602 => '1',
		7603 => '0',
		7604 => '1',
		7605 => '0',
		7606 => '1',
		7607 => '0',
		7608 => '1',
		7609 => '0',
		7610 => '1',
		7611 => '0',
		7612 => '1',
		7613 => '0',
		7614 => '1',
		7615 => '0',
		7616 => '1',
		7617 => '0',
		7618 => '1',
		7619 => '0',
		7620 => '1',
		7621 => '0',
		7622 => '1',
		7623 => '0',
		7624 => '1',
		7625 => '0',
		7626 => '1',
		7627 => '0',
		7628 => '1',
		7629 => '0',
		7630 => '1',
		7631 => '0',
		7632 => '1',
		7633 => '0',
		7634 => '1',
		7635 => '0',
		7636 => '1',
		7637 => '0',
		7638 => '1',
		7639 => '0',
		7640 => '1',
		7641 => '0',
		7642 => '1',
		7643 => '0',
		7644 => '1',
		7645 => '0',
		7646 => '1',
		7647 => '0',
		7648 => '1',
		7649 => '0',
		7650 => '1',
		7651 => '0',
		7652 => '1',
		7653 => '0',
		7654 => '1',
		7655 => '0',
		7656 => '1',
		7657 => '0',
		7658 => '1',
		7659 => '0',
		7660 => '1',
		7661 => '0',
		7662 => '1',
		7663 => '0',
		7664 => '1',
		7665 => '0',
		7666 => '1',
		7667 => '0',
		7668 => '1',
		7669 => '0',
		7670 => '1',
		7671 => '0',
		7680 => '0',
		7681 => '1',
		7682 => '0',
		7683 => '1',
		7684 => '0',
		7685 => '1',
		7686 => '0',
		7687 => '1',
		7688 => '0',
		7689 => '1',
		7690 => '0',
		7691 => '1',
		7692 => '0',
		7693 => '1',
		7694 => '0',
		7695 => '1',
		7696 => '0',
		7697 => '1',
		7698 => '0',
		7699 => '1',
		7700 => '0',
		7701 => '1',
		7702 => '0',
		7703 => '1',
		7704 => '0',
		7705 => '1',
		7706 => '0',
		7707 => '1',
		7708 => '0',
		7709 => '1',
		7710 => '0',
		7711 => '1',
		7712 => '0',
		7713 => '1',
		7714 => '0',
		7715 => '1',
		7716 => '0',
		7717 => '1',
		7718 => '0',
		7719 => '1',
		7720 => '0',
		7721 => '1',
		7722 => '0',
		7723 => '1',
		7724 => '0',
		7725 => '1',
		7726 => '0',
		7727 => '1',
		7728 => '0',
		7729 => '1',
		7730 => '0',
		7731 => '1',
		7732 => '0',
		7733 => '1',
		7734 => '0',
		7735 => '1',
		7736 => '0',
		7737 => '1',
		7738 => '0',
		7739 => '1',
		7740 => '0',
		7741 => '1',
		7742 => '0',
		7743 => '1',
		7744 => '0',
		7745 => '1',
		7746 => '0',
		7747 => '1',
		7748 => '0',
		7749 => '1',
		7750 => '0',
		7751 => '1',
		7752 => '0',
		7753 => '1',
		7754 => '0',
		7755 => '1',
		7756 => '0',
		7757 => '1',
		7758 => '0',
		7759 => '1',
		7760 => '0',
		7761 => '1',
		7762 => '0',
		7763 => '1',
		7764 => '0',
		7765 => '1',
		7766 => '0',
		7767 => '1',
		7768 => '0',
		7769 => '1',
		7770 => '0',
		7771 => '1',
		7772 => '0',
		7773 => '1',
		7774 => '0',
		7775 => '1',
		7776 => '0',
		7777 => '1',
		7778 => '0',
		7779 => '1',
		7780 => '0',
		7781 => '1',
		7782 => '0',
		7783 => '1',
		7784 => '0',
		7785 => '1',
		7786 => '0',
		7787 => '1',
		7788 => '0',
		7789 => '1',
		7790 => '0',
		7791 => '1',
		7792 => '0',
		7793 => '1',
		7794 => '0',
		7795 => '1',
		7796 => '0',
		7797 => '1',
		7798 => '0',
		7799 => '1',
		7808 => '1',
		7809 => '0',
		7810 => '1',
		7811 => '0',
		7812 => '1',
		7813 => '0',
		7814 => '1',
		7815 => '0',
		7816 => '1',
		7817 => '0',
		7818 => '1',
		7819 => '0',
		7820 => '1',
		7821 => '0',
		7822 => '1',
		7823 => '0',
		7824 => '1',
		7825 => '0',
		7826 => '1',
		7827 => '0',
		7828 => '1',
		7829 => '0',
		7830 => '1',
		7831 => '0',
		7832 => '1',
		7833 => '0',
		7834 => '1',
		7835 => '0',
		7836 => '1',
		7837 => '0',
		7838 => '1',
		7839 => '0',
		7840 => '1',
		7841 => '0',
		7842 => '1',
		7843 => '0',
		7844 => '1',
		7845 => '0',
		7846 => '1',
		7847 => '0',
		7848 => '1',
		7849 => '0',
		7850 => '1',
		7851 => '0',
		7852 => '1',
		7853 => '0',
		7854 => '1',
		7855 => '0',
		7856 => '1',
		7857 => '0',
		7858 => '1',
		7859 => '0',
		7860 => '1',
		7861 => '0',
		7862 => '1',
		7863 => '0',
		7864 => '1',
		7865 => '0',
		7866 => '1',
		7867 => '0',
		7868 => '1',
		7869 => '0',
		7870 => '1',
		7871 => '0',
		7872 => '1',
		7873 => '0',
		7874 => '1',
		7875 => '0',
		7876 => '1',
		7877 => '0',
		7878 => '1',
		7879 => '0',
		7880 => '1',
		7881 => '0',
		7882 => '1',
		7883 => '0',
		7884 => '1',
		7885 => '0',
		7886 => '1',
		7887 => '0',
		7888 => '1',
		7889 => '0',
		7890 => '1',
		7891 => '0',
		7892 => '1',
		7893 => '0',
		7894 => '1',
		7895 => '0',
		7896 => '1',
		7897 => '0',
		7898 => '1',
		7899 => '0',
		7900 => '1',
		7901 => '0',
		7902 => '1',
		7903 => '0',
		7904 => '1',
		7905 => '0',
		7906 => '1',
		7907 => '0',
		7908 => '1',
		7909 => '0',
		7910 => '1',
		7911 => '0',
		7912 => '1',
		7913 => '0',
		7914 => '1',
		7915 => '0',
		7916 => '1',
		7917 => '0',
		7918 => '1',
		7919 => '0',
		7920 => '1',
		7921 => '0',
		7922 => '1',
		7923 => '0',
		7924 => '1',
		7925 => '0',
		7926 => '1',
		7927 => '0',
		7936 => '0',
		7937 => '1',
		7938 => '0',
		7939 => '1',
		7940 => '0',
		7941 => '1',
		7942 => '0',
		7943 => '1',
		7944 => '0',
		7945 => '1',
		7946 => '0',
		7947 => '1',
		7948 => '0',
		7949 => '1',
		7950 => '0',
		7951 => '1',
		7952 => '0',
		7953 => '1',
		7954 => '0',
		7955 => '1',
		7956 => '0',
		7957 => '1',
		7958 => '0',
		7959 => '1',
		7960 => '0',
		7961 => '1',
		7962 => '0',
		7963 => '1',
		7964 => '0',
		7965 => '1',
		7966 => '0',
		7967 => '1',
		7968 => '0',
		7969 => '1',
		7970 => '0',
		7971 => '1',
		7972 => '0',
		7973 => '1',
		7974 => '0',
		7975 => '1',
		7976 => '0',
		7977 => '1',
		7978 => '0',
		7979 => '1',
		7980 => '0',
		7981 => '1',
		7982 => '0',
		7983 => '1',
		7984 => '0',
		7985 => '1',
		7986 => '0',
		7987 => '1',
		7988 => '0',
		7989 => '1',
		7990 => '0',
		7991 => '1',
		7992 => '0',
		7993 => '1',
		7994 => '0',
		7995 => '1',
		7996 => '0',
		7997 => '1',
		7998 => '0',
		7999 => '1',
		8000 => '0',
		8001 => '1',
		8002 => '0',
		8003 => '1',
		8004 => '0',
		8005 => '1',
		8006 => '0',
		8007 => '1',
		8008 => '0',
		8009 => '1',
		8010 => '0',
		8011 => '1',
		8012 => '0',
		8013 => '1',
		8014 => '0',
		8015 => '1',
		8016 => '0',
		8017 => '1',
		8018 => '0',
		8019 => '1',
		8020 => '0',
		8021 => '1',
		8022 => '0',
		8023 => '1',
		8024 => '0',
		8025 => '1',
		8026 => '0',
		8027 => '1',
		8028 => '0',
		8029 => '1',
		8030 => '0',
		8031 => '1',
		8032 => '0',
		8033 => '1',
		8034 => '0',
		8035 => '1',
		8036 => '0',
		8037 => '1',
		8038 => '0',
		8039 => '1',
		8040 => '0',
		8041 => '1',
		8042 => '0',
		8043 => '1',
		8044 => '0',
		8045 => '1',
		8046 => '0',
		8047 => '1',
		8048 => '0',
		8049 => '1',
		8050 => '0',
		8051 => '1',
		8052 => '0',
		8053 => '1',
		8054 => '0',
		8055 => '1',
		8064 => '1',
		8065 => '0',
		8066 => '1',
		8067 => '0',
		8068 => '1',
		8069 => '0',
		8070 => '1',
		8071 => '0',
		8072 => '1',
		8073 => '0',
		8074 => '1',
		8075 => '0',
		8076 => '1',
		8077 => '0',
		8078 => '1',
		8079 => '0',
		8080 => '1',
		8081 => '0',
		8082 => '1',
		8083 => '0',
		8084 => '1',
		8085 => '0',
		8086 => '1',
		8087 => '0',
		8088 => '1',
		8089 => '0',
		8090 => '1',
		8091 => '0',
		8092 => '1',
		8093 => '0',
		8094 => '1',
		8095 => '0',
		8096 => '1',
		8097 => '0',
		8098 => '1',
		8099 => '0',
		8100 => '1',
		8101 => '0',
		8102 => '1',
		8103 => '0',
		8104 => '1',
		8105 => '0',
		8106 => '1',
		8107 => '0',
		8108 => '1',
		8109 => '0',
		8110 => '1',
		8111 => '0',
		8112 => '1',
		8113 => '0',
		8114 => '1',
		8115 => '0',
		8116 => '1',
		8117 => '0',
		8118 => '1',
		8119 => '0',
		8120 => '1',
		8121 => '0',
		8122 => '1',
		8123 => '0',
		8124 => '1',
		8125 => '0',
		8126 => '1',
		8127 => '0',
		8128 => '1',
		8129 => '0',
		8130 => '1',
		8131 => '0',
		8132 => '1',
		8133 => '0',
		8134 => '1',
		8135 => '0',
		8136 => '1',
		8137 => '0',
		8138 => '1',
		8139 => '0',
		8140 => '1',
		8141 => '0',
		8142 => '1',
		8143 => '0',
		8144 => '1',
		8145 => '0',
		8146 => '1',
		8147 => '0',
		8148 => '1',
		8149 => '0',
		8150 => '1',
		8151 => '0',
		8152 => '1',
		8153 => '0',
		8154 => '1',
		8155 => '0',
		8156 => '1',
		8157 => '0',
		8158 => '1',
		8159 => '0',
		8160 => '1',
		8161 => '0',
		8162 => '1',
		8163 => '0',
		8164 => '1',
		8165 => '0',
		8166 => '1',
		8167 => '0',
		8168 => '1',
		8169 => '0',
		8170 => '1',
		8171 => '0',
		8172 => '1',
		8173 => '0',
		8174 => '1',
		8175 => '0',
		8176 => '1',
		8177 => '0',
		8178 => '1',
		8179 => '0',
		8180 => '1',
		8181 => '0',
		8182 => '1',
		8183 => '0',
		8192 => '0',
		8193 => '1',
		8194 => '0',
		8195 => '1',
		8196 => '0',
		8197 => '1',
		8198 => '0',
		8199 => '1',
		8200 => '0',
		8201 => '1',
		8202 => '0',
		8203 => '1',
		8204 => '0',
		8205 => '1',
		8206 => '0',
		8207 => '1',
		8208 => '0',
		8209 => '1',
		8210 => '0',
		8211 => '1',
		8212 => '0',
		8213 => '1',
		8214 => '0',
		8215 => '1',
		8216 => '0',
		8217 => '1',
		8218 => '0',
		8219 => '1',
		8220 => '0',
		8221 => '1',
		8222 => '0',
		8223 => '1',
		8224 => '0',
		8225 => '1',
		8226 => '0',
		8227 => '1',
		8228 => '0',
		8229 => '1',
		8230 => '0',
		8231 => '1',
		8232 => '0',
		8233 => '1',
		8234 => '0',
		8235 => '1',
		8236 => '0',
		8237 => '1',
		8238 => '0',
		8239 => '1',
		8240 => '0',
		8241 => '1',
		8242 => '0',
		8243 => '1',
		8244 => '0',
		8245 => '1',
		8246 => '0',
		8247 => '1',
		8248 => '0',
		8249 => '1',
		8250 => '0',
		8251 => '1',
		8252 => '0',
		8253 => '1',
		8254 => '0',
		8255 => '1',
		8256 => '0',
		8257 => '1',
		8258 => '0',
		8259 => '1',
		8260 => '0',
		8261 => '1',
		8262 => '0',
		8263 => '1',
		8264 => '0',
		8265 => '1',
		8266 => '0',
		8267 => '1',
		8268 => '0',
		8269 => '1',
		8270 => '0',
		8271 => '1',
		8272 => '0',
		8273 => '1',
		8274 => '0',
		8275 => '1',
		8276 => '0',
		8277 => '1',
		8278 => '0',
		8279 => '1',
		8280 => '0',
		8281 => '1',
		8282 => '0',
		8283 => '1',
		8284 => '0',
		8285 => '1',
		8286 => '0',
		8287 => '1',
		8288 => '0',
		8289 => '1',
		8290 => '0',
		8291 => '1',
		8292 => '0',
		8293 => '1',
		8294 => '0',
		8295 => '1',
		8296 => '0',
		8297 => '1',
		8298 => '0',
		8299 => '1',
		8300 => '0',
		8301 => '1',
		8302 => '0',
		8303 => '1',
		8304 => '0',
		8305 => '1',
		8306 => '0',
		8307 => '1',
		8308 => '0',
		8309 => '1',
		8310 => '0',
		8311 => '1',
		8320 => '1',
		8321 => '0',
		8322 => '1',
		8323 => '0',
		8324 => '1',
		8325 => '0',
		8326 => '1',
		8327 => '0',
		8328 => '1',
		8329 => '0',
		8330 => '1',
		8331 => '0',
		8332 => '1',
		8333 => '0',
		8334 => '1',
		8335 => '0',
		8336 => '1',
		8337 => '0',
		8338 => '1',
		8339 => '0',
		8340 => '1',
		8341 => '0',
		8342 => '1',
		8343 => '0',
		8344 => '1',
		8345 => '0',
		8346 => '1',
		8347 => '0',
		8348 => '1',
		8349 => '0',
		8350 => '1',
		8351 => '0',
		8352 => '1',
		8353 => '0',
		8354 => '1',
		8355 => '0',
		8356 => '1',
		8357 => '0',
		8358 => '1',
		8359 => '0',
		8360 => '1',
		8361 => '0',
		8362 => '1',
		8363 => '0',
		8364 => '1',
		8365 => '0',
		8366 => '1',
		8367 => '0',
		8368 => '1',
		8369 => '0',
		8370 => '1',
		8371 => '0',
		8372 => '1',
		8373 => '0',
		8374 => '1',
		8375 => '0',
		8376 => '1',
		8377 => '0',
		8378 => '1',
		8379 => '0',
		8380 => '1',
		8381 => '0',
		8382 => '1',
		8383 => '0',
		8384 => '1',
		8385 => '0',
		8386 => '1',
		8387 => '0',
		8388 => '1',
		8389 => '0',
		8390 => '1',
		8391 => '0',
		8392 => '1',
		8393 => '0',
		8394 => '1',
		8395 => '0',
		8396 => '1',
		8397 => '0',
		8398 => '1',
		8399 => '0',
		8400 => '1',
		8401 => '0',
		8402 => '1',
		8403 => '0',
		8404 => '1',
		8405 => '0',
		8406 => '1',
		8407 => '0',
		8408 => '1',
		8409 => '0',
		8410 => '1',
		8411 => '0',
		8412 => '1',
		8413 => '0',
		8414 => '1',
		8415 => '0',
		8416 => '1',
		8417 => '0',
		8418 => '1',
		8419 => '0',
		8420 => '1',
		8421 => '0',
		8422 => '1',
		8423 => '0',
		8424 => '1',
		8425 => '0',
		8426 => '1',
		8427 => '0',
		8428 => '1',
		8429 => '0',
		8430 => '1',
		8431 => '0',
		8432 => '1',
		8433 => '0',
		8434 => '1',
		8435 => '0',
		8436 => '1',
		8437 => '0',
		8438 => '1',
		8439 => '0',
		8448 => '0',
		8449 => '1',
		8450 => '0',
		8451 => '1',
		8452 => '0',
		8453 => '1',
		8454 => '0',
		8455 => '1',
		8456 => '0',
		8457 => '1',
		8458 => '0',
		8459 => '1',
		8460 => '0',
		8461 => '1',
		8462 => '0',
		8463 => '1',
		8464 => '0',
		8465 => '1',
		8466 => '0',
		8467 => '1',
		8468 => '0',
		8469 => '1',
		8470 => '0',
		8471 => '1',
		8472 => '0',
		8473 => '1',
		8474 => '0',
		8475 => '1',
		8476 => '0',
		8477 => '1',
		8478 => '0',
		8479 => '1',
		8480 => '0',
		8481 => '1',
		8482 => '0',
		8483 => '1',
		8484 => '0',
		8485 => '1',
		8486 => '0',
		8487 => '1',
		8488 => '0',
		8489 => '1',
		8490 => '0',
		8491 => '1',
		8492 => '0',
		8493 => '1',
		8494 => '0',
		8495 => '1',
		8496 => '0',
		8497 => '1',
		8498 => '0',
		8499 => '1',
		8500 => '0',
		8501 => '1',
		8502 => '0',
		8503 => '1',
		8504 => '0',
		8505 => '1',
		8506 => '0',
		8507 => '1',
		8508 => '0',
		8509 => '1',
		8510 => '0',
		8511 => '1',
		8512 => '0',
		8513 => '1',
		8514 => '0',
		8515 => '1',
		8516 => '0',
		8517 => '1',
		8518 => '0',
		8519 => '1',
		8520 => '0',
		8521 => '1',
		8522 => '0',
		8523 => '1',
		8524 => '0',
		8525 => '1',
		8526 => '0',
		8527 => '1',
		8528 => '0',
		8529 => '1',
		8530 => '0',
		8531 => '1',
		8532 => '0',
		8533 => '1',
		8534 => '0',
		8535 => '1',
		8536 => '0',
		8537 => '1',
		8538 => '0',
		8539 => '1',
		8540 => '0',
		8541 => '1',
		8542 => '0',
		8543 => '1',
		8544 => '0',
		8545 => '1',
		8546 => '0',
		8547 => '1',
		8548 => '0',
		8549 => '1',
		8550 => '0',
		8551 => '1',
		8552 => '0',
		8553 => '1',
		8554 => '0',
		8555 => '1',
		8556 => '0',
		8557 => '1',
		8558 => '0',
		8559 => '1',
		8560 => '0',
		8561 => '1',
		8562 => '0',
		8563 => '1',
		8564 => '0',
		8565 => '1',
		8566 => '0',
		8567 => '1',
		8576 => '1',
		8577 => '0',
		8578 => '1',
		8579 => '0',
		8580 => '1',
		8581 => '0',
		8582 => '1',
		8583 => '0',
		8584 => '1',
		8585 => '0',
		8586 => '1',
		8587 => '0',
		8588 => '1',
		8589 => '0',
		8590 => '1',
		8591 => '0',
		8592 => '1',
		8593 => '0',
		8594 => '1',
		8595 => '0',
		8596 => '1',
		8597 => '0',
		8598 => '1',
		8599 => '0',
		8600 => '1',
		8601 => '0',
		8602 => '1',
		8603 => '0',
		8604 => '1',
		8605 => '0',
		8606 => '1',
		8607 => '0',
		8608 => '1',
		8609 => '0',
		8610 => '1',
		8611 => '0',
		8612 => '1',
		8613 => '0',
		8614 => '1',
		8615 => '0',
		8616 => '1',
		8617 => '0',
		8618 => '1',
		8619 => '0',
		8620 => '1',
		8621 => '0',
		8622 => '1',
		8623 => '0',
		8624 => '1',
		8625 => '0',
		8626 => '1',
		8627 => '0',
		8628 => '1',
		8629 => '0',
		8630 => '1',
		8631 => '0',
		8632 => '1',
		8633 => '0',
		8634 => '1',
		8635 => '0',
		8636 => '1',
		8637 => '0',
		8638 => '1',
		8639 => '0',
		8640 => '1',
		8641 => '0',
		8642 => '1',
		8643 => '0',
		8644 => '1',
		8645 => '0',
		8646 => '1',
		8647 => '0',
		8648 => '1',
		8649 => '0',
		8650 => '1',
		8651 => '0',
		8652 => '1',
		8653 => '0',
		8654 => '1',
		8655 => '0',
		8656 => '1',
		8657 => '0',
		8658 => '1',
		8659 => '0',
		8660 => '1',
		8661 => '0',
		8662 => '1',
		8663 => '0',
		8664 => '1',
		8665 => '0',
		8666 => '1',
		8667 => '0',
		8668 => '1',
		8669 => '0',
		8670 => '1',
		8671 => '0',
		8672 => '1',
		8673 => '0',
		8674 => '1',
		8675 => '0',
		8676 => '1',
		8677 => '0',
		8678 => '1',
		8679 => '0',
		8680 => '1',
		8681 => '0',
		8682 => '1',
		8683 => '0',
		8684 => '1',
		8685 => '0',
		8686 => '1',
		8687 => '0',
		8688 => '1',
		8689 => '0',
		8690 => '1',
		8691 => '0',
		8692 => '1',
		8693 => '0',
		8694 => '1',
		8695 => '0',
		8704 => '0',
		8705 => '1',
		8706 => '0',
		8707 => '1',
		8708 => '0',
		8709 => '1',
		8710 => '0',
		8711 => '1',
		8712 => '0',
		8713 => '1',
		8714 => '0',
		8715 => '1',
		8716 => '0',
		8717 => '1',
		8718 => '0',
		8719 => '1',
		8720 => '0',
		8721 => '1',
		8722 => '0',
		8723 => '1',
		8724 => '0',
		8725 => '1',
		8726 => '0',
		8727 => '1',
		8728 => '0',
		8729 => '1',
		8730 => '0',
		8731 => '1',
		8732 => '0',
		8733 => '1',
		8734 => '0',
		8735 => '1',
		8736 => '0',
		8737 => '1',
		8738 => '0',
		8739 => '1',
		8740 => '0',
		8741 => '1',
		8742 => '0',
		8743 => '1',
		8744 => '0',
		8745 => '1',
		8746 => '0',
		8747 => '1',
		8748 => '0',
		8749 => '1',
		8750 => '0',
		8751 => '1',
		8752 => '0',
		8753 => '1',
		8754 => '0',
		8755 => '1',
		8756 => '0',
		8757 => '1',
		8758 => '0',
		8759 => '1',
		8760 => '0',
		8761 => '1',
		8762 => '0',
		8763 => '1',
		8764 => '0',
		8765 => '1',
		8766 => '0',
		8767 => '1',
		8768 => '0',
		8769 => '1',
		8770 => '0',
		8771 => '1',
		8772 => '0',
		8773 => '1',
		8774 => '0',
		8775 => '1',
		8776 => '0',
		8777 => '1',
		8778 => '0',
		8779 => '1',
		8780 => '0',
		8781 => '1',
		8782 => '0',
		8783 => '1',
		8784 => '0',
		8785 => '1',
		8786 => '0',
		8787 => '1',
		8788 => '0',
		8789 => '1',
		8790 => '0',
		8791 => '1',
		8792 => '0',
		8793 => '1',
		8794 => '0',
		8795 => '1',
		8796 => '0',
		8797 => '1',
		8798 => '0',
		8799 => '1',
		8800 => '0',
		8801 => '1',
		8802 => '0',
		8803 => '1',
		8804 => '0',
		8805 => '1',
		8806 => '0',
		8807 => '1',
		8808 => '0',
		8809 => '1',
		8810 => '0',
		8811 => '1',
		8812 => '0',
		8813 => '1',
		8814 => '0',
		8815 => '1',
		8816 => '0',
		8817 => '1',
		8818 => '0',
		8819 => '1',
		8820 => '0',
		8821 => '1',
		8822 => '0',
		8823 => '1',
		8832 => '1',
		8833 => '0',
		8834 => '1',
		8835 => '0',
		8836 => '1',
		8837 => '0',
		8838 => '1',
		8839 => '0',
		8840 => '1',
		8841 => '0',
		8842 => '1',
		8843 => '0',
		8844 => '1',
		8845 => '0',
		8846 => '1',
		8847 => '0',
		8848 => '1',
		8849 => '0',
		8850 => '1',
		8851 => '0',
		8852 => '1',
		8853 => '0',
		8854 => '1',
		8855 => '0',
		8856 => '1',
		8857 => '0',
		8858 => '1',
		8859 => '0',
		8860 => '1',
		8861 => '0',
		8862 => '1',
		8863 => '0',
		8864 => '1',
		8865 => '0',
		8866 => '1',
		8867 => '0',
		8868 => '1',
		8869 => '0',
		8870 => '1',
		8871 => '0',
		8872 => '1',
		8873 => '0',
		8874 => '1',
		8875 => '0',
		8876 => '1',
		8877 => '0',
		8878 => '1',
		8879 => '0',
		8880 => '1',
		8881 => '0',
		8882 => '1',
		8883 => '0',
		8884 => '1',
		8885 => '0',
		8886 => '1',
		8887 => '0',
		8888 => '1',
		8889 => '0',
		8890 => '1',
		8891 => '0',
		8892 => '1',
		8893 => '0',
		8894 => '1',
		8895 => '0',
		8896 => '1',
		8897 => '0',
		8898 => '1',
		8899 => '0',
		8900 => '1',
		8901 => '0',
		8902 => '1',
		8903 => '0',
		8904 => '1',
		8905 => '0',
		8906 => '1',
		8907 => '0',
		8908 => '1',
		8909 => '0',
		8910 => '1',
		8911 => '0',
		8912 => '1',
		8913 => '0',
		8914 => '1',
		8915 => '0',
		8916 => '1',
		8917 => '0',
		8918 => '1',
		8919 => '0',
		8920 => '1',
		8921 => '0',
		8922 => '1',
		8923 => '0',
		8924 => '1',
		8925 => '0',
		8926 => '1',
		8927 => '0',
		8928 => '1',
		8929 => '0',
		8930 => '1',
		8931 => '0',
		8932 => '1',
		8933 => '0',
		8934 => '1',
		8935 => '0',
		8936 => '1',
		8937 => '0',
		8938 => '1',
		8939 => '0',
		8940 => '1',
		8941 => '0',
		8942 => '1',
		8943 => '0',
		8944 => '1',
		8945 => '0',
		8946 => '1',
		8947 => '0',
		8948 => '1',
		8949 => '0',
		8950 => '1',
		8951 => '0',
		8960 => '0',
		8961 => '1',
		8962 => '0',
		8963 => '1',
		8964 => '0',
		8965 => '1',
		8966 => '0',
		8967 => '1',
		8968 => '0',
		8969 => '1',
		8970 => '0',
		8971 => '1',
		8972 => '0',
		8973 => '1',
		8974 => '0',
		8975 => '1',
		8976 => '0',
		8977 => '1',
		8978 => '0',
		8979 => '1',
		8980 => '0',
		8981 => '1',
		8982 => '0',
		8983 => '1',
		8984 => '0',
		8985 => '1',
		8986 => '0',
		8987 => '1',
		8988 => '0',
		8989 => '1',
		8990 => '0',
		8991 => '1',
		8992 => '0',
		8993 => '1',
		8994 => '0',
		8995 => '1',
		8996 => '0',
		8997 => '1',
		8998 => '0',
		8999 => '1',
		9000 => '0',
		9001 => '1',
		9002 => '0',
		9003 => '1',
		9004 => '0',
		9005 => '1',
		9006 => '0',
		9007 => '1',
		9008 => '0',
		9009 => '1',
		9010 => '0',
		9011 => '1',
		9012 => '0',
		9013 => '1',
		9014 => '0',
		9015 => '1',
		9016 => '0',
		9017 => '1',
		9018 => '0',
		9019 => '1',
		9020 => '0',
		9021 => '1',
		9022 => '0',
		9023 => '1',
		9024 => '0',
		9025 => '1',
		9026 => '0',
		9027 => '1',
		9028 => '0',
		9029 => '1',
		9030 => '0',
		9031 => '1',
		9032 => '0',
		9033 => '1',
		9034 => '0',
		9035 => '1',
		9036 => '0',
		9037 => '1',
		9038 => '0',
		9039 => '1',
		9040 => '0',
		9041 => '1',
		9042 => '0',
		9043 => '1',
		9044 => '0',
		9045 => '1',
		9046 => '0',
		9047 => '1',
		9048 => '0',
		9049 => '1',
		9050 => '0',
		9051 => '1',
		9052 => '0',
		9053 => '1',
		9054 => '0',
		9055 => '1',
		9056 => '0',
		9057 => '1',
		9058 => '0',
		9059 => '1',
		9060 => '0',
		9061 => '1',
		9062 => '0',
		9063 => '1',
		9064 => '0',
		9065 => '1',
		9066 => '0',
		9067 => '1',
		9068 => '0',
		9069 => '1',
		9070 => '0',
		9071 => '1',
		9072 => '0',
		9073 => '1',
		9074 => '0',
		9075 => '1',
		9076 => '0',
		9077 => '1',
		9078 => '0',
		9079 => '1',
		9088 => '1',
		9089 => '0',
		9090 => '1',
		9091 => '0',
		9092 => '1',
		9093 => '0',
		9094 => '1',
		9095 => '0',
		9096 => '1',
		9097 => '0',
		9098 => '1',
		9099 => '0',
		9100 => '1',
		9101 => '0',
		9102 => '1',
		9103 => '0',
		9104 => '1',
		9105 => '0',
		9106 => '1',
		9107 => '0',
		9108 => '1',
		9109 => '0',
		9110 => '1',
		9111 => '0',
		9112 => '1',
		9113 => '0',
		9114 => '1',
		9115 => '0',
		9116 => '1',
		9117 => '0',
		9118 => '1',
		9119 => '0',
		9120 => '1',
		9121 => '0',
		9122 => '1',
		9123 => '0',
		9124 => '1',
		9125 => '0',
		9126 => '1',
		9127 => '0',
		9128 => '1',
		9129 => '0',
		9130 => '1',
		9131 => '0',
		9132 => '1',
		9133 => '0',
		9134 => '1',
		9135 => '0',
		9136 => '1',
		9137 => '0',
		9138 => '1',
		9139 => '0',
		9140 => '1',
		9141 => '0',
		9142 => '1',
		9143 => '0',
		9144 => '1',
		9145 => '0',
		9146 => '1',
		9147 => '0',
		9148 => '1',
		9149 => '0',
		9150 => '1',
		9151 => '0',
		9152 => '1',
		9153 => '0',
		9154 => '1',
		9155 => '0',
		9156 => '1',
		9157 => '0',
		9158 => '1',
		9159 => '0',
		9160 => '1',
		9161 => '0',
		9162 => '1',
		9163 => '0',
		9164 => '1',
		9165 => '0',
		9166 => '1',
		9167 => '0',
		9168 => '1',
		9169 => '0',
		9170 => '1',
		9171 => '0',
		9172 => '1',
		9173 => '0',
		9174 => '1',
		9175 => '0',
		9176 => '1',
		9177 => '0',
		9178 => '1',
		9179 => '0',
		9180 => '1',
		9181 => '0',
		9182 => '1',
		9183 => '0',
		9184 => '1',
		9185 => '0',
		9186 => '1',
		9187 => '0',
		9188 => '1',
		9189 => '0',
		9190 => '1',
		9191 => '0',
		9192 => '1',
		9193 => '0',
		9194 => '1',
		9195 => '0',
		9196 => '1',
		9197 => '0',
		9198 => '1',
		9199 => '0',
		9200 => '1',
		9201 => '0',
		9202 => '1',
		9203 => '0',
		9204 => '1',
		9205 => '0',
		9206 => '1',
		9207 => '0',
		9216 => '0',
		9217 => '1',
		9218 => '0',
		9219 => '1',
		9220 => '0',
		9221 => '1',
		9222 => '0',
		9223 => '1',
		9224 => '0',
		9225 => '1',
		9226 => '0',
		9227 => '1',
		9228 => '0',
		9229 => '1',
		9230 => '0',
		9231 => '1',
		9232 => '0',
		9233 => '1',
		9234 => '0',
		9235 => '1',
		9236 => '0',
		9237 => '1',
		9238 => '0',
		9239 => '1',
		9240 => '0',
		9241 => '1',
		9242 => '0',
		9243 => '1',
		9244 => '0',
		9245 => '1',
		9246 => '0',
		9247 => '1',
		9248 => '0',
		9249 => '1',
		9250 => '0',
		9251 => '1',
		9252 => '0',
		9253 => '1',
		9254 => '0',
		9255 => '1',
		9256 => '0',
		9257 => '1',
		9258 => '0',
		9259 => '1',
		9260 => '0',
		9261 => '1',
		9262 => '0',
		9263 => '1',
		9264 => '0',
		9265 => '1',
		9266 => '0',
		9267 => '1',
		9268 => '0',
		9269 => '1',
		9270 => '0',
		9271 => '1',
		9272 => '0',
		9273 => '1',
		9274 => '0',
		9275 => '1',
		9276 => '0',
		9277 => '1',
		9278 => '0',
		9279 => '1',
		9280 => '0',
		9281 => '1',
		9282 => '0',
		9283 => '1',
		9284 => '0',
		9285 => '1',
		9286 => '0',
		9287 => '1',
		9288 => '0',
		9289 => '1',
		9290 => '0',
		9291 => '1',
		9292 => '0',
		9293 => '1',
		9294 => '0',
		9295 => '1',
		9296 => '0',
		9297 => '1',
		9298 => '0',
		9299 => '1',
		9300 => '0',
		9301 => '1',
		9302 => '0',
		9303 => '1',
		9304 => '0',
		9305 => '1',
		9306 => '0',
		9307 => '1',
		9308 => '0',
		9309 => '1',
		9310 => '0',
		9311 => '1',
		9312 => '0',
		9313 => '1',
		9314 => '0',
		9315 => '1',
		9316 => '0',
		9317 => '1',
		9318 => '0',
		9319 => '1',
		9320 => '0',
		9321 => '1',
		9322 => '0',
		9323 => '1',
		9324 => '0',
		9325 => '1',
		9326 => '0',
		9327 => '1',
		9328 => '0',
		9329 => '1',
		9330 => '0',
		9331 => '1',
		9332 => '0',
		9333 => '1',
		9334 => '0',
		9335 => '1',
		9344 => '1',
		9345 => '0',
		9346 => '1',
		9347 => '0',
		9348 => '1',
		9349 => '0',
		9350 => '1',
		9351 => '0',
		9352 => '1',
		9353 => '0',
		9354 => '1',
		9355 => '0',
		9356 => '1',
		9357 => '0',
		9358 => '1',
		9359 => '0',
		9360 => '1',
		9361 => '0',
		9362 => '1',
		9363 => '0',
		9364 => '1',
		9365 => '0',
		9366 => '1',
		9367 => '0',
		9368 => '1',
		9369 => '0',
		9370 => '1',
		9371 => '0',
		9372 => '1',
		9373 => '0',
		9374 => '1',
		9375 => '0',
		9376 => '1',
		9377 => '0',
		9378 => '1',
		9379 => '0',
		9380 => '1',
		9381 => '0',
		9382 => '1',
		9383 => '0',
		9384 => '1',
		9385 => '0',
		9386 => '1',
		9387 => '0',
		9388 => '1',
		9389 => '0',
		9390 => '1',
		9391 => '0',
		9392 => '1',
		9393 => '0',
		9394 => '1',
		9395 => '0',
		9396 => '1',
		9397 => '0',
		9398 => '1',
		9399 => '0',
		9400 => '1',
		9401 => '0',
		9402 => '1',
		9403 => '0',
		9404 => '1',
		9405 => '0',
		9406 => '1',
		9407 => '0',
		9408 => '1',
		9409 => '0',
		9410 => '1',
		9411 => '0',
		9412 => '1',
		9413 => '0',
		9414 => '1',
		9415 => '0',
		9416 => '1',
		9417 => '0',
		9418 => '1',
		9419 => '0',
		9420 => '1',
		9421 => '0',
		9422 => '1',
		9423 => '0',
		9424 => '1',
		9425 => '0',
		9426 => '1',
		9427 => '0',
		9428 => '1',
		9429 => '0',
		9430 => '1',
		9431 => '0',
		9432 => '1',
		9433 => '0',
		9434 => '1',
		9435 => '0',
		9436 => '1',
		9437 => '0',
		9438 => '1',
		9439 => '0',
		9440 => '1',
		9441 => '0',
		9442 => '1',
		9443 => '0',
		9444 => '1',
		9445 => '0',
		9446 => '1',
		9447 => '0',
		9448 => '1',
		9449 => '0',
		9450 => '1',
		9451 => '0',
		9452 => '1',
		9453 => '0',
		9454 => '1',
		9455 => '0',
		9456 => '1',
		9457 => '0',
		9458 => '1',
		9459 => '0',
		9460 => '1',
		9461 => '0',
		9462 => '1',
		9463 => '0',
		9472 => '0',
		9473 => '1',
		9474 => '0',
		9475 => '1',
		9476 => '0',
		9477 => '1',
		9478 => '0',
		9479 => '1',
		9480 => '0',
		9481 => '1',
		9482 => '0',
		9483 => '1',
		9484 => '0',
		9485 => '1',
		9486 => '0',
		9487 => '1',
		9488 => '0',
		9489 => '1',
		9490 => '0',
		9491 => '1',
		9492 => '0',
		9493 => '1',
		9494 => '0',
		9495 => '1',
		9496 => '0',
		9497 => '1',
		9498 => '0',
		9499 => '1',
		9500 => '0',
		9501 => '1',
		9502 => '0',
		9503 => '1',
		9504 => '0',
		9505 => '1',
		9506 => '0',
		9507 => '1',
		9508 => '0',
		9509 => '1',
		9510 => '0',
		9511 => '1',
		9512 => '0',
		9513 => '1',
		9514 => '0',
		9515 => '1',
		9516 => '0',
		9517 => '1',
		9518 => '0',
		9519 => '1',
		9520 => '0',
		9521 => '1',
		9522 => '0',
		9523 => '1',
		9524 => '0',
		9525 => '1',
		9526 => '0',
		9527 => '1',
		9528 => '0',
		9529 => '1',
		9530 => '0',
		9531 => '1',
		9532 => '0',
		9533 => '1',
		9534 => '0',
		9535 => '1',
		9536 => '0',
		9537 => '1',
		9538 => '0',
		9539 => '1',
		9540 => '0',
		9541 => '1',
		9542 => '0',
		9543 => '1',
		9544 => '0',
		9545 => '1',
		9546 => '0',
		9547 => '1',
		9548 => '0',
		9549 => '1',
		9550 => '0',
		9551 => '1',
		9552 => '0',
		9553 => '1',
		9554 => '0',
		9555 => '1',
		9556 => '0',
		9557 => '1',
		9558 => '0',
		9559 => '1',
		9560 => '0',
		9561 => '1',
		9562 => '0',
		9563 => '1',
		9564 => '0',
		9565 => '1',
		9566 => '0',
		9567 => '1',
		9568 => '0',
		9569 => '1',
		9570 => '0',
		9571 => '1',
		9572 => '0',
		9573 => '1',
		9574 => '0',
		9575 => '1',
		9576 => '0',
		9577 => '1',
		9578 => '0',
		9579 => '1',
		9580 => '0',
		9581 => '1',
		9582 => '0',
		9583 => '1',
		9584 => '0',
		9585 => '1',
		9586 => '0',
		9587 => '1',
		9588 => '0',
		9589 => '1',
		9590 => '0',
		9591 => '1',
		9600 => '1',
		9601 => '0',
		9602 => '1',
		9603 => '0',
		9604 => '1',
		9605 => '0',
		9606 => '1',
		9607 => '0',
		9608 => '1',
		9609 => '0',
		9610 => '1',
		9611 => '0',
		9612 => '1',
		9613 => '0',
		9614 => '1',
		9615 => '0',
		9616 => '1',
		9617 => '0',
		9618 => '1',
		9619 => '0',
		9620 => '1',
		9621 => '0',
		9622 => '1',
		9623 => '0',
		9624 => '1',
		9625 => '0',
		9626 => '1',
		9627 => '0',
		9628 => '1',
		9629 => '0',
		9630 => '1',
		9631 => '0',
		9632 => '1',
		9633 => '0',
		9634 => '1',
		9635 => '0',
		9636 => '1',
		9637 => '0',
		9638 => '1',
		9639 => '0',
		9640 => '1',
		9641 => '0',
		9642 => '1',
		9643 => '0',
		9644 => '1',
		9645 => '0',
		9646 => '1',
		9647 => '0',
		9648 => '1',
		9649 => '0',
		9650 => '1',
		9651 => '0',
		9652 => '1',
		9653 => '0',
		9654 => '1',
		9655 => '0',
		9656 => '1',
		9657 => '0',
		9658 => '1',
		9659 => '0',
		9660 => '1',
		9661 => '0',
		9662 => '1',
		9663 => '0',
		9664 => '1',
		9665 => '0',
		9666 => '1',
		9667 => '0',
		9668 => '1',
		9669 => '0',
		9670 => '1',
		9671 => '0',
		9672 => '1',
		9673 => '0',
		9674 => '1',
		9675 => '0',
		9676 => '1',
		9677 => '0',
		9678 => '1',
		9679 => '0',
		9680 => '1',
		9681 => '0',
		9682 => '1',
		9683 => '0',
		9684 => '1',
		9685 => '0',
		9686 => '1',
		9687 => '0',
		9688 => '1',
		9689 => '0',
		9690 => '1',
		9691 => '0',
		9692 => '1',
		9693 => '0',
		9694 => '1',
		9695 => '0',
		9696 => '1',
		9697 => '0',
		9698 => '1',
		9699 => '0',
		9700 => '1',
		9701 => '0',
		9702 => '1',
		9703 => '0',
		9704 => '1',
		9705 => '0',
		9706 => '1',
		9707 => '0',
		9708 => '1',
		9709 => '0',
		9710 => '1',
		9711 => '0',
		9712 => '1',
		9713 => '0',
		9714 => '1',
		9715 => '0',
		9716 => '1',
		9717 => '0',
		9718 => '1',
		9719 => '0',
		9728 => '0',
		9729 => '1',
		9730 => '0',
		9731 => '1',
		9732 => '0',
		9733 => '1',
		9734 => '0',
		9735 => '1',
		9736 => '0',
		9737 => '1',
		9738 => '0',
		9739 => '1',
		9740 => '0',
		9741 => '1',
		9742 => '0',
		9743 => '1',
		9744 => '0',
		9745 => '1',
		9746 => '0',
		9747 => '1',
		9748 => '0',
		9749 => '1',
		9750 => '0',
		9751 => '1',
		9752 => '0',
		9753 => '1',
		9754 => '0',
		9755 => '1',
		9756 => '0',
		9757 => '1',
		9758 => '0',
		9759 => '1',
		9760 => '0',
		9761 => '1',
		9762 => '0',
		9763 => '1',
		9764 => '0',
		9765 => '1',
		9766 => '0',
		9767 => '1',
		9768 => '0',
		9769 => '1',
		9770 => '0',
		9771 => '1',
		9772 => '0',
		9773 => '1',
		9774 => '0',
		9775 => '1',
		9776 => '0',
		9777 => '1',
		9778 => '0',
		9779 => '1',
		9780 => '0',
		9781 => '1',
		9782 => '0',
		9783 => '1',
		9784 => '0',
		9785 => '1',
		9786 => '0',
		9787 => '1',
		9788 => '0',
		9789 => '1',
		9790 => '0',
		9791 => '1',
		9792 => '0',
		9793 => '1',
		9794 => '0',
		9795 => '1',
		9796 => '0',
		9797 => '1',
		9798 => '0',
		9799 => '1',
		9800 => '0',
		9801 => '1',
		9802 => '0',
		9803 => '1',
		9804 => '0',
		9805 => '1',
		9806 => '0',
		9807 => '1',
		9808 => '0',
		9809 => '1',
		9810 => '0',
		9811 => '1',
		9812 => '0',
		9813 => '1',
		9814 => '0',
		9815 => '1',
		9816 => '0',
		9817 => '1',
		9818 => '0',
		9819 => '1',
		9820 => '0',
		9821 => '1',
		9822 => '0',
		9823 => '1',
		9824 => '0',
		9825 => '1',
		9826 => '0',
		9827 => '1',
		9828 => '0',
		9829 => '1',
		9830 => '0',
		9831 => '1',
		9832 => '0',
		9833 => '1',
		9834 => '0',
		9835 => '1',
		9836 => '0',
		9837 => '1',
		9838 => '0',
		9839 => '1',
		9840 => '0',
		9841 => '1',
		9842 => '0',
		9843 => '1',
		9844 => '0',
		9845 => '1',
		9846 => '0',
		9847 => '1',
		9856 => '1',
		9857 => '0',
		9858 => '1',
		9859 => '0',
		9860 => '1',
		9861 => '0',
		9862 => '1',
		9863 => '0',
		9864 => '1',
		9865 => '0',
		9866 => '1',
		9867 => '0',
		9868 => '1',
		9869 => '0',
		9870 => '1',
		9871 => '0',
		9872 => '1',
		9873 => '0',
		9874 => '1',
		9875 => '0',
		9876 => '1',
		9877 => '0',
		9878 => '1',
		9879 => '0',
		9880 => '1',
		9881 => '0',
		9882 => '1',
		9883 => '0',
		9884 => '1',
		9885 => '0',
		9886 => '1',
		9887 => '0',
		9888 => '1',
		9889 => '0',
		9890 => '1',
		9891 => '0',
		9892 => '1',
		9893 => '0',
		9894 => '1',
		9895 => '0',
		9896 => '1',
		9897 => '0',
		9898 => '1',
		9899 => '0',
		9900 => '1',
		9901 => '0',
		9902 => '1',
		9903 => '0',
		9904 => '1',
		9905 => '0',
		9906 => '1',
		9907 => '0',
		9908 => '1',
		9909 => '0',
		9910 => '1',
		9911 => '0',
		9912 => '1',
		9913 => '0',
		9914 => '1',
		9915 => '0',
		9916 => '1',
		9917 => '0',
		9918 => '1',
		9919 => '0',
		9920 => '1',
		9921 => '0',
		9922 => '1',
		9923 => '0',
		9924 => '1',
		9925 => '0',
		9926 => '1',
		9927 => '0',
		9928 => '1',
		9929 => '0',
		9930 => '1',
		9931 => '0',
		9932 => '1',
		9933 => '0',
		9934 => '1',
		9935 => '0',
		9936 => '1',
		9937 => '0',
		9938 => '1',
		9939 => '0',
		9940 => '1',
		9941 => '0',
		9942 => '1',
		9943 => '0',
		9944 => '1',
		9945 => '0',
		9946 => '1',
		9947 => '0',
		9948 => '1',
		9949 => '0',
		9950 => '1',
		9951 => '0',
		9952 => '1',
		9953 => '0',
		9954 => '1',
		9955 => '0',
		9956 => '1',
		9957 => '0',
		9958 => '1',
		9959 => '0',
		9960 => '1',
		9961 => '0',
		9962 => '1',
		9963 => '0',
		9964 => '1',
		9965 => '0',
		9966 => '1',
		9967 => '0',
		9968 => '1',
		9969 => '0',
		9970 => '1',
		9971 => '0',
		9972 => '1',
		9973 => '0',
		9974 => '1',
		9975 => '0',
		9984 => '0',
		9985 => '1',
		9986 => '0',
		9987 => '1',
		9988 => '0',
		9989 => '1',
		9990 => '0',
		9991 => '1',
		9992 => '0',
		9993 => '1',
		9994 => '0',
		9995 => '1',
		9996 => '0',
		9997 => '1',
		9998 => '0',
		9999 => '1',
		10000 => '0',
		10001 => '1',
		10002 => '0',
		10003 => '1',
		10004 => '0',
		10005 => '1',
		10006 => '0',
		10007 => '1',
		10008 => '0',
		10009 => '1',
		10010 => '0',
		10011 => '1',
		10012 => '0',
		10013 => '1',
		10014 => '0',
		10015 => '1',
		10016 => '0',
		10017 => '1',
		10018 => '0',
		10019 => '1',
		10020 => '0',
		10021 => '1',
		10022 => '0',
		10023 => '1',
		10024 => '0',
		10025 => '1',
		10026 => '0',
		10027 => '1',
		10028 => '0',
		10029 => '1',
		10030 => '0',
		10031 => '1',
		10032 => '0',
		10033 => '1',
		10034 => '0',
		10035 => '1',
		10036 => '0',
		10037 => '1',
		10038 => '0',
		10039 => '1',
		10040 => '0',
		10041 => '1',
		10042 => '0',
		10043 => '1',
		10044 => '0',
		10045 => '1',
		10046 => '0',
		10047 => '1',
		10048 => '0',
		10049 => '1',
		10050 => '0',
		10051 => '1',
		10052 => '0',
		10053 => '1',
		10054 => '0',
		10055 => '1',
		10056 => '0',
		10057 => '1',
		10058 => '0',
		10059 => '1',
		10060 => '0',
		10061 => '1',
		10062 => '0',
		10063 => '1',
		10064 => '0',
		10065 => '1',
		10066 => '0',
		10067 => '1',
		10068 => '0',
		10069 => '1',
		10070 => '0',
		10071 => '1',
		10072 => '0',
		10073 => '1',
		10074 => '0',
		10075 => '1',
		10076 => '0',
		10077 => '1',
		10078 => '0',
		10079 => '1',
		10080 => '0',
		10081 => '1',
		10082 => '0',
		10083 => '1',
		10084 => '0',
		10085 => '1',
		10086 => '0',
		10087 => '1',
		10088 => '0',
		10089 => '1',
		10090 => '0',
		10091 => '1',
		10092 => '0',
		10093 => '1',
		10094 => '0',
		10095 => '1',
		10096 => '0',
		10097 => '1',
		10098 => '0',
		10099 => '1',
		10100 => '0',
		10101 => '1',
		10102 => '0',
		10103 => '1',
		10112 => '1',
		10113 => '0',
		10114 => '1',
		10115 => '0',
		10116 => '1',
		10117 => '0',
		10118 => '1',
		10119 => '0',
		10120 => '1',
		10121 => '0',
		10122 => '1',
		10123 => '0',
		10124 => '1',
		10125 => '0',
		10126 => '1',
		10127 => '0',
		10128 => '1',
		10129 => '0',
		10130 => '1',
		10131 => '0',
		10132 => '1',
		10133 => '0',
		10134 => '1',
		10135 => '0',
		10136 => '1',
		10137 => '0',
		10138 => '1',
		10139 => '0',
		10140 => '1',
		10141 => '0',
		10142 => '1',
		10143 => '0',
		10144 => '1',
		10145 => '0',
		10146 => '1',
		10147 => '0',
		10148 => '1',
		10149 => '0',
		10150 => '1',
		10151 => '0',
		10152 => '1',
		10153 => '0',
		10154 => '1',
		10155 => '0',
		10156 => '1',
		10157 => '0',
		10158 => '1',
		10159 => '0',
		10160 => '1',
		10161 => '0',
		10162 => '1',
		10163 => '0',
		10164 => '1',
		10165 => '0',
		10166 => '1',
		10167 => '0',
		10168 => '1',
		10169 => '0',
		10170 => '1',
		10171 => '0',
		10172 => '1',
		10173 => '0',
		10174 => '1',
		10175 => '0',
		10176 => '1',
		10177 => '0',
		10178 => '1',
		10179 => '0',
		10180 => '1',
		10181 => '0',
		10182 => '1',
		10183 => '0',
		10184 => '1',
		10185 => '0',
		10186 => '1',
		10187 => '0',
		10188 => '1',
		10189 => '0',
		10190 => '1',
		10191 => '0',
		10192 => '1',
		10193 => '0',
		10194 => '1',
		10195 => '0',
		10196 => '1',
		10197 => '0',
		10198 => '1',
		10199 => '0',
		10200 => '1',
		10201 => '0',
		10202 => '1',
		10203 => '0',
		10204 => '1',
		10205 => '0',
		10206 => '1',
		10207 => '0',
		10208 => '1',
		10209 => '0',
		10210 => '1',
		10211 => '0',
		10212 => '1',
		10213 => '0',
		10214 => '1',
		10215 => '0',
		10216 => '1',
		10217 => '0',
		10218 => '1',
		10219 => '0',
		10220 => '1',
		10221 => '0',
		10222 => '1',
		10223 => '0',
		10224 => '1',
		10225 => '0',
		10226 => '1',
		10227 => '0',
		10228 => '1',
		10229 => '0',
		10230 => '1',
		10231 => '0',
		10240 => '0',
		10241 => '1',
		10242 => '0',
		10243 => '1',
		10244 => '0',
		10245 => '1',
		10246 => '0',
		10247 => '1',
		10248 => '0',
		10249 => '1',
		10250 => '0',
		10251 => '1',
		10252 => '0',
		10253 => '1',
		10254 => '0',
		10255 => '1',
		10256 => '0',
		10257 => '1',
		10258 => '0',
		10259 => '1',
		10260 => '0',
		10261 => '1',
		10262 => '0',
		10263 => '1',
		10264 => '0',
		10265 => '1',
		10266 => '0',
		10267 => '1',
		10268 => '0',
		10269 => '1',
		10270 => '0',
		10271 => '1',
		10272 => '0',
		10273 => '1',
		10274 => '0',
		10275 => '1',
		10276 => '0',
		10277 => '1',
		10278 => '0',
		10279 => '1',
		10280 => '0',
		10281 => '1',
		10282 => '0',
		10283 => '1',
		10284 => '0',
		10285 => '1',
		10286 => '0',
		10287 => '1',
		10288 => '0',
		10289 => '1',
		10290 => '0',
		10291 => '1',
		10292 => '0',
		10293 => '1',
		10294 => '0',
		10295 => '1',
		10296 => '0',
		10297 => '1',
		10298 => '0',
		10299 => '1',
		10300 => '0',
		10301 => '1',
		10302 => '0',
		10303 => '1',
		10304 => '0',
		10305 => '1',
		10306 => '0',
		10307 => '1',
		10308 => '0',
		10309 => '1',
		10310 => '0',
		10311 => '1',
		10312 => '0',
		10313 => '1',
		10314 => '0',
		10315 => '1',
		10316 => '0',
		10317 => '1',
		10318 => '0',
		10319 => '1',
		10320 => '0',
		10321 => '1',
		10322 => '0',
		10323 => '1',
		10324 => '0',
		10325 => '1',
		10326 => '0',
		10327 => '1',
		10328 => '0',
		10329 => '1',
		10330 => '0',
		10331 => '1',
		10332 => '0',
		10333 => '1',
		10334 => '0',
		10335 => '1',
		10336 => '0',
		10337 => '1',
		10338 => '0',
		10339 => '1',
		10340 => '0',
		10341 => '1',
		10342 => '0',
		10343 => '1',
		10344 => '0',
		10345 => '1',
		10346 => '0',
		10347 => '1',
		10348 => '0',
		10349 => '1',
		10350 => '0',
		10351 => '1',
		10352 => '0',
		10353 => '1',
		10354 => '0',
		10355 => '1',
		10356 => '0',
		10357 => '1',
		10358 => '0',
		10359 => '1',
		10368 => '1',
		10369 => '0',
		10370 => '1',
		10371 => '0',
		10372 => '1',
		10373 => '0',
		10374 => '1',
		10375 => '0',
		10376 => '1',
		10377 => '0',
		10378 => '1',
		10379 => '0',
		10380 => '1',
		10381 => '0',
		10382 => '1',
		10383 => '0',
		10384 => '1',
		10385 => '0',
		10386 => '1',
		10387 => '0',
		10388 => '1',
		10389 => '0',
		10390 => '1',
		10391 => '0',
		10392 => '1',
		10393 => '0',
		10394 => '1',
		10395 => '0',
		10396 => '1',
		10397 => '0',
		10398 => '1',
		10399 => '0',
		10400 => '1',
		10401 => '0',
		10402 => '1',
		10403 => '0',
		10404 => '1',
		10405 => '0',
		10406 => '1',
		10407 => '0',
		10408 => '1',
		10409 => '0',
		10410 => '1',
		10411 => '0',
		10412 => '1',
		10413 => '0',
		10414 => '1',
		10415 => '0',
		10416 => '1',
		10417 => '0',
		10418 => '1',
		10419 => '0',
		10420 => '1',
		10421 => '0',
		10422 => '1',
		10423 => '0',
		10424 => '1',
		10425 => '0',
		10426 => '1',
		10427 => '0',
		10428 => '1',
		10429 => '0',
		10430 => '1',
		10431 => '0',
		10432 => '1',
		10433 => '0',
		10434 => '1',
		10435 => '0',
		10436 => '1',
		10437 => '0',
		10438 => '1',
		10439 => '0',
		10440 => '1',
		10441 => '0',
		10442 => '1',
		10443 => '0',
		10444 => '1',
		10445 => '0',
		10446 => '1',
		10447 => '0',
		10448 => '1',
		10449 => '0',
		10450 => '1',
		10451 => '0',
		10452 => '1',
		10453 => '0',
		10454 => '1',
		10455 => '0',
		10456 => '1',
		10457 => '0',
		10458 => '1',
		10459 => '0',
		10460 => '1',
		10461 => '0',
		10462 => '1',
		10463 => '0',
		10464 => '1',
		10465 => '0',
		10466 => '1',
		10467 => '0',
		10468 => '1',
		10469 => '0',
		10470 => '1',
		10471 => '0',
		10472 => '1',
		10473 => '0',
		10474 => '1',
		10475 => '0',
		10476 => '1',
		10477 => '0',
		10478 => '1',
		10479 => '0',
		10480 => '1',
		10481 => '0',
		10482 => '1',
		10483 => '0',
		10484 => '1',
		10485 => '0',
		10486 => '1',
		10487 => '0',
		10496 => '0',
		10497 => '1',
		10498 => '0',
		10499 => '1',
		10500 => '0',
		10501 => '1',
		10502 => '0',
		10503 => '1',
		10504 => '0',
		10505 => '1',
		10506 => '0',
		10507 => '1',
		10508 => '0',
		10509 => '1',
		10510 => '0',
		10511 => '1',
		10512 => '0',
		10513 => '1',
		10514 => '0',
		10515 => '1',
		10516 => '0',
		10517 => '1',
		10518 => '0',
		10519 => '1',
		10520 => '0',
		10521 => '1',
		10522 => '0',
		10523 => '1',
		10524 => '0',
		10525 => '1',
		10526 => '0',
		10527 => '1',
		10528 => '0',
		10529 => '1',
		10530 => '0',
		10531 => '1',
		10532 => '0',
		10533 => '1',
		10534 => '0',
		10535 => '1',
		10536 => '0',
		10537 => '1',
		10538 => '0',
		10539 => '1',
		10540 => '0',
		10541 => '1',
		10542 => '0',
		10543 => '1',
		10544 => '0',
		10545 => '1',
		10546 => '0',
		10547 => '1',
		10548 => '0',
		10549 => '1',
		10550 => '0',
		10551 => '1',
		10552 => '0',
		10553 => '1',
		10554 => '0',
		10555 => '1',
		10556 => '0',
		10557 => '1',
		10558 => '0',
		10559 => '1',
		10560 => '0',
		10561 => '1',
		10562 => '0',
		10563 => '1',
		10564 => '0',
		10565 => '1',
		10566 => '0',
		10567 => '1',
		10568 => '0',
		10569 => '1',
		10570 => '0',
		10571 => '1',
		10572 => '0',
		10573 => '1',
		10574 => '0',
		10575 => '1',
		10576 => '0',
		10577 => '1',
		10578 => '0',
		10579 => '1',
		10580 => '0',
		10581 => '1',
		10582 => '0',
		10583 => '1',
		10584 => '0',
		10585 => '1',
		10586 => '0',
		10587 => '1',
		10588 => '0',
		10589 => '1',
		10590 => '0',
		10591 => '1',
		10592 => '0',
		10593 => '1',
		10594 => '0',
		10595 => '1',
		10596 => '0',
		10597 => '1',
		10598 => '0',
		10599 => '1',
		10600 => '0',
		10601 => '1',
		10602 => '0',
		10603 => '1',
		10604 => '0',
		10605 => '1',
		10606 => '0',
		10607 => '1',
		10608 => '0',
		10609 => '1',
		10610 => '0',
		10611 => '1',
		10612 => '0',
		10613 => '1',
		10614 => '0',
		10615 => '1',
		10624 => '1',
		10625 => '0',
		10626 => '1',
		10627 => '0',
		10628 => '1',
		10629 => '0',
		10630 => '1',
		10631 => '0',
		10632 => '1',
		10633 => '0',
		10634 => '1',
		10635 => '0',
		10636 => '1',
		10637 => '0',
		10638 => '1',
		10639 => '0',
		10640 => '1',
		10641 => '0',
		10642 => '1',
		10643 => '0',
		10644 => '1',
		10645 => '0',
		10646 => '1',
		10647 => '0',
		10648 => '1',
		10649 => '0',
		10650 => '1',
		10651 => '0',
		10652 => '1',
		10653 => '0',
		10654 => '1',
		10655 => '0',
		10656 => '1',
		10657 => '0',
		10658 => '1',
		10659 => '0',
		10660 => '1',
		10661 => '0',
		10662 => '1',
		10663 => '0',
		10664 => '1',
		10665 => '0',
		10666 => '1',
		10667 => '0',
		10668 => '1',
		10669 => '0',
		10670 => '1',
		10671 => '0',
		10672 => '1',
		10673 => '0',
		10674 => '1',
		10675 => '0',
		10676 => '1',
		10677 => '0',
		10678 => '1',
		10679 => '0',
		10680 => '1',
		10681 => '0',
		10682 => '1',
		10683 => '0',
		10684 => '1',
		10685 => '0',
		10686 => '1',
		10687 => '0',
		10688 => '1',
		10689 => '0',
		10690 => '1',
		10691 => '0',
		10692 => '1',
		10693 => '0',
		10694 => '1',
		10695 => '0',
		10696 => '1',
		10697 => '0',
		10698 => '1',
		10699 => '0',
		10700 => '1',
		10701 => '0',
		10702 => '1',
		10703 => '0',
		10704 => '1',
		10705 => '0',
		10706 => '1',
		10707 => '0',
		10708 => '1',
		10709 => '0',
		10710 => '1',
		10711 => '0',
		10712 => '1',
		10713 => '0',
		10714 => '1',
		10715 => '0',
		10716 => '1',
		10717 => '0',
		10718 => '1',
		10719 => '0',
		10720 => '1',
		10721 => '0',
		10722 => '1',
		10723 => '0',
		10724 => '1',
		10725 => '0',
		10726 => '1',
		10727 => '0',
		10728 => '1',
		10729 => '0',
		10730 => '1',
		10731 => '0',
		10732 => '1',
		10733 => '0',
		10734 => '1',
		10735 => '0',
		10736 => '1',
		10737 => '0',
		10738 => '1',
		10739 => '0',
		10740 => '1',
		10741 => '0',
		10742 => '1',
		10743 => '0',
		10752 => '0',
		10753 => '1',
		10754 => '0',
		10755 => '1',
		10756 => '0',
		10757 => '1',
		10758 => '0',
		10759 => '1',
		10760 => '0',
		10761 => '1',
		10762 => '0',
		10763 => '1',
		10764 => '0',
		10765 => '1',
		10766 => '0',
		10767 => '1',
		10768 => '0',
		10769 => '1',
		10770 => '0',
		10771 => '1',
		10772 => '0',
		10773 => '1',
		10774 => '0',
		10775 => '1',
		10776 => '0',
		10777 => '1',
		10778 => '0',
		10779 => '1',
		10780 => '0',
		10781 => '1',
		10782 => '0',
		10783 => '1',
		10784 => '0',
		10785 => '1',
		10786 => '0',
		10787 => '1',
		10788 => '0',
		10789 => '1',
		10790 => '0',
		10791 => '1',
		10792 => '0',
		10793 => '1',
		10794 => '0',
		10795 => '1',
		10796 => '0',
		10797 => '1',
		10798 => '0',
		10799 => '1',
		10800 => '0',
		10801 => '1',
		10802 => '0',
		10803 => '1',
		10804 => '0',
		10805 => '1',
		10806 => '0',
		10807 => '1',
		10808 => '0',
		10809 => '1',
		10810 => '0',
		10811 => '1',
		10812 => '0',
		10813 => '1',
		10814 => '0',
		10815 => '1',
		10816 => '0',
		10817 => '1',
		10818 => '0',
		10819 => '1',
		10820 => '0',
		10821 => '1',
		10822 => '0',
		10823 => '1',
		10824 => '0',
		10825 => '1',
		10826 => '0',
		10827 => '1',
		10828 => '0',
		10829 => '1',
		10830 => '0',
		10831 => '1',
		10832 => '0',
		10833 => '1',
		10834 => '0',
		10835 => '1',
		10836 => '0',
		10837 => '1',
		10838 => '0',
		10839 => '1',
		10840 => '0',
		10841 => '1',
		10842 => '0',
		10843 => '1',
		10844 => '0',
		10845 => '1',
		10846 => '0',
		10847 => '1',
		10848 => '0',
		10849 => '1',
		10850 => '0',
		10851 => '1',
		10852 => '0',
		10853 => '1',
		10854 => '0',
		10855 => '1',
		10856 => '0',
		10857 => '1',
		10858 => '0',
		10859 => '1',
		10860 => '0',
		10861 => '1',
		10862 => '0',
		10863 => '1',
		10864 => '0',
		10865 => '1',
		10866 => '0',
		10867 => '1',
		10868 => '0',
		10869 => '1',
		10870 => '0',
		10871 => '1',
		10880 => '1',
		10881 => '0',
		10882 => '1',
		10883 => '0',
		10884 => '1',
		10885 => '0',
		10886 => '1',
		10887 => '0',
		10888 => '1',
		10889 => '0',
		10890 => '1',
		10891 => '0',
		10892 => '1',
		10893 => '0',
		10894 => '1',
		10895 => '0',
		10896 => '1',
		10897 => '0',
		10898 => '1',
		10899 => '0',
		10900 => '1',
		10901 => '0',
		10902 => '1',
		10903 => '0',
		10904 => '1',
		10905 => '0',
		10906 => '1',
		10907 => '0',
		10908 => '1',
		10909 => '0',
		10910 => '1',
		10911 => '0',
		10912 => '1',
		10913 => '0',
		10914 => '1',
		10915 => '0',
		10916 => '1',
		10917 => '0',
		10918 => '1',
		10919 => '0',
		10920 => '1',
		10921 => '0',
		10922 => '1',
		10923 => '0',
		10924 => '1',
		10925 => '0',
		10926 => '1',
		10927 => '0',
		10928 => '1',
		10929 => '0',
		10930 => '1',
		10931 => '0',
		10932 => '1',
		10933 => '0',
		10934 => '1',
		10935 => '0',
		10936 => '1',
		10937 => '0',
		10938 => '1',
		10939 => '0',
		10940 => '1',
		10941 => '0',
		10942 => '1',
		10943 => '0',
		10944 => '1',
		10945 => '0',
		10946 => '1',
		10947 => '0',
		10948 => '1',
		10949 => '0',
		10950 => '1',
		10951 => '0',
		10952 => '1',
		10953 => '0',
		10954 => '1',
		10955 => '0',
		10956 => '1',
		10957 => '0',
		10958 => '1',
		10959 => '0',
		10960 => '1',
		10961 => '0',
		10962 => '1',
		10963 => '0',
		10964 => '1',
		10965 => '0',
		10966 => '1',
		10967 => '0',
		10968 => '1',
		10969 => '0',
		10970 => '1',
		10971 => '0',
		10972 => '1',
		10973 => '0',
		10974 => '1',
		10975 => '0',
		10976 => '1',
		10977 => '0',
		10978 => '1',
		10979 => '0',
		10980 => '1',
		10981 => '0',
		10982 => '1',
		10983 => '0',
		10984 => '1',
		10985 => '0',
		10986 => '1',
		10987 => '0',
		10988 => '1',
		10989 => '0',
		10990 => '1',
		10991 => '0',
		10992 => '1',
		10993 => '0',
		10994 => '1',
		10995 => '0',
		10996 => '1',
		10997 => '0',
		10998 => '1',
		10999 => '0',
		11008 => '0',
		11009 => '1',
		11010 => '0',
		11011 => '1',
		11012 => '0',
		11013 => '1',
		11014 => '0',
		11015 => '1',
		11016 => '0',
		11017 => '1',
		11018 => '0',
		11019 => '1',
		11020 => '0',
		11021 => '1',
		11022 => '0',
		11023 => '1',
		11024 => '0',
		11025 => '1',
		11026 => '0',
		11027 => '1',
		11028 => '0',
		11029 => '1',
		11030 => '0',
		11031 => '1',
		11032 => '0',
		11033 => '1',
		11034 => '0',
		11035 => '1',
		11036 => '0',
		11037 => '1',
		11038 => '0',
		11039 => '1',
		11040 => '0',
		11041 => '1',
		11042 => '0',
		11043 => '1',
		11044 => '0',
		11045 => '1',
		11046 => '0',
		11047 => '1',
		11048 => '0',
		11049 => '1',
		11050 => '0',
		11051 => '1',
		11052 => '0',
		11053 => '1',
		11054 => '0',
		11055 => '1',
		11056 => '0',
		11057 => '1',
		11058 => '0',
		11059 => '1',
		11060 => '0',
		11061 => '1',
		11062 => '0',
		11063 => '1',
		11064 => '0',
		11065 => '1',
		11066 => '0',
		11067 => '1',
		11068 => '0',
		11069 => '1',
		11070 => '0',
		11071 => '1',
		11072 => '0',
		11073 => '1',
		11074 => '0',
		11075 => '1',
		11076 => '0',
		11077 => '1',
		11078 => '0',
		11079 => '1',
		11080 => '0',
		11081 => '1',
		11082 => '0',
		11083 => '1',
		11084 => '0',
		11085 => '1',
		11086 => '0',
		11087 => '1',
		11088 => '0',
		11089 => '1',
		11090 => '0',
		11091 => '1',
		11092 => '0',
		11093 => '1',
		11094 => '0',
		11095 => '1',
		11096 => '0',
		11097 => '1',
		11098 => '0',
		11099 => '1',
		11100 => '0',
		11101 => '1',
		11102 => '0',
		11103 => '1',
		11104 => '0',
		11105 => '1',
		11106 => '0',
		11107 => '1',
		11108 => '0',
		11109 => '1',
		11110 => '0',
		11111 => '1',
		11112 => '0',
		11113 => '1',
		11114 => '0',
		11115 => '1',
		11116 => '0',
		11117 => '1',
		11118 => '0',
		11119 => '1',
		11120 => '0',
		11121 => '1',
		11122 => '0',
		11123 => '1',
		11124 => '0',
		11125 => '1',
		11126 => '0',
		11127 => '1',
		11136 => '1',
		11137 => '0',
		11138 => '1',
		11139 => '0',
		11140 => '1',
		11141 => '0',
		11142 => '1',
		11143 => '0',
		11144 => '1',
		11145 => '0',
		11146 => '1',
		11147 => '0',
		11148 => '1',
		11149 => '0',
		11150 => '1',
		11151 => '0',
		11152 => '1',
		11153 => '0',
		11154 => '1',
		11155 => '0',
		11156 => '1',
		11157 => '0',
		11158 => '1',
		11159 => '0',
		11160 => '1',
		11161 => '0',
		11162 => '1',
		11163 => '0',
		11164 => '1',
		11165 => '0',
		11166 => '1',
		11167 => '0',
		11168 => '1',
		11169 => '0',
		11170 => '1',
		11171 => '0',
		11172 => '1',
		11173 => '0',
		11174 => '1',
		11175 => '0',
		11176 => '1',
		11177 => '0',
		11178 => '1',
		11179 => '0',
		11180 => '1',
		11181 => '0',
		11182 => '1',
		11183 => '0',
		11184 => '1',
		11185 => '0',
		11186 => '1',
		11187 => '0',
		11188 => '1',
		11189 => '0',
		11190 => '1',
		11191 => '0',
		11192 => '1',
		11193 => '0',
		11194 => '1',
		11195 => '0',
		11196 => '1',
		11197 => '0',
		11198 => '1',
		11199 => '0',
		11200 => '1',
		11201 => '0',
		11202 => '1',
		11203 => '0',
		11204 => '1',
		11205 => '0',
		11206 => '1',
		11207 => '0',
		11208 => '1',
		11209 => '0',
		11210 => '1',
		11211 => '0',
		11212 => '1',
		11213 => '0',
		11214 => '1',
		11215 => '0',
		11216 => '1',
		11217 => '0',
		11218 => '1',
		11219 => '0',
		11220 => '1',
		11221 => '0',
		11222 => '1',
		11223 => '0',
		11224 => '1',
		11225 => '0',
		11226 => '1',
		11227 => '0',
		11228 => '1',
		11229 => '0',
		11230 => '1',
		11231 => '0',
		11232 => '1',
		11233 => '0',
		11234 => '1',
		11235 => '0',
		11236 => '1',
		11237 => '0',
		11238 => '1',
		11239 => '0',
		11240 => '1',
		11241 => '0',
		11242 => '1',
		11243 => '0',
		11244 => '1',
		11245 => '0',
		11246 => '1',
		11247 => '0',
		11248 => '1',
		11249 => '0',
		11250 => '1',
		11251 => '0',
		11252 => '1',
		11253 => '0',
		11254 => '1',
		11255 => '0',
		11264 => '0',
		11265 => '1',
		11266 => '0',
		11267 => '1',
		11268 => '0',
		11269 => '1',
		11270 => '0',
		11271 => '1',
		11272 => '0',
		11273 => '1',
		11274 => '0',
		11275 => '1',
		11276 => '0',
		11277 => '1',
		11278 => '0',
		11279 => '1',
		11280 => '0',
		11281 => '1',
		11282 => '0',
		11283 => '1',
		11284 => '0',
		11285 => '1',
		11286 => '0',
		11287 => '1',
		11288 => '0',
		11289 => '1',
		11290 => '0',
		11291 => '1',
		11292 => '0',
		11293 => '1',
		11294 => '0',
		11295 => '1',
		11296 => '0',
		11297 => '1',
		11298 => '0',
		11299 => '1',
		11300 => '0',
		11301 => '1',
		11302 => '0',
		11303 => '1',
		11304 => '0',
		11305 => '1',
		11306 => '0',
		11307 => '1',
		11308 => '0',
		11309 => '1',
		11310 => '0',
		11311 => '1',
		11312 => '0',
		11313 => '1',
		11314 => '0',
		11315 => '1',
		11316 => '0',
		11317 => '1',
		11318 => '0',
		11319 => '1',
		11320 => '0',
		11321 => '1',
		11322 => '0',
		11323 => '1',
		11324 => '0',
		11325 => '1',
		11326 => '0',
		11327 => '1',
		11328 => '0',
		11329 => '1',
		11330 => '0',
		11331 => '1',
		11332 => '0',
		11333 => '1',
		11334 => '0',
		11335 => '1',
		11336 => '0',
		11337 => '1',
		11338 => '0',
		11339 => '1',
		11340 => '0',
		11341 => '1',
		11342 => '0',
		11343 => '1',
		11344 => '0',
		11345 => '1',
		11346 => '0',
		11347 => '1',
		11348 => '0',
		11349 => '1',
		11350 => '0',
		11351 => '1',
		11352 => '0',
		11353 => '1',
		11354 => '0',
		11355 => '1',
		11356 => '0',
		11357 => '1',
		11358 => '0',
		11359 => '1',
		11360 => '0',
		11361 => '1',
		11362 => '0',
		11363 => '1',
		11364 => '0',
		11365 => '1',
		11366 => '0',
		11367 => '1',
		11368 => '0',
		11369 => '1',
		11370 => '0',
		11371 => '1',
		11372 => '0',
		11373 => '1',
		11374 => '0',
		11375 => '1',
		11376 => '0',
		11377 => '1',
		11378 => '0',
		11379 => '1',
		11380 => '0',
		11381 => '1',
		11382 => '0',
		11383 => '1',
		11392 => '1',
		11393 => '0',
		11394 => '1',
		11395 => '0',
		11396 => '1',
		11397 => '0',
		11398 => '1',
		11399 => '0',
		11400 => '1',
		11401 => '0',
		11402 => '1',
		11403 => '0',
		11404 => '1',
		11405 => '0',
		11406 => '1',
		11407 => '0',
		11408 => '1',
		11409 => '0',
		11410 => '1',
		11411 => '0',
		11412 => '1',
		11413 => '0',
		11414 => '1',
		11415 => '0',
		11416 => '1',
		11417 => '0',
		11418 => '1',
		11419 => '0',
		11420 => '1',
		11421 => '0',
		11422 => '1',
		11423 => '0',
		11424 => '1',
		11425 => '0',
		11426 => '1',
		11427 => '0',
		11428 => '1',
		11429 => '0',
		11430 => '1',
		11431 => '0',
		11432 => '1',
		11433 => '0',
		11434 => '1',
		11435 => '0',
		11436 => '1',
		11437 => '0',
		11438 => '1',
		11439 => '0',
		11440 => '1',
		11441 => '0',
		11442 => '1',
		11443 => '0',
		11444 => '1',
		11445 => '0',
		11446 => '1',
		11447 => '0',
		11448 => '1',
		11449 => '0',
		11450 => '1',
		11451 => '0',
		11452 => '1',
		11453 => '0',
		11454 => '1',
		11455 => '0',
		11456 => '1',
		11457 => '0',
		11458 => '1',
		11459 => '0',
		11460 => '1',
		11461 => '0',
		11462 => '1',
		11463 => '0',
		11464 => '1',
		11465 => '0',
		11466 => '1',
		11467 => '0',
		11468 => '1',
		11469 => '0',
		11470 => '1',
		11471 => '0',
		11472 => '1',
		11473 => '0',
		11474 => '1',
		11475 => '0',
		11476 => '1',
		11477 => '0',
		11478 => '1',
		11479 => '0',
		11480 => '1',
		11481 => '0',
		11482 => '1',
		11483 => '0',
		11484 => '1',
		11485 => '0',
		11486 => '1',
		11487 => '0',
		11488 => '1',
		11489 => '0',
		11490 => '1',
		11491 => '0',
		11492 => '1',
		11493 => '0',
		11494 => '1',
		11495 => '0',
		11496 => '1',
		11497 => '0',
		11498 => '1',
		11499 => '0',
		11500 => '1',
		11501 => '0',
		11502 => '1',
		11503 => '0',
		11504 => '1',
		11505 => '0',
		11506 => '1',
		11507 => '0',
		11508 => '1',
		11509 => '0',
		11510 => '1',
		11511 => '0',
		11520 => '0',
		11521 => '1',
		11522 => '0',
		11523 => '1',
		11524 => '0',
		11525 => '1',
		11526 => '0',
		11527 => '1',
		11528 => '0',
		11529 => '1',
		11530 => '0',
		11531 => '1',
		11532 => '0',
		11533 => '1',
		11534 => '0',
		11535 => '1',
		11536 => '0',
		11537 => '1',
		11538 => '0',
		11539 => '1',
		11540 => '0',
		11541 => '1',
		11542 => '0',
		11543 => '1',
		11544 => '0',
		11545 => '1',
		11546 => '0',
		11547 => '1',
		11548 => '0',
		11549 => '1',
		11550 => '0',
		11551 => '1',
		11552 => '0',
		11553 => '1',
		11554 => '0',
		11555 => '1',
		11556 => '0',
		11557 => '1',
		11558 => '0',
		11559 => '1',
		11560 => '0',
		11561 => '1',
		11562 => '0',
		11563 => '1',
		11564 => '0',
		11565 => '1',
		11566 => '0',
		11567 => '1',
		11568 => '0',
		11569 => '1',
		11570 => '0',
		11571 => '1',
		11572 => '0',
		11573 => '1',
		11574 => '0',
		11575 => '1',
		11576 => '0',
		11577 => '1',
		11578 => '0',
		11579 => '1',
		11580 => '0',
		11581 => '1',
		11582 => '0',
		11583 => '1',
		11584 => '0',
		11585 => '1',
		11586 => '0',
		11587 => '1',
		11588 => '0',
		11589 => '1',
		11590 => '0',
		11591 => '1',
		11592 => '0',
		11593 => '1',
		11594 => '0',
		11595 => '1',
		11596 => '0',
		11597 => '1',
		11598 => '0',
		11599 => '1',
		11600 => '0',
		11601 => '1',
		11602 => '0',
		11603 => '1',
		11604 => '0',
		11605 => '1',
		11606 => '0',
		11607 => '1',
		11608 => '0',
		11609 => '1',
		11610 => '0',
		11611 => '1',
		11612 => '0',
		11613 => '1',
		11614 => '0',
		11615 => '1',
		11616 => '0',
		11617 => '1',
		11618 => '0',
		11619 => '1',
		11620 => '0',
		11621 => '1',
		11622 => '0',
		11623 => '1',
		11624 => '0',
		11625 => '1',
		11626 => '0',
		11627 => '1',
		11628 => '0',
		11629 => '1',
		11630 => '0',
		11631 => '1',
		11632 => '0',
		11633 => '1',
		11634 => '0',
		11635 => '1',
		11636 => '0',
		11637 => '1',
		11638 => '0',
		11639 => '1',
		11648 => '1',
		11649 => '0',
		11650 => '1',
		11651 => '0',
		11652 => '1',
		11653 => '0',
		11654 => '1',
		11655 => '0',
		11656 => '1',
		11657 => '0',
		11658 => '1',
		11659 => '0',
		11660 => '1',
		11661 => '0',
		11662 => '1',
		11663 => '0',
		11664 => '1',
		11665 => '0',
		11666 => '1',
		11667 => '0',
		11668 => '1',
		11669 => '0',
		11670 => '1',
		11671 => '0',
		11672 => '1',
		11673 => '0',
		11674 => '1',
		11675 => '0',
		11676 => '1',
		11677 => '0',
		11678 => '1',
		11679 => '0',
		11680 => '1',
		11681 => '0',
		11682 => '1',
		11683 => '0',
		11684 => '1',
		11685 => '0',
		11686 => '1',
		11687 => '0',
		11688 => '1',
		11689 => '0',
		11690 => '1',
		11691 => '0',
		11692 => '1',
		11693 => '0',
		11694 => '1',
		11695 => '0',
		11696 => '1',
		11697 => '0',
		11698 => '1',
		11699 => '0',
		11700 => '1',
		11701 => '0',
		11702 => '1',
		11703 => '0',
		11704 => '1',
		11705 => '0',
		11706 => '1',
		11707 => '0',
		11708 => '1',
		11709 => '0',
		11710 => '1',
		11711 => '0',
		11712 => '1',
		11713 => '0',
		11714 => '1',
		11715 => '0',
		11716 => '1',
		11717 => '0',
		11718 => '1',
		11719 => '0',
		11720 => '1',
		11721 => '0',
		11722 => '1',
		11723 => '0',
		11724 => '1',
		11725 => '0',
		11726 => '1',
		11727 => '0',
		11728 => '1',
		11729 => '0',
		11730 => '1',
		11731 => '0',
		11732 => '1',
		11733 => '0',
		11734 => '1',
		11735 => '0',
		11736 => '1',
		11737 => '0',
		11738 => '1',
		11739 => '0',
		11740 => '1',
		11741 => '0',
		11742 => '1',
		11743 => '0',
		11744 => '1',
		11745 => '0',
		11746 => '1',
		11747 => '0',
		11748 => '1',
		11749 => '0',
		11750 => '1',
		11751 => '0',
		11752 => '1',
		11753 => '0',
		11754 => '1',
		11755 => '0',
		11756 => '1',
		11757 => '0',
		11758 => '1',
		11759 => '0',
		11760 => '1',
		11761 => '0',
		11762 => '1',
		11763 => '0',
		11764 => '1',
		11765 => '0',
		11766 => '1',
		11767 => '0',
		11776 => '0',
		11777 => '1',
		11778 => '0',
		11779 => '1',
		11780 => '0',
		11781 => '1',
		11782 => '0',
		11783 => '1',
		11784 => '0',
		11785 => '1',
		11786 => '0',
		11787 => '1',
		11788 => '0',
		11789 => '1',
		11790 => '0',
		11791 => '1',
		11792 => '0',
		11793 => '1',
		11794 => '0',
		11795 => '1',
		11796 => '0',
		11797 => '1',
		11798 => '0',
		11799 => '1',
		11800 => '0',
		11801 => '1',
		11802 => '0',
		11803 => '1',
		11804 => '0',
		11805 => '1',
		11806 => '0',
		11807 => '1',
		11808 => '0',
		11809 => '1',
		11810 => '0',
		11811 => '1',
		11812 => '0',
		11813 => '1',
		11814 => '0',
		11815 => '1',
		11816 => '0',
		11817 => '1',
		11818 => '0',
		11819 => '1',
		11820 => '0',
		11821 => '1',
		11822 => '0',
		11823 => '1',
		11824 => '0',
		11825 => '1',
		11826 => '0',
		11827 => '1',
		11828 => '0',
		11829 => '1',
		11830 => '0',
		11831 => '1',
		11832 => '0',
		11833 => '1',
		11834 => '0',
		11835 => '1',
		11836 => '0',
		11837 => '1',
		11838 => '0',
		11839 => '1',
		11840 => '0',
		11841 => '1',
		11842 => '0',
		11843 => '1',
		11844 => '0',
		11845 => '1',
		11846 => '0',
		11847 => '1',
		11848 => '0',
		11849 => '1',
		11850 => '0',
		11851 => '1',
		11852 => '0',
		11853 => '1',
		11854 => '0',
		11855 => '1',
		11856 => '0',
		11857 => '1',
		11858 => '0',
		11859 => '1',
		11860 => '0',
		11861 => '1',
		11862 => '0',
		11863 => '1',
		11864 => '0',
		11865 => '1',
		11866 => '0',
		11867 => '1',
		11868 => '0',
		11869 => '1',
		11870 => '0',
		11871 => '1',
		11872 => '0',
		11873 => '1',
		11874 => '0',
		11875 => '1',
		11876 => '0',
		11877 => '1',
		11878 => '0',
		11879 => '1',
		11880 => '0',
		11881 => '1',
		11882 => '0',
		11883 => '1',
		11884 => '0',
		11885 => '1',
		11886 => '0',
		11887 => '1',
		11888 => '0',
		11889 => '1',
		11890 => '0',
		11891 => '1',
		11892 => '0',
		11893 => '1',
		11894 => '0',
		11895 => '1',
		11904 => '1',
		11905 => '0',
		11906 => '1',
		11907 => '0',
		11908 => '1',
		11909 => '0',
		11910 => '1',
		11911 => '0',
		11912 => '1',
		11913 => '0',
		11914 => '1',
		11915 => '0',
		11916 => '1',
		11917 => '0',
		11918 => '1',
		11919 => '0',
		11920 => '1',
		11921 => '0',
		11922 => '1',
		11923 => '0',
		11924 => '1',
		11925 => '0',
		11926 => '1',
		11927 => '0',
		11928 => '1',
		11929 => '0',
		11930 => '1',
		11931 => '0',
		11932 => '1',
		11933 => '0',
		11934 => '1',
		11935 => '0',
		11936 => '1',
		11937 => '0',
		11938 => '1',
		11939 => '0',
		11940 => '1',
		11941 => '0',
		11942 => '1',
		11943 => '0',
		11944 => '1',
		11945 => '0',
		11946 => '1',
		11947 => '0',
		11948 => '1',
		11949 => '0',
		11950 => '1',
		11951 => '0',
		11952 => '1',
		11953 => '0',
		11954 => '1',
		11955 => '0',
		11956 => '1',
		11957 => '0',
		11958 => '1',
		11959 => '0',
		11960 => '1',
		11961 => '0',
		11962 => '1',
		11963 => '0',
		11964 => '1',
		11965 => '0',
		11966 => '1',
		11967 => '0',
		11968 => '1',
		11969 => '0',
		11970 => '1',
		11971 => '0',
		11972 => '1',
		11973 => '0',
		11974 => '1',
		11975 => '0',
		11976 => '1',
		11977 => '0',
		11978 => '1',
		11979 => '0',
		11980 => '1',
		11981 => '0',
		11982 => '1',
		11983 => '0',
		11984 => '1',
		11985 => '0',
		11986 => '1',
		11987 => '0',
		11988 => '1',
		11989 => '0',
		11990 => '1',
		11991 => '0',
		11992 => '1',
		11993 => '0',
		11994 => '1',
		11995 => '0',
		11996 => '1',
		11997 => '0',
		11998 => '1',
		11999 => '0',
		12000 => '1',
		12001 => '0',
		12002 => '1',
		12003 => '0',
		12004 => '1',
		12005 => '0',
		12006 => '1',
		12007 => '0',
		12008 => '1',
		12009 => '0',
		12010 => '1',
		12011 => '0',
		12012 => '1',
		12013 => '0',
		12014 => '1',
		12015 => '0',
		12016 => '1',
		12017 => '0',
		12018 => '1',
		12019 => '0',
		12020 => '1',
		12021 => '0',
		12022 => '1',
		12023 => '0',
		12032 => '0',
		12033 => '1',
		12034 => '0',
		12035 => '1',
		12036 => '0',
		12037 => '1',
		12038 => '0',
		12039 => '1',
		12040 => '0',
		12041 => '1',
		12042 => '0',
		12043 => '1',
		12044 => '0',
		12045 => '1',
		12046 => '0',
		12047 => '1',
		12048 => '0',
		12049 => '1',
		12050 => '0',
		12051 => '1',
		12052 => '0',
		12053 => '1',
		12054 => '0',
		12055 => '1',
		12056 => '0',
		12057 => '1',
		12058 => '0',
		12059 => '1',
		12060 => '0',
		12061 => '1',
		12062 => '0',
		12063 => '1',
		12064 => '0',
		12065 => '1',
		12066 => '0',
		12067 => '1',
		12068 => '0',
		12069 => '1',
		12070 => '0',
		12071 => '1',
		12072 => '0',
		12073 => '1',
		12074 => '0',
		12075 => '1',
		12076 => '0',
		12077 => '1',
		12078 => '0',
		12079 => '1',
		12080 => '0',
		12081 => '1',
		12082 => '0',
		12083 => '1',
		12084 => '0',
		12085 => '1',
		12086 => '0',
		12087 => '1',
		12088 => '0',
		12089 => '1',
		12090 => '0',
		12091 => '1',
		12092 => '0',
		12093 => '1',
		12094 => '0',
		12095 => '1',
		12096 => '0',
		12097 => '1',
		12098 => '0',
		12099 => '1',
		12100 => '0',
		12101 => '1',
		12102 => '0',
		12103 => '1',
		12104 => '0',
		12105 => '1',
		12106 => '0',
		12107 => '1',
		12108 => '0',
		12109 => '1',
		12110 => '0',
		12111 => '1',
		12112 => '0',
		12113 => '1',
		12114 => '0',
		12115 => '1',
		12116 => '0',
		12117 => '1',
		12118 => '0',
		12119 => '1',
		12120 => '0',
		12121 => '1',
		12122 => '0',
		12123 => '1',
		12124 => '0',
		12125 => '1',
		12126 => '0',
		12127 => '1',
		12128 => '0',
		12129 => '1',
		12130 => '0',
		12131 => '1',
		12132 => '0',
		12133 => '1',
		12134 => '0',
		12135 => '1',
		12136 => '0',
		12137 => '1',
		12138 => '0',
		12139 => '1',
		12140 => '0',
		12141 => '1',
		12142 => '0',
		12143 => '1',
		12144 => '0',
		12145 => '1',
		12146 => '0',
		12147 => '1',
		12148 => '0',
		12149 => '1',
		12150 => '0',
		12151 => '1',
		12160 => '1',
		12161 => '0',
		12162 => '1',
		12163 => '0',
		12164 => '1',
		12165 => '0',
		12166 => '1',
		12167 => '0',
		12168 => '1',
		12169 => '0',
		12170 => '1',
		12171 => '0',
		12172 => '1',
		12173 => '0',
		12174 => '1',
		12175 => '0',
		12176 => '1',
		12177 => '0',
		12178 => '1',
		12179 => '0',
		12180 => '1',
		12181 => '0',
		12182 => '1',
		12183 => '0',
		12184 => '1',
		12185 => '0',
		12186 => '1',
		12187 => '0',
		12188 => '1',
		12189 => '0',
		12190 => '1',
		12191 => '0',
		12192 => '1',
		12193 => '0',
		12194 => '1',
		12195 => '0',
		12196 => '1',
		12197 => '0',
		12198 => '1',
		12199 => '0',
		12200 => '1',
		12201 => '0',
		12202 => '1',
		12203 => '0',
		12204 => '1',
		12205 => '0',
		12206 => '1',
		12207 => '0',
		12208 => '1',
		12209 => '0',
		12210 => '1',
		12211 => '0',
		12212 => '1',
		12213 => '0',
		12214 => '1',
		12215 => '0',
		12216 => '1',
		12217 => '0',
		12218 => '1',
		12219 => '0',
		12220 => '1',
		12221 => '0',
		12222 => '1',
		12223 => '0',
		12224 => '1',
		12225 => '0',
		12226 => '1',
		12227 => '0',
		12228 => '1',
		12229 => '0',
		12230 => '1',
		12231 => '0',
		12232 => '1',
		12233 => '0',
		12234 => '1',
		12235 => '0',
		12236 => '1',
		12237 => '0',
		12238 => '1',
		12239 => '0',
		12240 => '1',
		12241 => '0',
		12242 => '1',
		12243 => '0',
		12244 => '1',
		12245 => '0',
		12246 => '1',
		12247 => '0',
		12248 => '1',
		12249 => '0',
		12250 => '1',
		12251 => '0',
		12252 => '1',
		12253 => '0',
		12254 => '1',
		12255 => '0',
		12256 => '1',
		12257 => '0',
		12258 => '1',
		12259 => '0',
		12260 => '1',
		12261 => '0',
		12262 => '1',
		12263 => '0',
		12264 => '1',
		12265 => '0',
		12266 => '1',
		12267 => '0',
		12268 => '1',
		12269 => '0',
		12270 => '1',
		12271 => '0',
		12272 => '1',
		12273 => '0',
		12274 => '1',
		12275 => '0',
		12276 => '1',
		12277 => '0',
		12278 => '1',
		12279 => '0',
		12288 => '0',
		12289 => '1',
		12290 => '0',
		12291 => '1',
		12292 => '0',
		12293 => '1',
		12294 => '0',
		12295 => '1',
		12296 => '0',
		12297 => '1',
		12298 => '0',
		12299 => '1',
		12300 => '0',
		12301 => '1',
		12302 => '0',
		12303 => '1',
		12304 => '0',
		12305 => '1',
		12306 => '0',
		12307 => '1',
		12308 => '0',
		12309 => '1',
		12310 => '0',
		12311 => '1',
		12312 => '0',
		12313 => '1',
		12314 => '0',
		12315 => '1',
		12316 => '0',
		12317 => '1',
		12318 => '0',
		12319 => '1',
		12320 => '0',
		12321 => '1',
		12322 => '0',
		12323 => '1',
		12324 => '0',
		12325 => '1',
		12326 => '0',
		12327 => '1',
		12328 => '0',
		12329 => '1',
		12330 => '0',
		12331 => '1',
		12332 => '0',
		12333 => '1',
		12334 => '0',
		12335 => '1',
		12336 => '0',
		12337 => '1',
		12338 => '0',
		12339 => '1',
		12340 => '0',
		12341 => '1',
		12342 => '0',
		12343 => '1',
		12344 => '0',
		12345 => '1',
		12346 => '0',
		12347 => '1',
		12348 => '0',
		12349 => '1',
		12350 => '0',
		12351 => '1',
		12352 => '0',
		12353 => '1',
		12354 => '0',
		12355 => '1',
		12356 => '0',
		12357 => '1',
		12358 => '0',
		12359 => '1',
		12360 => '0',
		12361 => '1',
		12362 => '0',
		12363 => '1',
		12364 => '0',
		12365 => '1',
		12366 => '0',
		12367 => '1',
		12368 => '0',
		12369 => '1',
		12370 => '0',
		12371 => '1',
		12372 => '0',
		12373 => '1',
		12374 => '0',
		12375 => '1',
		12376 => '0',
		12377 => '1',
		12378 => '0',
		12379 => '1',
		12380 => '0',
		12381 => '1',
		12382 => '0',
		12383 => '1',
		12384 => '0',
		12385 => '1',
		12386 => '0',
		12387 => '1',
		12388 => '0',
		12389 => '1',
		12390 => '0',
		12391 => '1',
		12392 => '0',
		12393 => '1',
		12394 => '0',
		12395 => '1',
		12396 => '0',
		12397 => '1',
		12398 => '0',
		12399 => '1',
		12400 => '0',
		12401 => '1',
		12402 => '0',
		12403 => '1',
		12404 => '0',
		12405 => '1',
		12406 => '0',
		12407 => '1',
		12416 => '1',
		12417 => '0',
		12418 => '1',
		12419 => '0',
		12420 => '1',
		12421 => '0',
		12422 => '1',
		12423 => '0',
		12424 => '1',
		12425 => '0',
		12426 => '1',
		12427 => '0',
		12428 => '1',
		12429 => '0',
		12430 => '1',
		12431 => '0',
		12432 => '1',
		12433 => '0',
		12434 => '1',
		12435 => '0',
		12436 => '1',
		12437 => '0',
		12438 => '1',
		12439 => '0',
		12440 => '1',
		12441 => '0',
		12442 => '1',
		12443 => '0',
		12444 => '1',
		12445 => '0',
		12446 => '1',
		12447 => '0',
		12448 => '1',
		12449 => '0',
		12450 => '1',
		12451 => '0',
		12452 => '1',
		12453 => '0',
		12454 => '1',
		12455 => '0',
		12456 => '1',
		12457 => '0',
		12458 => '1',
		12459 => '0',
		12460 => '1',
		12461 => '0',
		12462 => '1',
		12463 => '0',
		12464 => '1',
		12465 => '0',
		12466 => '1',
		12467 => '0',
		12468 => '1',
		12469 => '0',
		12470 => '1',
		12471 => '0',
		12472 => '1',
		12473 => '0',
		12474 => '1',
		12475 => '0',
		12476 => '1',
		12477 => '0',
		12478 => '1',
		12479 => '0',
		12480 => '1',
		12481 => '0',
		12482 => '1',
		12483 => '0',
		12484 => '1',
		12485 => '0',
		12486 => '1',
		12487 => '0',
		12488 => '1',
		12489 => '0',
		12490 => '1',
		12491 => '0',
		12492 => '1',
		12493 => '0',
		12494 => '1',
		12495 => '0',
		12496 => '1',
		12497 => '0',
		12498 => '1',
		12499 => '0',
		12500 => '1',
		12501 => '0',
		12502 => '1',
		12503 => '0',
		12504 => '1',
		12505 => '0',
		12506 => '1',
		12507 => '0',
		12508 => '1',
		12509 => '0',
		12510 => '1',
		12511 => '0',
		12512 => '1',
		12513 => '0',
		12514 => '1',
		12515 => '0',
		12516 => '1',
		12517 => '0',
		12518 => '1',
		12519 => '0',
		12520 => '1',
		12521 => '0',
		12522 => '1',
		12523 => '0',
		12524 => '1',
		12525 => '0',
		12526 => '1',
		12527 => '0',
		12528 => '1',
		12529 => '0',
		12530 => '1',
		12531 => '0',
		12532 => '1',
		12533 => '0',
		12534 => '1',
		12535 => '0',
		12544 => '0',
		12545 => '1',
		12546 => '0',
		12547 => '1',
		12548 => '0',
		12549 => '1',
		12550 => '0',
		12551 => '1',
		12552 => '0',
		12553 => '1',
		12554 => '0',
		12555 => '1',
		12556 => '0',
		12557 => '1',
		12558 => '0',
		12559 => '1',
		12560 => '0',
		12561 => '1',
		12562 => '0',
		12563 => '1',
		12564 => '0',
		12565 => '1',
		12566 => '0',
		12567 => '1',
		12568 => '0',
		12569 => '1',
		12570 => '0',
		12571 => '1',
		12572 => '0',
		12573 => '1',
		12574 => '0',
		12575 => '1',
		12576 => '0',
		12577 => '1',
		12578 => '0',
		12579 => '1',
		12580 => '0',
		12581 => '1',
		12582 => '0',
		12583 => '1',
		12584 => '0',
		12585 => '1',
		12586 => '0',
		12587 => '1',
		12588 => '0',
		12589 => '1',
		12590 => '0',
		12591 => '1',
		12592 => '0',
		12593 => '1',
		12594 => '0',
		12595 => '1',
		12596 => '0',
		12597 => '1',
		12598 => '0',
		12599 => '1',
		12600 => '0',
		12601 => '1',
		12602 => '0',
		12603 => '1',
		12604 => '0',
		12605 => '1',
		12606 => '0',
		12607 => '1',
		12608 => '0',
		12609 => '1',
		12610 => '0',
		12611 => '1',
		12612 => '0',
		12613 => '1',
		12614 => '0',
		12615 => '1',
		12616 => '0',
		12617 => '1',
		12618 => '0',
		12619 => '1',
		12620 => '0',
		12621 => '1',
		12622 => '0',
		12623 => '1',
		12624 => '0',
		12625 => '1',
		12626 => '0',
		12627 => '1',
		12628 => '0',
		12629 => '1',
		12630 => '0',
		12631 => '1',
		12632 => '0',
		12633 => '1',
		12634 => '0',
		12635 => '1',
		12636 => '0',
		12637 => '1',
		12638 => '0',
		12639 => '1',
		12640 => '0',
		12641 => '1',
		12642 => '0',
		12643 => '1',
		12644 => '0',
		12645 => '1',
		12646 => '0',
		12647 => '1',
		12648 => '0',
		12649 => '1',
		12650 => '0',
		12651 => '1',
		12652 => '0',
		12653 => '1',
		12654 => '0',
		12655 => '1',
		12656 => '0',
		12657 => '1',
		12658 => '0',
		12659 => '1',
		12660 => '0',
		12661 => '1',
		12662 => '0',
		12663 => '1',
		12672 => '1',
		12673 => '0',
		12674 => '1',
		12675 => '0',
		12676 => '1',
		12677 => '0',
		12678 => '1',
		12679 => '0',
		12680 => '1',
		12681 => '0',
		12682 => '1',
		12683 => '0',
		12684 => '1',
		12685 => '0',
		12686 => '1',
		12687 => '0',
		12688 => '1',
		12689 => '0',
		12690 => '1',
		12691 => '0',
		12692 => '1',
		12693 => '0',
		12694 => '1',
		12695 => '0',
		12696 => '1',
		12697 => '0',
		12698 => '1',
		12699 => '0',
		12700 => '1',
		12701 => '0',
		12702 => '1',
		12703 => '0',
		12704 => '1',
		12705 => '0',
		12706 => '1',
		12707 => '0',
		12708 => '1',
		12709 => '0',
		12710 => '1',
		12711 => '0',
		12712 => '1',
		12713 => '0',
		12714 => '1',
		12715 => '0',
		12716 => '1',
		12717 => '0',
		12718 => '1',
		12719 => '0',
		12720 => '1',
		12721 => '0',
		12722 => '1',
		12723 => '0',
		12724 => '1',
		12725 => '0',
		12726 => '1',
		12727 => '0',
		12728 => '1',
		12729 => '0',
		12730 => '1',
		12731 => '0',
		12732 => '1',
		12733 => '0',
		12734 => '1',
		12735 => '0',
		12736 => '1',
		12737 => '0',
		12738 => '1',
		12739 => '0',
		12740 => '1',
		12741 => '0',
		12742 => '1',
		12743 => '0',
		12744 => '1',
		12745 => '0',
		12746 => '1',
		12747 => '0',
		12748 => '1',
		12749 => '0',
		12750 => '1',
		12751 => '0',
		12752 => '1',
		12753 => '0',
		12754 => '1',
		12755 => '0',
		12756 => '1',
		12757 => '0',
		12758 => '1',
		12759 => '0',
		12760 => '1',
		12761 => '0',
		12762 => '1',
		12763 => '0',
		12764 => '1',
		12765 => '0',
		12766 => '1',
		12767 => '0',
		12768 => '1',
		12769 => '0',
		12770 => '1',
		12771 => '0',
		12772 => '1',
		12773 => '0',
		12774 => '1',
		12775 => '0',
		12776 => '1',
		12777 => '0',
		12778 => '1',
		12779 => '0',
		12780 => '1',
		12781 => '0',
		12782 => '1',
		12783 => '0',
		12784 => '1',
		12785 => '0',
		12786 => '1',
		12787 => '0',
		12788 => '1',
		12789 => '0',
		12790 => '1',
		12791 => '0',
		12800 => '0',
		12801 => '1',
		12802 => '0',
		12803 => '1',
		12804 => '0',
		12805 => '1',
		12806 => '0',
		12807 => '1',
		12808 => '0',
		12809 => '1',
		12810 => '0',
		12811 => '1',
		12812 => '0',
		12813 => '1',
		12814 => '0',
		12815 => '1',
		12816 => '0',
		12817 => '1',
		12818 => '0',
		12819 => '1',
		12820 => '0',
		12821 => '1',
		12822 => '0',
		12823 => '1',
		12824 => '0',
		12825 => '1',
		12826 => '0',
		12827 => '1',
		12828 => '0',
		12829 => '1',
		12830 => '0',
		12831 => '1',
		12832 => '0',
		12833 => '1',
		12834 => '0',
		12835 => '1',
		12836 => '0',
		12837 => '1',
		12838 => '0',
		12839 => '1',
		12840 => '0',
		12841 => '1',
		12842 => '0',
		12843 => '1',
		12844 => '0',
		12845 => '1',
		12846 => '0',
		12847 => '1',
		12848 => '0',
		12849 => '1',
		12850 => '0',
		12851 => '1',
		12852 => '0',
		12853 => '1',
		12854 => '0',
		12855 => '1',
		12856 => '0',
		12857 => '1',
		12858 => '0',
		12859 => '1',
		12860 => '0',
		12861 => '1',
		12862 => '0',
		12863 => '1',
		12864 => '0',
		12865 => '1',
		12866 => '0',
		12867 => '1',
		12868 => '0',
		12869 => '1',
		12870 => '0',
		12871 => '1',
		12872 => '0',
		12873 => '1',
		12874 => '0',
		12875 => '1',
		12876 => '0',
		12877 => '1',
		12878 => '0',
		12879 => '1',
		12880 => '0',
		12881 => '1',
		12882 => '0',
		12883 => '1',
		12884 => '0',
		12885 => '1',
		12886 => '0',
		12887 => '1',
		12888 => '0',
		12889 => '1',
		12890 => '0',
		12891 => '1',
		12892 => '0',
		12893 => '1',
		12894 => '0',
		12895 => '1',
		12896 => '0',
		12897 => '1',
		12898 => '0',
		12899 => '1',
		12900 => '0',
		12901 => '1',
		12902 => '0',
		12903 => '1',
		12904 => '0',
		12905 => '1',
		12906 => '0',
		12907 => '1',
		12908 => '0',
		12909 => '1',
		12910 => '0',
		12911 => '1',
		12912 => '0',
		12913 => '1',
		12914 => '0',
		12915 => '1',
		12916 => '0',
		12917 => '1',
		12918 => '0',
		12919 => '1',
		12928 => '1',
		12929 => '0',
		12930 => '1',
		12931 => '0',
		12932 => '1',
		12933 => '0',
		12934 => '1',
		12935 => '0',
		12936 => '1',
		12937 => '0',
		12938 => '1',
		12939 => '0',
		12940 => '1',
		12941 => '0',
		12942 => '1',
		12943 => '0',
		12944 => '1',
		12945 => '0',
		12946 => '1',
		12947 => '0',
		12948 => '1',
		12949 => '0',
		12950 => '1',
		12951 => '0',
		12952 => '1',
		12953 => '0',
		12954 => '1',
		12955 => '0',
		12956 => '1',
		12957 => '0',
		12958 => '1',
		12959 => '0',
		12960 => '1',
		12961 => '0',
		12962 => '1',
		12963 => '0',
		12964 => '1',
		12965 => '0',
		12966 => '1',
		12967 => '0',
		12968 => '1',
		12969 => '0',
		12970 => '1',
		12971 => '0',
		12972 => '1',
		12973 => '0',
		12974 => '1',
		12975 => '0',
		12976 => '1',
		12977 => '0',
		12978 => '1',
		12979 => '0',
		12980 => '1',
		12981 => '0',
		12982 => '1',
		12983 => '0',
		12984 => '1',
		12985 => '0',
		12986 => '1',
		12987 => '0',
		12988 => '1',
		12989 => '0',
		12990 => '1',
		12991 => '0',
		12992 => '1',
		12993 => '0',
		12994 => '1',
		12995 => '0',
		12996 => '1',
		12997 => '0',
		12998 => '1',
		12999 => '0',
		13000 => '1',
		13001 => '0',
		13002 => '1',
		13003 => '0',
		13004 => '1',
		13005 => '0',
		13006 => '1',
		13007 => '0',
		13008 => '1',
		13009 => '0',
		13010 => '1',
		13011 => '0',
		13012 => '1',
		13013 => '0',
		13014 => '1',
		13015 => '0',
		13016 => '1',
		13017 => '0',
		13018 => '1',
		13019 => '0',
		13020 => '1',
		13021 => '0',
		13022 => '1',
		13023 => '0',
		13024 => '1',
		13025 => '0',
		13026 => '1',
		13027 => '0',
		13028 => '1',
		13029 => '0',
		13030 => '1',
		13031 => '0',
		13032 => '1',
		13033 => '0',
		13034 => '1',
		13035 => '0',
		13036 => '1',
		13037 => '0',
		13038 => '1',
		13039 => '0',
		13040 => '1',
		13041 => '0',
		13042 => '1',
		13043 => '0',
		13044 => '1',
		13045 => '0',
		13046 => '1',
		13047 => '0',
		13056 => '0',
		13057 => '1',
		13058 => '0',
		13059 => '1',
		13060 => '0',
		13061 => '1',
		13062 => '0',
		13063 => '1',
		13064 => '0',
		13065 => '1',
		13066 => '0',
		13067 => '1',
		13068 => '0',
		13069 => '1',
		13070 => '0',
		13071 => '1',
		13072 => '0',
		13073 => '1',
		13074 => '0',
		13075 => '1',
		13076 => '0',
		13077 => '1',
		13078 => '0',
		13079 => '1',
		13080 => '0',
		13081 => '1',
		13082 => '0',
		13083 => '1',
		13084 => '0',
		13085 => '1',
		13086 => '0',
		13087 => '1',
		13088 => '0',
		13089 => '1',
		13090 => '0',
		13091 => '1',
		13092 => '0',
		13093 => '1',
		13094 => '0',
		13095 => '1',
		13096 => '0',
		13097 => '1',
		13098 => '0',
		13099 => '1',
		13100 => '0',
		13101 => '1',
		13102 => '0',
		13103 => '1',
		13104 => '0',
		13105 => '1',
		13106 => '0',
		13107 => '1',
		13108 => '0',
		13109 => '1',
		13110 => '0',
		13111 => '1',
		13112 => '0',
		13113 => '1',
		13114 => '0',
		13115 => '1',
		13116 => '0',
		13117 => '1',
		13118 => '0',
		13119 => '1',
		13120 => '0',
		13121 => '1',
		13122 => '0',
		13123 => '1',
		13124 => '0',
		13125 => '1',
		13126 => '0',
		13127 => '1',
		13128 => '0',
		13129 => '1',
		13130 => '0',
		13131 => '1',
		13132 => '0',
		13133 => '1',
		13134 => '0',
		13135 => '1',
		13136 => '0',
		13137 => '1',
		13138 => '0',
		13139 => '1',
		13140 => '0',
		13141 => '1',
		13142 => '0',
		13143 => '1',
		13144 => '0',
		13145 => '1',
		13146 => '0',
		13147 => '1',
		13148 => '0',
		13149 => '1',
		13150 => '0',
		13151 => '1',
		13152 => '0',
		13153 => '1',
		13154 => '0',
		13155 => '1',
		13156 => '0',
		13157 => '1',
		13158 => '0',
		13159 => '1',
		13160 => '0',
		13161 => '1',
		13162 => '0',
		13163 => '1',
		13164 => '0',
		13165 => '1',
		13166 => '0',
		13167 => '1',
		13168 => '0',
		13169 => '1',
		13170 => '0',
		13171 => '1',
		13172 => '0',
		13173 => '1',
		13174 => '0',
		13175 => '1',
		13184 => '1',
		13185 => '0',
		13186 => '1',
		13187 => '0',
		13188 => '1',
		13189 => '0',
		13190 => '1',
		13191 => '0',
		13192 => '1',
		13193 => '0',
		13194 => '1',
		13195 => '0',
		13196 => '1',
		13197 => '0',
		13198 => '1',
		13199 => '0',
		13200 => '1',
		13201 => '0',
		13202 => '1',
		13203 => '0',
		13204 => '1',
		13205 => '0',
		13206 => '1',
		13207 => '0',
		13208 => '1',
		13209 => '0',
		13210 => '1',
		13211 => '0',
		13212 => '1',
		13213 => '0',
		13214 => '1',
		13215 => '0',
		13216 => '1',
		13217 => '0',
		13218 => '1',
		13219 => '0',
		13220 => '1',
		13221 => '0',
		13222 => '1',
		13223 => '0',
		13224 => '1',
		13225 => '0',
		13226 => '1',
		13227 => '0',
		13228 => '1',
		13229 => '0',
		13230 => '1',
		13231 => '0',
		13232 => '1',
		13233 => '0',
		13234 => '1',
		13235 => '0',
		13236 => '1',
		13237 => '0',
		13238 => '1',
		13239 => '0',
		13240 => '1',
		13241 => '0',
		13242 => '1',
		13243 => '0',
		13244 => '1',
		13245 => '0',
		13246 => '1',
		13247 => '0',
		13248 => '1',
		13249 => '0',
		13250 => '1',
		13251 => '0',
		13252 => '1',
		13253 => '0',
		13254 => '1',
		13255 => '0',
		13256 => '1',
		13257 => '0',
		13258 => '1',
		13259 => '0',
		13260 => '1',
		13261 => '0',
		13262 => '1',
		13263 => '0',
		13264 => '1',
		13265 => '0',
		13266 => '1',
		13267 => '0',
		13268 => '1',
		13269 => '0',
		13270 => '1',
		13271 => '0',
		13272 => '1',
		13273 => '0',
		13274 => '1',
		13275 => '0',
		13276 => '1',
		13277 => '0',
		13278 => '1',
		13279 => '0',
		13280 => '1',
		13281 => '0',
		13282 => '1',
		13283 => '0',
		13284 => '1',
		13285 => '0',
		13286 => '1',
		13287 => '0',
		13288 => '1',
		13289 => '0',
		13290 => '1',
		13291 => '0',
		13292 => '1',
		13293 => '0',
		13294 => '1',
		13295 => '0',
		13296 => '1',
		13297 => '0',
		13298 => '1',
		13299 => '0',
		13300 => '1',
		13301 => '0',
		13302 => '1',
		13303 => '0',
		13312 => '0',
		13313 => '1',
		13314 => '0',
		13315 => '1',
		13316 => '0',
		13317 => '1',
		13318 => '0',
		13319 => '1',
		13320 => '0',
		13321 => '1',
		13322 => '0',
		13323 => '1',
		13324 => '0',
		13325 => '1',
		13326 => '0',
		13327 => '1',
		13328 => '0',
		13329 => '1',
		13330 => '0',
		13331 => '1',
		13332 => '0',
		13333 => '1',
		13334 => '0',
		13335 => '1',
		13336 => '0',
		13337 => '1',
		13338 => '0',
		13339 => '1',
		13340 => '0',
		13341 => '1',
		13342 => '0',
		13343 => '1',
		13344 => '0',
		13345 => '1',
		13346 => '0',
		13347 => '1',
		13348 => '0',
		13349 => '1',
		13350 => '0',
		13351 => '1',
		13352 => '0',
		13353 => '1',
		13354 => '0',
		13355 => '1',
		13356 => '0',
		13357 => '1',
		13358 => '0',
		13359 => '1',
		13360 => '0',
		13361 => '1',
		13362 => '0',
		13363 => '1',
		13364 => '0',
		13365 => '1',
		13366 => '0',
		13367 => '1',
		13368 => '0',
		13369 => '1',
		13370 => '0',
		13371 => '1',
		13372 => '0',
		13373 => '1',
		13374 => '0',
		13375 => '1',
		13376 => '0',
		13377 => '1',
		13378 => '0',
		13379 => '1',
		13380 => '0',
		13381 => '1',
		13382 => '0',
		13383 => '1',
		13384 => '0',
		13385 => '1',
		13386 => '0',
		13387 => '1',
		13388 => '0',
		13389 => '1',
		13390 => '0',
		13391 => '1',
		13392 => '0',
		13393 => '1',
		13394 => '0',
		13395 => '1',
		13396 => '0',
		13397 => '1',
		13398 => '0',
		13399 => '1',
		13400 => '0',
		13401 => '1',
		13402 => '0',
		13403 => '1',
		13404 => '0',
		13405 => '1',
		13406 => '0',
		13407 => '1',
		13408 => '0',
		13409 => '1',
		13410 => '0',
		13411 => '1',
		13412 => '0',
		13413 => '1',
		13414 => '0',
		13415 => '1',
		13416 => '0',
		13417 => '1',
		13418 => '0',
		13419 => '1',
		13420 => '0',
		13421 => '1',
		13422 => '0',
		13423 => '1',
		13424 => '0',
		13425 => '1',
		13426 => '0',
		13427 => '1',
		13428 => '0',
		13429 => '1',
		13430 => '0',
		13431 => '1',
		13440 => '1',
		13441 => '0',
		13442 => '1',
		13443 => '0',
		13444 => '1',
		13445 => '0',
		13446 => '1',
		13447 => '0',
		13448 => '1',
		13449 => '0',
		13450 => '1',
		13451 => '0',
		13452 => '1',
		13453 => '0',
		13454 => '1',
		13455 => '0',
		13456 => '1',
		13457 => '0',
		13458 => '1',
		13459 => '0',
		13460 => '1',
		13461 => '0',
		13462 => '1',
		13463 => '0',
		13464 => '1',
		13465 => '0',
		13466 => '1',
		13467 => '0',
		13468 => '1',
		13469 => '0',
		13470 => '1',
		13471 => '0',
		13472 => '1',
		13473 => '0',
		13474 => '1',
		13475 => '0',
		13476 => '1',
		13477 => '0',
		13478 => '1',
		13479 => '0',
		13480 => '1',
		13481 => '0',
		13482 => '1',
		13483 => '0',
		13484 => '1',
		13485 => '0',
		13486 => '1',
		13487 => '0',
		13488 => '1',
		13489 => '0',
		13490 => '1',
		13491 => '0',
		13492 => '1',
		13493 => '0',
		13494 => '1',
		13495 => '0',
		13496 => '1',
		13497 => '0',
		13498 => '1',
		13499 => '0',
		13500 => '1',
		13501 => '0',
		13502 => '1',
		13503 => '0',
		13504 => '1',
		13505 => '0',
		13506 => '1',
		13507 => '0',
		13508 => '1',
		13509 => '0',
		13510 => '1',
		13511 => '0',
		13512 => '1',
		13513 => '0',
		13514 => '1',
		13515 => '0',
		13516 => '1',
		13517 => '0',
		13518 => '1',
		13519 => '0',
		13520 => '1',
		13521 => '0',
		13522 => '1',
		13523 => '0',
		13524 => '1',
		13525 => '0',
		13526 => '1',
		13527 => '0',
		13528 => '1',
		13529 => '0',
		13530 => '1',
		13531 => '0',
		13532 => '1',
		13533 => '0',
		13534 => '1',
		13535 => '0',
		13536 => '1',
		13537 => '0',
		13538 => '1',
		13539 => '0',
		13540 => '1',
		13541 => '0',
		13542 => '1',
		13543 => '0',
		13544 => '1',
		13545 => '0',
		13546 => '1',
		13547 => '0',
		13548 => '1',
		13549 => '0',
		13550 => '1',
		13551 => '0',
		13552 => '1',
		13553 => '0',
		13554 => '1',
		13555 => '0',
		13556 => '1',
		13557 => '0',
		13558 => '1',
		13559 => '0',
		13568 => '0',
		13569 => '1',
		13570 => '0',
		13571 => '1',
		13572 => '0',
		13573 => '1',
		13574 => '0',
		13575 => '1',
		13576 => '0',
		13577 => '1',
		13578 => '0',
		13579 => '1',
		13580 => '0',
		13581 => '1',
		13582 => '0',
		13583 => '1',
		13584 => '0',
		13585 => '1',
		13586 => '0',
		13587 => '1',
		13588 => '0',
		13589 => '1',
		13590 => '0',
		13591 => '1',
		13592 => '0',
		13593 => '1',
		13594 => '0',
		13595 => '1',
		13596 => '0',
		13597 => '1',
		13598 => '0',
		13599 => '1',
		13600 => '0',
		13601 => '1',
		13602 => '0',
		13603 => '1',
		13604 => '0',
		13605 => '1',
		13606 => '0',
		13607 => '1',
		13608 => '0',
		13609 => '1',
		13610 => '0',
		13611 => '1',
		13612 => '0',
		13613 => '1',
		13614 => '0',
		13615 => '1',
		13616 => '0',
		13617 => '1',
		13618 => '0',
		13619 => '1',
		13620 => '0',
		13621 => '1',
		13622 => '0',
		13623 => '1',
		13624 => '0',
		13625 => '1',
		13626 => '0',
		13627 => '1',
		13628 => '0',
		13629 => '1',
		13630 => '0',
		13631 => '1',
		13632 => '0',
		13633 => '1',
		13634 => '0',
		13635 => '1',
		13636 => '0',
		13637 => '1',
		13638 => '0',
		13639 => '1',
		13640 => '0',
		13641 => '1',
		13642 => '0',
		13643 => '1',
		13644 => '0',
		13645 => '1',
		13646 => '0',
		13647 => '1',
		13648 => '0',
		13649 => '1',
		13650 => '0',
		13651 => '1',
		13652 => '0',
		13653 => '1',
		13654 => '0',
		13655 => '1',
		13656 => '0',
		13657 => '1',
		13658 => '0',
		13659 => '1',
		13660 => '0',
		13661 => '1',
		13662 => '0',
		13663 => '1',
		13664 => '0',
		13665 => '1',
		13666 => '0',
		13667 => '1',
		13668 => '0',
		13669 => '1',
		13670 => '0',
		13671 => '1',
		13672 => '0',
		13673 => '1',
		13674 => '0',
		13675 => '1',
		13676 => '0',
		13677 => '1',
		13678 => '0',
		13679 => '1',
		13680 => '0',
		13681 => '1',
		13682 => '0',
		13683 => '1',
		13684 => '0',
		13685 => '1',
		13686 => '0',
		13687 => '1',
		13696 => '1',
		13697 => '0',
		13698 => '1',
		13699 => '0',
		13700 => '1',
		13701 => '0',
		13702 => '1',
		13703 => '0',
		13704 => '1',
		13705 => '0',
		13706 => '1',
		13707 => '0',
		13708 => '1',
		13709 => '0',
		13710 => '1',
		13711 => '0',
		13712 => '1',
		13713 => '0',
		13714 => '1',
		13715 => '0',
		13716 => '1',
		13717 => '0',
		13718 => '1',
		13719 => '0',
		13720 => '1',
		13721 => '0',
		13722 => '1',
		13723 => '0',
		13724 => '1',
		13725 => '0',
		13726 => '1',
		13727 => '0',
		13728 => '1',
		13729 => '0',
		13730 => '1',
		13731 => '0',
		13732 => '1',
		13733 => '0',
		13734 => '1',
		13735 => '0',
		13736 => '1',
		13737 => '0',
		13738 => '1',
		13739 => '0',
		13740 => '1',
		13741 => '0',
		13742 => '1',
		13743 => '0',
		13744 => '1',
		13745 => '0',
		13746 => '1',
		13747 => '0',
		13748 => '1',
		13749 => '0',
		13750 => '1',
		13751 => '0',
		13752 => '1',
		13753 => '0',
		13754 => '1',
		13755 => '0',
		13756 => '1',
		13757 => '0',
		13758 => '1',
		13759 => '0',
		13760 => '1',
		13761 => '0',
		13762 => '1',
		13763 => '0',
		13764 => '1',
		13765 => '0',
		13766 => '1',
		13767 => '0',
		13768 => '1',
		13769 => '0',
		13770 => '1',
		13771 => '0',
		13772 => '1',
		13773 => '0',
		13774 => '1',
		13775 => '0',
		13776 => '1',
		13777 => '0',
		13778 => '1',
		13779 => '0',
		13780 => '1',
		13781 => '0',
		13782 => '1',
		13783 => '0',
		13784 => '1',
		13785 => '0',
		13786 => '1',
		13787 => '0',
		13788 => '1',
		13789 => '0',
		13790 => '1',
		13791 => '0',
		13792 => '1',
		13793 => '0',
		13794 => '1',
		13795 => '0',
		13796 => '1',
		13797 => '0',
		13798 => '1',
		13799 => '0',
		13800 => '1',
		13801 => '0',
		13802 => '1',
		13803 => '0',
		13804 => '1',
		13805 => '0',
		13806 => '1',
		13807 => '0',
		13808 => '1',
		13809 => '0',
		13810 => '1',
		13811 => '0',
		13812 => '1',
		13813 => '0',
		13814 => '1',
		13815 => '0',
		13824 => '0',
		13825 => '1',
		13826 => '0',
		13827 => '1',
		13828 => '0',
		13829 => '1',
		13830 => '0',
		13831 => '1',
		13832 => '0',
		13833 => '1',
		13834 => '0',
		13835 => '1',
		13836 => '0',
		13837 => '1',
		13838 => '0',
		13839 => '1',
		13840 => '0',
		13841 => '1',
		13842 => '0',
		13843 => '1',
		13844 => '0',
		13845 => '1',
		13846 => '0',
		13847 => '1',
		13848 => '0',
		13849 => '1',
		13850 => '0',
		13851 => '1',
		13852 => '0',
		13853 => '1',
		13854 => '0',
		13855 => '1',
		13856 => '0',
		13857 => '1',
		13858 => '0',
		13859 => '1',
		13860 => '0',
		13861 => '1',
		13862 => '0',
		13863 => '1',
		13864 => '0',
		13865 => '1',
		13866 => '0',
		13867 => '1',
		13868 => '0',
		13869 => '1',
		13870 => '0',
		13871 => '1',
		13872 => '0',
		13873 => '1',
		13874 => '0',
		13875 => '1',
		13876 => '0',
		13877 => '1',
		13878 => '0',
		13879 => '1',
		13880 => '0',
		13881 => '1',
		13882 => '0',
		13883 => '1',
		13884 => '0',
		13885 => '1',
		13886 => '0',
		13887 => '1',
		13888 => '0',
		13889 => '1',
		13890 => '0',
		13891 => '1',
		13892 => '0',
		13893 => '1',
		13894 => '0',
		13895 => '1',
		13896 => '0',
		13897 => '1',
		13898 => '0',
		13899 => '1',
		13900 => '0',
		13901 => '1',
		13902 => '0',
		13903 => '1',
		13904 => '0',
		13905 => '1',
		13906 => '0',
		13907 => '1',
		13908 => '0',
		13909 => '1',
		13910 => '0',
		13911 => '1',
		13912 => '0',
		13913 => '1',
		13914 => '0',
		13915 => '1',
		13916 => '0',
		13917 => '1',
		13918 => '0',
		13919 => '1',
		13920 => '0',
		13921 => '1',
		13922 => '0',
		13923 => '1',
		13924 => '0',
		13925 => '1',
		13926 => '0',
		13927 => '1',
		13928 => '0',
		13929 => '1',
		13930 => '0',
		13931 => '1',
		13932 => '0',
		13933 => '1',
		13934 => '0',
		13935 => '1',
		13936 => '0',
		13937 => '1',
		13938 => '0',
		13939 => '1',
		13940 => '0',
		13941 => '1',
		13942 => '0',
		13943 => '1',
		13952 => '1',
		13953 => '0',
		13954 => '1',
		13955 => '0',
		13956 => '1',
		13957 => '0',
		13958 => '1',
		13959 => '0',
		13960 => '1',
		13961 => '0',
		13962 => '1',
		13963 => '0',
		13964 => '1',
		13965 => '0',
		13966 => '1',
		13967 => '0',
		13968 => '1',
		13969 => '0',
		13970 => '1',
		13971 => '0',
		13972 => '1',
		13973 => '0',
		13974 => '1',
		13975 => '0',
		13976 => '1',
		13977 => '0',
		13978 => '1',
		13979 => '0',
		13980 => '1',
		13981 => '0',
		13982 => '1',
		13983 => '0',
		13984 => '1',
		13985 => '0',
		13986 => '1',
		13987 => '0',
		13988 => '1',
		13989 => '0',
		13990 => '1',
		13991 => '0',
		13992 => '1',
		13993 => '0',
		13994 => '1',
		13995 => '0',
		13996 => '1',
		13997 => '0',
		13998 => '1',
		13999 => '0',
		14000 => '1',
		14001 => '0',
		14002 => '1',
		14003 => '0',
		14004 => '1',
		14005 => '0',
		14006 => '1',
		14007 => '0',
		14008 => '1',
		14009 => '0',
		14010 => '1',
		14011 => '0',
		14012 => '1',
		14013 => '0',
		14014 => '1',
		14015 => '0',
		14016 => '1',
		14017 => '0',
		14018 => '1',
		14019 => '0',
		14020 => '1',
		14021 => '0',
		14022 => '1',
		14023 => '0',
		14024 => '1',
		14025 => '0',
		14026 => '1',
		14027 => '0',
		14028 => '1',
		14029 => '0',
		14030 => '1',
		14031 => '0',
		14032 => '1',
		14033 => '0',
		14034 => '1',
		14035 => '0',
		14036 => '1',
		14037 => '0',
		14038 => '1',
		14039 => '0',
		14040 => '1',
		14041 => '0',
		14042 => '1',
		14043 => '0',
		14044 => '1',
		14045 => '0',
		14046 => '1',
		14047 => '0',
		14048 => '1',
		14049 => '0',
		14050 => '1',
		14051 => '0',
		14052 => '1',
		14053 => '0',
		14054 => '1',
		14055 => '0',
		14056 => '1',
		14057 => '0',
		14058 => '1',
		14059 => '0',
		14060 => '1',
		14061 => '0',
		14062 => '1',
		14063 => '0',
		14064 => '1',
		14065 => '0',
		14066 => '1',
		14067 => '0',
		14068 => '1',
		14069 => '0',
		14070 => '1',
		14071 => '0',
		14080 => '0',
		14081 => '1',
		14082 => '0',
		14083 => '1',
		14084 => '0',
		14085 => '1',
		14086 => '0',
		14087 => '1',
		14088 => '0',
		14089 => '1',
		14090 => '0',
		14091 => '1',
		14092 => '0',
		14093 => '1',
		14094 => '0',
		14095 => '1',
		14096 => '0',
		14097 => '1',
		14098 => '0',
		14099 => '1',
		14100 => '0',
		14101 => '1',
		14102 => '0',
		14103 => '1',
		14104 => '0',
		14105 => '1',
		14106 => '0',
		14107 => '1',
		14108 => '0',
		14109 => '1',
		14110 => '0',
		14111 => '1',
		14112 => '0',
		14113 => '1',
		14114 => '0',
		14115 => '1',
		14116 => '0',
		14117 => '1',
		14118 => '0',
		14119 => '1',
		14120 => '0',
		14121 => '1',
		14122 => '0',
		14123 => '1',
		14124 => '0',
		14125 => '1',
		14126 => '0',
		14127 => '1',
		14128 => '0',
		14129 => '1',
		14130 => '0',
		14131 => '1',
		14132 => '0',
		14133 => '1',
		14134 => '0',
		14135 => '1',
		14136 => '0',
		14137 => '1',
		14138 => '0',
		14139 => '1',
		14140 => '0',
		14141 => '1',
		14142 => '0',
		14143 => '1',
		14144 => '0',
		14145 => '1',
		14146 => '0',
		14147 => '1',
		14148 => '0',
		14149 => '1',
		14150 => '0',
		14151 => '1',
		14152 => '0',
		14153 => '1',
		14154 => '0',
		14155 => '1',
		14156 => '0',
		14157 => '1',
		14158 => '0',
		14159 => '1',
		14160 => '0',
		14161 => '1',
		14162 => '0',
		14163 => '1',
		14164 => '0',
		14165 => '1',
		14166 => '0',
		14167 => '1',
		14168 => '0',
		14169 => '1',
		14170 => '0',
		14171 => '1',
		14172 => '0',
		14173 => '1',
		14174 => '0',
		14175 => '1',
		14176 => '0',
		14177 => '1',
		14178 => '0',
		14179 => '1',
		14180 => '0',
		14181 => '1',
		14182 => '0',
		14183 => '1',
		14184 => '0',
		14185 => '1',
		14186 => '0',
		14187 => '1',
		14188 => '0',
		14189 => '1',
		14190 => '0',
		14191 => '1',
		14192 => '0',
		14193 => '1',
		14194 => '0',
		14195 => '1',
		14196 => '0',
		14197 => '1',
		14198 => '0',
		14199 => '1',
		14208 => '1',
		14209 => '0',
		14210 => '1',
		14211 => '0',
		14212 => '1',
		14213 => '0',
		14214 => '1',
		14215 => '0',
		14216 => '1',
		14217 => '0',
		14218 => '1',
		14219 => '0',
		14220 => '1',
		14221 => '0',
		14222 => '1',
		14223 => '0',
		14224 => '1',
		14225 => '0',
		14226 => '1',
		14227 => '0',
		14228 => '1',
		14229 => '0',
		14230 => '1',
		14231 => '0',
		14232 => '1',
		14233 => '0',
		14234 => '1',
		14235 => '0',
		14236 => '1',
		14237 => '0',
		14238 => '1',
		14239 => '0',
		14240 => '1',
		14241 => '0',
		14242 => '1',
		14243 => '0',
		14244 => '1',
		14245 => '0',
		14246 => '1',
		14247 => '0',
		14248 => '1',
		14249 => '0',
		14250 => '1',
		14251 => '0',
		14252 => '1',
		14253 => '0',
		14254 => '1',
		14255 => '0',
		14256 => '1',
		14257 => '0',
		14258 => '1',
		14259 => '0',
		14260 => '1',
		14261 => '0',
		14262 => '1',
		14263 => '0',
		14264 => '1',
		14265 => '0',
		14266 => '1',
		14267 => '0',
		14268 => '1',
		14269 => '0',
		14270 => '1',
		14271 => '0',
		14272 => '1',
		14273 => '0',
		14274 => '1',
		14275 => '0',
		14276 => '1',
		14277 => '0',
		14278 => '1',
		14279 => '0',
		14280 => '1',
		14281 => '0',
		14282 => '1',
		14283 => '0',
		14284 => '1',
		14285 => '0',
		14286 => '1',
		14287 => '0',
		14288 => '1',
		14289 => '0',
		14290 => '1',
		14291 => '0',
		14292 => '1',
		14293 => '0',
		14294 => '1',
		14295 => '0',
		14296 => '1',
		14297 => '0',
		14298 => '1',
		14299 => '0',
		14300 => '1',
		14301 => '0',
		14302 => '1',
		14303 => '0',
		14304 => '1',
		14305 => '0',
		14306 => '1',
		14307 => '0',
		14308 => '1',
		14309 => '0',
		14310 => '1',
		14311 => '0',
		14312 => '1',
		14313 => '0',
		14314 => '1',
		14315 => '0',
		14316 => '1',
		14317 => '0',
		14318 => '1',
		14319 => '0',
		14320 => '1',
		14321 => '0',
		14322 => '1',
		14323 => '0',
		14324 => '1',
		14325 => '0',
		14326 => '1',
		14327 => '0',
		14336 => '0',
		14337 => '1',
		14338 => '0',
		14339 => '1',
		14340 => '0',
		14341 => '1',
		14342 => '0',
		14343 => '1',
		14344 => '0',
		14345 => '1',
		14346 => '0',
		14347 => '1',
		14348 => '0',
		14349 => '1',
		14350 => '0',
		14351 => '1',
		14352 => '0',
		14353 => '1',
		14354 => '0',
		14355 => '1',
		14356 => '0',
		14357 => '1',
		14358 => '0',
		14359 => '1',
		14360 => '0',
		14361 => '1',
		14362 => '0',
		14363 => '1',
		14364 => '0',
		14365 => '1',
		14366 => '0',
		14367 => '1',
		14368 => '0',
		14369 => '1',
		14370 => '0',
		14371 => '1',
		14372 => '0',
		14373 => '1',
		14374 => '0',
		14375 => '1',
		14376 => '0',
		14377 => '1',
		14378 => '0',
		14379 => '1',
		14380 => '0',
		14381 => '1',
		14382 => '0',
		14383 => '1',
		14384 => '0',
		14385 => '1',
		14386 => '0',
		14387 => '1',
		14388 => '0',
		14389 => '1',
		14390 => '0',
		14391 => '1',
		14392 => '0',
		14393 => '1',
		14394 => '0',
		14395 => '1',
		14396 => '0',
		14397 => '1',
		14398 => '0',
		14399 => '1',
		14400 => '0',
		14401 => '1',
		14402 => '0',
		14403 => '1',
		14404 => '0',
		14405 => '1',
		14406 => '0',
		14407 => '1',
		14408 => '0',
		14409 => '1',
		14410 => '0',
		14411 => '1',
		14412 => '0',
		14413 => '1',
		14414 => '0',
		14415 => '1',
		14416 => '0',
		14417 => '1',
		14418 => '0',
		14419 => '1',
		14420 => '0',
		14421 => '1',
		14422 => '0',
		14423 => '1',
		14424 => '0',
		14425 => '1',
		14426 => '0',
		14427 => '1',
		14428 => '0',
		14429 => '1',
		14430 => '0',
		14431 => '1',
		14432 => '0',
		14433 => '1',
		14434 => '0',
		14435 => '1',
		14436 => '0',
		14437 => '1',
		14438 => '0',
		14439 => '1',
		14440 => '0',
		14441 => '1',
		14442 => '0',
		14443 => '1',
		14444 => '0',
		14445 => '1',
		14446 => '0',
		14447 => '1',
		14448 => '0',
		14449 => '1',
		14450 => '0',
		14451 => '1',
		14452 => '0',
		14453 => '1',
		14454 => '0',
		14455 => '1',
		14464 => '1',
		14465 => '0',
		14466 => '1',
		14467 => '0',
		14468 => '1',
		14469 => '0',
		14470 => '1',
		14471 => '0',
		14472 => '1',
		14473 => '0',
		14474 => '1',
		14475 => '0',
		14476 => '1',
		14477 => '0',
		14478 => '1',
		14479 => '0',
		14480 => '1',
		14481 => '0',
		14482 => '1',
		14483 => '0',
		14484 => '1',
		14485 => '0',
		14486 => '1',
		14487 => '0',
		14488 => '1',
		14489 => '0',
		14490 => '1',
		14491 => '0',
		14492 => '1',
		14493 => '0',
		14494 => '1',
		14495 => '0',
		14496 => '1',
		14497 => '0',
		14498 => '1',
		14499 => '0',
		14500 => '1',
		14501 => '0',
		14502 => '1',
		14503 => '0',
		14504 => '1',
		14505 => '0',
		14506 => '1',
		14507 => '0',
		14508 => '1',
		14509 => '0',
		14510 => '1',
		14511 => '0',
		14512 => '1',
		14513 => '0',
		14514 => '1',
		14515 => '0',
		14516 => '1',
		14517 => '0',
		14518 => '1',
		14519 => '0',
		14520 => '1',
		14521 => '0',
		14522 => '1',
		14523 => '0',
		14524 => '1',
		14525 => '0',
		14526 => '1',
		14527 => '0',
		14528 => '1',
		14529 => '0',
		14530 => '1',
		14531 => '0',
		14532 => '1',
		14533 => '0',
		14534 => '1',
		14535 => '0',
		14536 => '1',
		14537 => '0',
		14538 => '1',
		14539 => '0',
		14540 => '1',
		14541 => '0',
		14542 => '1',
		14543 => '0',
		14544 => '1',
		14545 => '0',
		14546 => '1',
		14547 => '0',
		14548 => '1',
		14549 => '0',
		14550 => '1',
		14551 => '0',
		14552 => '1',
		14553 => '0',
		14554 => '1',
		14555 => '0',
		14556 => '1',
		14557 => '0',
		14558 => '1',
		14559 => '0',
		14560 => '1',
		14561 => '0',
		14562 => '1',
		14563 => '0',
		14564 => '1',
		14565 => '0',
		14566 => '1',
		14567 => '0',
		14568 => '1',
		14569 => '0',
		14570 => '1',
		14571 => '0',
		14572 => '1',
		14573 => '0',
		14574 => '1',
		14575 => '0',
		14576 => '1',
		14577 => '0',
		14578 => '1',
		14579 => '0',
		14580 => '1',
		14581 => '0',
		14582 => '1',
		14583 => '0',
		14592 => '0',
		14593 => '1',
		14594 => '0',
		14595 => '1',
		14596 => '0',
		14597 => '1',
		14598 => '0',
		14599 => '1',
		14600 => '0',
		14601 => '1',
		14602 => '0',
		14603 => '1',
		14604 => '0',
		14605 => '1',
		14606 => '0',
		14607 => '1',
		14608 => '0',
		14609 => '1',
		14610 => '0',
		14611 => '1',
		14612 => '0',
		14613 => '1',
		14614 => '0',
		14615 => '1',
		14616 => '0',
		14617 => '1',
		14618 => '0',
		14619 => '1',
		14620 => '0',
		14621 => '1',
		14622 => '0',
		14623 => '1',
		14624 => '0',
		14625 => '1',
		14626 => '0',
		14627 => '1',
		14628 => '0',
		14629 => '1',
		14630 => '0',
		14631 => '1',
		14632 => '0',
		14633 => '1',
		14634 => '0',
		14635 => '1',
		14636 => '0',
		14637 => '1',
		14638 => '0',
		14639 => '1',
		14640 => '0',
		14641 => '1',
		14642 => '0',
		14643 => '1',
		14644 => '0',
		14645 => '1',
		14646 => '0',
		14647 => '1',
		14648 => '0',
		14649 => '1',
		14650 => '0',
		14651 => '1',
		14652 => '0',
		14653 => '1',
		14654 => '0',
		14655 => '1',
		14656 => '0',
		14657 => '1',
		14658 => '0',
		14659 => '1',
		14660 => '0',
		14661 => '1',
		14662 => '0',
		14663 => '1',
		14664 => '0',
		14665 => '1',
		14666 => '0',
		14667 => '1',
		14668 => '0',
		14669 => '1',
		14670 => '0',
		14671 => '1',
		14672 => '0',
		14673 => '1',
		14674 => '0',
		14675 => '1',
		14676 => '0',
		14677 => '1',
		14678 => '0',
		14679 => '1',
		14680 => '0',
		14681 => '1',
		14682 => '0',
		14683 => '1',
		14684 => '0',
		14685 => '1',
		14686 => '0',
		14687 => '1',
		14688 => '0',
		14689 => '1',
		14690 => '0',
		14691 => '1',
		14692 => '0',
		14693 => '1',
		14694 => '0',
		14695 => '1',
		14696 => '0',
		14697 => '1',
		14698 => '0',
		14699 => '1',
		14700 => '0',
		14701 => '1',
		14702 => '0',
		14703 => '1',
		14704 => '0',
		14705 => '1',
		14706 => '0',
		14707 => '1',
		14708 => '0',
		14709 => '1',
		14710 => '0',
		14711 => '1',
		14720 => '1',
		14721 => '0',
		14722 => '1',
		14723 => '0',
		14724 => '1',
		14725 => '0',
		14726 => '1',
		14727 => '0',
		14728 => '1',
		14729 => '0',
		14730 => '1',
		14731 => '0',
		14732 => '1',
		14733 => '0',
		14734 => '1',
		14735 => '0',
		14736 => '1',
		14737 => '0',
		14738 => '1',
		14739 => '0',
		14740 => '1',
		14741 => '0',
		14742 => '1',
		14743 => '0',
		14744 => '1',
		14745 => '0',
		14746 => '1',
		14747 => '0',
		14748 => '1',
		14749 => '0',
		14750 => '1',
		14751 => '0',
		14752 => '1',
		14753 => '0',
		14754 => '1',
		14755 => '0',
		14756 => '1',
		14757 => '0',
		14758 => '1',
		14759 => '0',
		14760 => '1',
		14761 => '0',
		14762 => '1',
		14763 => '0',
		14764 => '1',
		14765 => '0',
		14766 => '1',
		14767 => '0',
		14768 => '1',
		14769 => '0',
		14770 => '1',
		14771 => '0',
		14772 => '1',
		14773 => '0',
		14774 => '1',
		14775 => '0',
		14776 => '1',
		14777 => '0',
		14778 => '1',
		14779 => '0',
		14780 => '1',
		14781 => '0',
		14782 => '1',
		14783 => '0',
		14784 => '1',
		14785 => '0',
		14786 => '1',
		14787 => '0',
		14788 => '1',
		14789 => '0',
		14790 => '1',
		14791 => '0',
		14792 => '1',
		14793 => '0',
		14794 => '1',
		14795 => '0',
		14796 => '1',
		14797 => '0',
		14798 => '1',
		14799 => '0',
		14800 => '1',
		14801 => '0',
		14802 => '1',
		14803 => '0',
		14804 => '1',
		14805 => '0',
		14806 => '1',
		14807 => '0',
		14808 => '1',
		14809 => '0',
		14810 => '1',
		14811 => '0',
		14812 => '1',
		14813 => '0',
		14814 => '1',
		14815 => '0',
		14816 => '1',
		14817 => '0',
		14818 => '1',
		14819 => '0',
		14820 => '1',
		14821 => '0',
		14822 => '1',
		14823 => '0',
		14824 => '1',
		14825 => '0',
		14826 => '1',
		14827 => '0',
		14828 => '1',
		14829 => '0',
		14830 => '1',
		14831 => '0',
		14832 => '1',
		14833 => '0',
		14834 => '1',
		14835 => '0',
		14836 => '1',
		14837 => '0',
		14838 => '1',
		14839 => '0',
		14848 => '0',
		14849 => '1',
		14850 => '0',
		14851 => '1',
		14852 => '0',
		14853 => '1',
		14854 => '0',
		14855 => '1',
		14856 => '0',
		14857 => '1',
		14858 => '0',
		14859 => '1',
		14860 => '0',
		14861 => '1',
		14862 => '0',
		14863 => '1',
		14864 => '0',
		14865 => '1',
		14866 => '0',
		14867 => '1',
		14868 => '0',
		14869 => '1',
		14870 => '0',
		14871 => '1',
		14872 => '0',
		14873 => '1',
		14874 => '0',
		14875 => '1',
		14876 => '0',
		14877 => '1',
		14878 => '0',
		14879 => '1',
		14880 => '0',
		14881 => '1',
		14882 => '0',
		14883 => '1',
		14884 => '0',
		14885 => '1',
		14886 => '0',
		14887 => '1',
		14888 => '0',
		14889 => '1',
		14890 => '0',
		14891 => '1',
		14892 => '0',
		14893 => '1',
		14894 => '0',
		14895 => '1',
		14896 => '0',
		14897 => '1',
		14898 => '0',
		14899 => '1',
		14900 => '0',
		14901 => '1',
		14902 => '0',
		14903 => '1',
		14904 => '0',
		14905 => '1',
		14906 => '0',
		14907 => '1',
		14908 => '0',
		14909 => '1',
		14910 => '0',
		14911 => '1',
		14912 => '0',
		14913 => '1',
		14914 => '0',
		14915 => '1',
		14916 => '0',
		14917 => '1',
		14918 => '0',
		14919 => '1',
		14920 => '0',
		14921 => '1',
		14922 => '0',
		14923 => '1',
		14924 => '0',
		14925 => '1',
		14926 => '0',
		14927 => '1',
		14928 => '0',
		14929 => '1',
		14930 => '0',
		14931 => '1',
		14932 => '0',
		14933 => '1',
		14934 => '0',
		14935 => '1',
		14936 => '0',
		14937 => '1',
		14938 => '0',
		14939 => '1',
		14940 => '0',
		14941 => '1',
		14942 => '0',
		14943 => '1',
		14944 => '0',
		14945 => '1',
		14946 => '0',
		14947 => '1',
		14948 => '0',
		14949 => '1',
		14950 => '0',
		14951 => '1',
		14952 => '0',
		14953 => '1',
		14954 => '0',
		14955 => '1',
		14956 => '0',
		14957 => '1',
		14958 => '0',
		14959 => '1',
		14960 => '0',
		14961 => '1',
		14962 => '0',
		14963 => '1',
		14964 => '0',
		14965 => '1',
		14966 => '0',
		14967 => '1',
		14976 => '1',
		14977 => '0',
		14978 => '1',
		14979 => '0',
		14980 => '1',
		14981 => '0',
		14982 => '1',
		14983 => '0',
		14984 => '1',
		14985 => '0',
		14986 => '1',
		14987 => '0',
		14988 => '1',
		14989 => '0',
		14990 => '1',
		14991 => '0',
		14992 => '1',
		14993 => '0',
		14994 => '1',
		14995 => '0',
		14996 => '1',
		14997 => '0',
		14998 => '1',
		14999 => '0',
		15000 => '1',
		15001 => '0',
		15002 => '1',
		15003 => '0',
		15004 => '1',
		15005 => '0',
		15006 => '1',
		15007 => '0',
		15008 => '1',
		15009 => '0',
		15010 => '1',
		15011 => '0',
		15012 => '1',
		15013 => '0',
		15014 => '1',
		15015 => '0',
		15016 => '1',
		15017 => '0',
		15018 => '1',
		15019 => '0',
		15020 => '1',
		15021 => '0',
		15022 => '1',
		15023 => '0',
		15024 => '1',
		15025 => '0',
		15026 => '1',
		15027 => '0',
		15028 => '1',
		15029 => '0',
		15030 => '1',
		15031 => '0',
		15032 => '1',
		15033 => '0',
		15034 => '1',
		15035 => '0',
		15036 => '1',
		15037 => '0',
		15038 => '1',
		15039 => '0',
		15040 => '1',
		15041 => '0',
		15042 => '1',
		15043 => '0',
		15044 => '1',
		15045 => '0',
		15046 => '1',
		15047 => '0',
		15048 => '1',
		15049 => '0',
		15050 => '1',
		15051 => '0',
		15052 => '1',
		15053 => '0',
		15054 => '1',
		15055 => '0',
		15056 => '1',
		15057 => '0',
		15058 => '1',
		15059 => '0',
		15060 => '1',
		15061 => '0',
		15062 => '1',
		15063 => '0',
		15064 => '1',
		15065 => '0',
		15066 => '1',
		15067 => '0',
		15068 => '1',
		15069 => '0',
		15070 => '1',
		15071 => '0',
		15072 => '1',
		15073 => '0',
		15074 => '1',
		15075 => '0',
		15076 => '1',
		15077 => '0',
		15078 => '1',
		15079 => '0',
		15080 => '1',
		15081 => '0',
		15082 => '1',
		15083 => '0',
		15084 => '1',
		15085 => '0',
		15086 => '1',
		15087 => '0',
		15088 => '1',
		15089 => '0',
		15090 => '1',
		15091 => '0',
		15092 => '1',
		15093 => '0',
		15094 => '1',
		15095 => '0',
		15104 => '0',
		15105 => '1',
		15106 => '0',
		15107 => '1',
		15108 => '0',
		15109 => '1',
		15110 => '0',
		15111 => '1',
		15112 => '0',
		15113 => '1',
		15114 => '0',
		15115 => '1',
		15116 => '0',
		15117 => '1',
		15118 => '0',
		15119 => '1',
		15120 => '0',
		15121 => '1',
		15122 => '0',
		15123 => '1',
		15124 => '0',
		15125 => '1',
		15126 => '0',
		15127 => '1',
		15128 => '0',
		15129 => '1',
		15130 => '0',
		15131 => '1',
		15132 => '0',
		15133 => '1',
		15134 => '0',
		15135 => '1',
		15136 => '0',
		15137 => '1',
		15138 => '0',
		15139 => '1',
		15140 => '0',
		15141 => '1',
		15142 => '0',
		15143 => '1',
		15144 => '0',
		15145 => '1',
		15146 => '0',
		15147 => '1',
		15148 => '0',
		15149 => '1',
		15150 => '0',
		15151 => '1',
		15152 => '0',
		15153 => '1',
		15154 => '0',
		15155 => '1',
		15156 => '0',
		15157 => '1',
		15158 => '0',
		15159 => '1',
		15160 => '0',
		15161 => '1',
		15162 => '0',
		15163 => '1',
		15164 => '0',
		15165 => '1',
		15166 => '0',
		15167 => '1',
		15168 => '0',
		15169 => '1',
		15170 => '0',
		15171 => '1',
		15172 => '0',
		15173 => '1',
		15174 => '0',
		15175 => '1',
		15176 => '0',
		15177 => '1',
		15178 => '0',
		15179 => '1',
		15180 => '0',
		15181 => '1',
		15182 => '0',
		15183 => '1',
		15184 => '0',
		15185 => '1',
		15186 => '0',
		15187 => '1',
		15188 => '0',
		15189 => '1',
		15190 => '0',
		15191 => '1',
		15192 => '0',
		15193 => '1',
		15194 => '0',
		15195 => '1',
		15196 => '0',
		15197 => '1',
		15198 => '0',
		15199 => '1',
		15200 => '0',
		15201 => '1',
		15202 => '0',
		15203 => '1',
		15204 => '0',
		15205 => '1',
		15206 => '0',
		15207 => '1',
		15208 => '0',
		15209 => '1',
		15210 => '0',
		15211 => '1',
		15212 => '0',
		15213 => '1',
		15214 => '0',
		15215 => '1',
		15216 => '0',
		15217 => '1',
		15218 => '0',
		15219 => '1',
		15220 => '0',
		15221 => '1',
		15222 => '0',
		15223 => '1',
		15232 => '1',
		15233 => '0',
		15234 => '1',
		15235 => '0',
		15236 => '1',
		15237 => '0',
		15238 => '1',
		15239 => '0',
		15240 => '1',
		15241 => '0',
		15242 => '1',
		15243 => '0',
		15244 => '1',
		15245 => '0',
		15246 => '1',
		15247 => '0',
		15248 => '1',
		15249 => '0',
		15250 => '1',
		15251 => '0',
		15252 => '1',
		15253 => '0',
		15254 => '1',
		15255 => '0',
		15256 => '1',
		15257 => '0',
		15258 => '1',
		15259 => '0',
		15260 => '1',
		15261 => '0',
		15262 => '1',
		15263 => '0',
		15264 => '1',
		15265 => '0',
		15266 => '1',
		15267 => '0',
		15268 => '1',
		15269 => '0',
		15270 => '1',
		15271 => '0',
		15272 => '1',
		15273 => '0',
		15274 => '1',
		15275 => '0',
		15276 => '1',
		15277 => '0',
		15278 => '1',
		15279 => '0',
		15280 => '1',
		15281 => '0',
		15282 => '1',
		15283 => '0',
		15284 => '1',
		15285 => '0',
		15286 => '1',
		15287 => '0',
		15288 => '1',
		15289 => '0',
		15290 => '1',
		15291 => '0',
		15292 => '1',
		15293 => '0',
		15294 => '1',
		15295 => '0',
		15296 => '1',
		15297 => '0',
		15298 => '1',
		15299 => '0',
		15300 => '1',
		15301 => '0',
		15302 => '1',
		15303 => '0',
		15304 => '1',
		15305 => '0',
		15306 => '1',
		15307 => '0',
		15308 => '1',
		15309 => '0',
		15310 => '1',
		15311 => '0',
		15312 => '1',
		15313 => '0',
		15314 => '1',
		15315 => '0',
		15316 => '1',
		15317 => '0',
		15318 => '1',
		15319 => '0',
		15320 => '1',
		15321 => '0',
		15322 => '1',
		15323 => '0',
		15324 => '1',
		15325 => '0',
		15326 => '1',
		15327 => '0',
		15328 => '1',
		15329 => '0',
		15330 => '1',
		15331 => '0',
		15332 => '1',
		15333 => '0',
		15334 => '1',
		15335 => '0',
		15336 => '1',
		15337 => '0',
		15338 => '1',
		15339 => '0',
		15340 => '1',
		15341 => '0',
		15342 => '1',
		15343 => '0',
		15344 => '1',
		15345 => '0',
		15346 => '1',
		15347 => '0',
		15348 => '1',
		15349 => '0',
		15350 => '1',
		15351 => '0',

	others => '0'
);

begin
	
	-- process ROM
	process (CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (EN = '1') then
				DATA <= ROM(to_integer(unsigned(ADDR)));
			end if;
		end if;
	end process;
	
end Behavioral;

