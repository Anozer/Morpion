library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM_vide is
	port (CLK : in std_logic;
		  EN : in std_logic;
		  ADDR : in std_logic_vector(11 downto 0);
		  DATA : out std_logic_vector(7 downto 0));
end ROM_vide;

architecture Behavioral of ROM_vide is

type zone_memoire is array ((2**12)-1 downto 0) of std_logic_vector (7 downto 0);
constant ROM: zone_memoire := (
	0 => "00000000",
	1 => "00000000",
	2 => "00000000",
	3 => "00000000",
	4 => "00000000",
	5 => "00000000",
	6 => "00000000",
	7 => "00000000",
	8 => "00000000",
	9 => "00000000",
	10 => "00000000",
	11 => "00000000",
	12 => "00000000",
	13 => "00000000",
	14 => "00000000",
	15 => "00000000",
	16 => "00000000",
	17 => "00000000",
	18 => "00000000",
	19 => "00000000",
	20 => "00000000",
	21 => "00000000",
	22 => "00000000",
	23 => "00000000",
	24 => "00000000",
	25 => "00000000",
	26 => "00000000",
	27 => "00000000",
	28 => "00000000",
	29 => "00000000",
	30 => "00000000",
	31 => "00000000",
	32 => "00000000",
	33 => "00000000",
	34 => "00000000",
	35 => "00000000",
	36 => "00000000",
	37 => "00000000",
	38 => "00000000",
	39 => "00000000",
	40 => "00000000",
	41 => "00000000",
	42 => "00000000",
	43 => "00000000",
	44 => "00000000",
	45 => "00000000",
	46 => "00000000",
	47 => "00000000",
	48 => "00000000",
	49 => "00000000",
	50 => "00000000",
	51 => "00000000",
	52 => "00000000",
	53 => "00000000",
	54 => "00000000",
	55 => "00000000",
	56 => "00000000",
	57 => "00000000",
	58 => "00000000",
	59 => "00000000",
	64 => "00000000",
	65 => "00000000",
	66 => "00000000",
	67 => "00000000",
	68 => "00000000",
	69 => "00000000",
	70 => "00000000",
	71 => "00000000",
	72 => "00000000",
	73 => "00000000",
	74 => "00000000",
	75 => "00000000",
	76 => "00000000",
	77 => "00000000",
	78 => "00000000",
	79 => "00000000",
	80 => "00000000",
	81 => "00000000",
	82 => "00000000",
	83 => "00000000",
	84 => "00000000",
	85 => "00000000",
	86 => "00000000",
	87 => "00000000",
	88 => "00000000",
	89 => "00000000",
	90 => "00000000",
	91 => "00000000",
	92 => "00000000",
	93 => "00000000",
	94 => "00000000",
	95 => "00000000",
	96 => "00000000",
	97 => "00000000",
	98 => "00000000",
	99 => "00000000",
	100 => "00000000",
	101 => "00000000",
	102 => "00000000",
	103 => "00000000",
	104 => "00000000",
	105 => "00000000",
	106 => "00000000",
	107 => "00000000",
	108 => "00000000",
	109 => "00000000",
	110 => "00000000",
	111 => "00000000",
	112 => "00000000",
	113 => "00000000",
	114 => "00000000",
	115 => "00000000",
	116 => "00000000",
	117 => "00000000",
	118 => "00000000",
	119 => "00000000",
	120 => "00000000",
	121 => "00000000",
	122 => "00000000",
	123 => "00000000",
	128 => "00000000",
	129 => "00000000",
	130 => "00000000",
	131 => "00000000",
	132 => "00000000",
	133 => "00000000",
	134 => "00000000",
	135 => "00000000",
	136 => "00000000",
	137 => "00000000",
	138 => "00000000",
	139 => "00000000",
	140 => "00000000",
	141 => "00000000",
	142 => "00000000",
	143 => "00000000",
	144 => "00000000",
	145 => "00000000",
	146 => "00000000",
	147 => "00000000",
	148 => "00000000",
	149 => "00000000",
	150 => "00000000",
	151 => "00000000",
	152 => "00000000",
	153 => "00000000",
	154 => "00000000",
	155 => "00000000",
	156 => "00000000",
	157 => "00000000",
	158 => "00000000",
	159 => "00000000",
	160 => "00000000",
	161 => "00000000",
	162 => "00000000",
	163 => "00000000",
	164 => "00000000",
	165 => "00000000",
	166 => "00000000",
	167 => "00000000",
	168 => "00000000",
	169 => "00000000",
	170 => "00000000",
	171 => "00000000",
	172 => "00000000",
	173 => "00000000",
	174 => "00000000",
	175 => "00000000",
	176 => "00000000",
	177 => "00000000",
	178 => "00000000",
	179 => "00000000",
	180 => "00000000",
	181 => "00000000",
	182 => "00000000",
	183 => "00000000",
	184 => "00000000",
	185 => "00000000",
	186 => "00000000",
	187 => "00000000",
	192 => "00000000",
	193 => "00000000",
	194 => "00000000",
	195 => "00000000",
	196 => "00000000",
	197 => "00000000",
	198 => "00000000",
	199 => "00000000",
	200 => "00000000",
	201 => "00000000",
	202 => "00000000",
	203 => "00000000",
	204 => "00000000",
	205 => "00000000",
	206 => "00000000",
	207 => "00000000",
	208 => "00000000",
	209 => "00000000",
	210 => "00000000",
	211 => "00000000",
	212 => "00000000",
	213 => "00000000",
	214 => "00000000",
	215 => "00000000",
	216 => "00000000",
	217 => "00000000",
	218 => "00000000",
	219 => "00000000",
	220 => "00000000",
	221 => "00000000",
	222 => "00000000",
	223 => "00000000",
	224 => "00000000",
	225 => "00000000",
	226 => "00000000",
	227 => "00000000",
	228 => "00000000",
	229 => "00000000",
	230 => "00000000",
	231 => "00000000",
	232 => "00000000",
	233 => "00000000",
	234 => "00000000",
	235 => "00000000",
	236 => "00000000",
	237 => "00000000",
	238 => "00000000",
	239 => "00000000",
	240 => "00000000",
	241 => "00000000",
	242 => "00000000",
	243 => "00000000",
	244 => "00000000",
	245 => "00000000",
	246 => "00000000",
	247 => "00000000",
	248 => "00000000",
	249 => "00000000",
	250 => "00000000",
	251 => "00000000",
	256 => "00000000",
	257 => "00000000",
	258 => "00000000",
	259 => "00000000",
	260 => "00000000",
	261 => "00000000",
	262 => "00000000",
	263 => "00000000",
	264 => "00000000",
	265 => "00000000",
	266 => "00000000",
	267 => "00000000",
	268 => "00000000",
	269 => "00000000",
	270 => "00000000",
	271 => "00000000",
	272 => "00000000",
	273 => "00000000",
	274 => "00000000",
	275 => "00000000",
	276 => "00000000",
	277 => "00000000",
	278 => "00000000",
	279 => "00000000",
	280 => "00000000",
	281 => "00000000",
	282 => "00000000",
	283 => "00000000",
	284 => "00000000",
	285 => "00000000",
	286 => "00000000",
	287 => "00000000",
	288 => "00000000",
	289 => "00000000",
	290 => "00000000",
	291 => "00000000",
	292 => "00000000",
	293 => "00000000",
	294 => "00000000",
	295 => "00000000",
	296 => "00000000",
	297 => "00000000",
	298 => "00000000",
	299 => "00000000",
	300 => "00000000",
	301 => "00000000",
	302 => "00000000",
	303 => "00000000",
	304 => "00000000",
	305 => "00000000",
	306 => "00000000",
	307 => "00000000",
	308 => "00000000",
	309 => "00000000",
	310 => "00000000",
	311 => "00000000",
	312 => "00000000",
	313 => "00000000",
	314 => "00000000",
	315 => "00000000",
	320 => "00000000",
	321 => "00000000",
	322 => "00000000",
	323 => "00000000",
	324 => "00000000",
	325 => "00000000",
	326 => "00000000",
	327 => "00000000",
	328 => "00000000",
	329 => "00000000",
	330 => "00000000",
	331 => "00000000",
	332 => "00000000",
	333 => "00000000",
	334 => "00000000",
	335 => "00000000",
	336 => "00000000",
	337 => "00000000",
	338 => "00000000",
	339 => "00000000",
	340 => "00000000",
	341 => "00000000",
	342 => "00000000",
	343 => "00000000",
	344 => "00000000",
	345 => "00000000",
	346 => "00000000",
	347 => "00000000",
	348 => "00000000",
	349 => "00000000",
	350 => "00000000",
	351 => "00000000",
	352 => "00000000",
	353 => "00000000",
	354 => "00000000",
	355 => "00000000",
	356 => "00000000",
	357 => "00000000",
	358 => "00000000",
	359 => "00000000",
	360 => "00000000",
	361 => "00000000",
	362 => "00000000",
	363 => "00000000",
	364 => "00000000",
	365 => "00000000",
	366 => "00000000",
	367 => "00000000",
	368 => "00000000",
	369 => "00000000",
	370 => "00000000",
	371 => "00000000",
	372 => "00000000",
	373 => "00000000",
	374 => "00000000",
	375 => "00000000",
	376 => "00000000",
	377 => "00000000",
	378 => "00000000",
	379 => "00000000",
	384 => "00000000",
	385 => "00000000",
	386 => "00000000",
	387 => "00000000",
	388 => "00000000",
	389 => "00000000",
	390 => "00000000",
	391 => "00000000",
	392 => "00000000",
	393 => "00000000",
	394 => "00000000",
	395 => "00000000",
	396 => "00000000",
	397 => "00000000",
	398 => "00000000",
	399 => "00000000",
	400 => "00000000",
	401 => "00000000",
	402 => "00000000",
	403 => "00000000",
	404 => "00000000",
	405 => "00000000",
	406 => "00000000",
	407 => "00000000",
	408 => "00000000",
	409 => "00000000",
	410 => "00000000",
	411 => "00000000",
	412 => "00000000",
	413 => "00000000",
	414 => "00000000",
	415 => "00000000",
	416 => "00000000",
	417 => "00000000",
	418 => "00000000",
	419 => "00000000",
	420 => "00000000",
	421 => "00000000",
	422 => "00000000",
	423 => "00000000",
	424 => "00000000",
	425 => "00000000",
	426 => "00000000",
	427 => "00000000",
	428 => "00000000",
	429 => "00000000",
	430 => "00000000",
	431 => "00000000",
	432 => "00000000",
	433 => "00000000",
	434 => "00000000",
	435 => "00000000",
	436 => "00000000",
	437 => "00000000",
	438 => "00000000",
	439 => "00000000",
	440 => "00000000",
	441 => "00000000",
	442 => "00000000",
	443 => "00000000",
	448 => "00000000",
	449 => "00000000",
	450 => "00000000",
	451 => "00000000",
	452 => "00000000",
	453 => "00000000",
	454 => "00000000",
	455 => "00000000",
	456 => "00000000",
	457 => "00000000",
	458 => "00000000",
	459 => "00000000",
	460 => "00000000",
	461 => "00000000",
	462 => "00000000",
	463 => "00000000",
	464 => "00000000",
	465 => "00000000",
	466 => "00000000",
	467 => "00000000",
	468 => "00000000",
	469 => "00000000",
	470 => "00000000",
	471 => "00000000",
	472 => "00000000",
	473 => "00000000",
	474 => "00000000",
	475 => "00000000",
	476 => "00000000",
	477 => "00000000",
	478 => "00000000",
	479 => "00000000",
	480 => "00000000",
	481 => "00000000",
	482 => "00000000",
	483 => "00000000",
	484 => "00000000",
	485 => "00000000",
	486 => "00000000",
	487 => "00000000",
	488 => "00000000",
	489 => "00000000",
	490 => "00000000",
	491 => "00000000",
	492 => "00000000",
	493 => "00000000",
	494 => "00000000",
	495 => "00000000",
	496 => "00000000",
	497 => "00000000",
	498 => "00000000",
	499 => "00000000",
	500 => "00000000",
	501 => "00000000",
	502 => "00000000",
	503 => "00000000",
	504 => "00000000",
	505 => "00000000",
	506 => "00000000",
	507 => "00000000",
	512 => "00000000",
	513 => "00000000",
	514 => "00000000",
	515 => "00000000",
	516 => "00000000",
	517 => "00000000",
	518 => "00000000",
	519 => "00000000",
	520 => "00000000",
	521 => "00000000",
	522 => "00000000",
	523 => "00000000",
	524 => "00000000",
	525 => "00000000",
	526 => "00000000",
	527 => "00000000",
	528 => "00000000",
	529 => "00000000",
	530 => "00000000",
	531 => "00000000",
	532 => "00000000",
	533 => "00000000",
	534 => "00000000",
	535 => "00000000",
	536 => "00000000",
	537 => "00000000",
	538 => "00000000",
	539 => "00000000",
	540 => "00000000",
	541 => "00000000",
	542 => "00000000",
	543 => "00000000",
	544 => "00000000",
	545 => "00000000",
	546 => "00000000",
	547 => "00000000",
	548 => "00000000",
	549 => "00000000",
	550 => "00000000",
	551 => "00000000",
	552 => "00000000",
	553 => "00000000",
	554 => "00000000",
	555 => "00000000",
	556 => "00000000",
	557 => "00000000",
	558 => "00000000",
	559 => "00000000",
	560 => "00000000",
	561 => "00000000",
	562 => "00000000",
	563 => "00000000",
	564 => "00000000",
	565 => "00000000",
	566 => "00000000",
	567 => "00000000",
	568 => "00000000",
	569 => "00000000",
	570 => "00000000",
	571 => "00000000",
	576 => "00000000",
	577 => "00000000",
	578 => "00000000",
	579 => "00000000",
	580 => "00000000",
	581 => "00000000",
	582 => "00000000",
	583 => "00000000",
	584 => "00000000",
	585 => "00000000",
	586 => "00000000",
	587 => "00000000",
	588 => "00000000",
	589 => "00000000",
	590 => "00000000",
	591 => "00000000",
	592 => "00000000",
	593 => "00000000",
	594 => "00000000",
	595 => "00000000",
	596 => "00000000",
	597 => "00000000",
	598 => "00000000",
	599 => "00000000",
	600 => "00000000",
	601 => "00000000",
	602 => "00000000",
	603 => "00000000",
	604 => "00000000",
	605 => "00000000",
	606 => "00000000",
	607 => "00000000",
	608 => "00000000",
	609 => "00000000",
	610 => "00000000",
	611 => "00000000",
	612 => "00000000",
	613 => "00000000",
	614 => "00000000",
	615 => "00000000",
	616 => "00000000",
	617 => "00000000",
	618 => "00000000",
	619 => "00000000",
	620 => "00000000",
	621 => "00000000",
	622 => "00000000",
	623 => "00000000",
	624 => "00000000",
	625 => "00000000",
	626 => "00000000",
	627 => "00000000",
	628 => "00000000",
	629 => "00000000",
	630 => "00000000",
	631 => "00000000",
	632 => "00000000",
	633 => "00000000",
	634 => "00000000",
	635 => "00000000",
	640 => "00000000",
	641 => "00000000",
	642 => "00000000",
	643 => "00000000",
	644 => "00000000",
	645 => "00000000",
	646 => "00000000",
	647 => "00000000",
	648 => "00000000",
	649 => "00000000",
	650 => "00000000",
	651 => "00000000",
	652 => "00000000",
	653 => "00000000",
	654 => "00000000",
	655 => "00000000",
	656 => "00000000",
	657 => "00000000",
	658 => "00000000",
	659 => "00000000",
	660 => "00000000",
	661 => "00000000",
	662 => "00000000",
	663 => "00000000",
	664 => "00000000",
	665 => "00000000",
	666 => "00000000",
	667 => "00000000",
	668 => "00000000",
	669 => "00000000",
	670 => "00000000",
	671 => "00000000",
	672 => "00000000",
	673 => "00000000",
	674 => "00000000",
	675 => "00000000",
	676 => "00000000",
	677 => "00000000",
	678 => "00000000",
	679 => "00000000",
	680 => "00000000",
	681 => "00000000",
	682 => "00000000",
	683 => "00000000",
	684 => "00000000",
	685 => "00000000",
	686 => "00000000",
	687 => "00000000",
	688 => "00000000",
	689 => "00000000",
	690 => "00000000",
	691 => "00000000",
	692 => "00000000",
	693 => "00000000",
	694 => "00000000",
	695 => "00000000",
	696 => "00000000",
	697 => "00000000",
	698 => "00000000",
	699 => "00000000",
	704 => "00000000",
	705 => "00000000",
	706 => "00000000",
	707 => "00000000",
	708 => "00000000",
	709 => "00000000",
	710 => "00000000",
	711 => "00000000",
	712 => "00000000",
	713 => "00000000",
	714 => "00000000",
	715 => "00000000",
	716 => "00000000",
	717 => "00000000",
	718 => "00000000",
	719 => "00000000",
	720 => "00000000",
	721 => "00000000",
	722 => "00000000",
	723 => "00000000",
	724 => "00000000",
	725 => "00000000",
	726 => "00000000",
	727 => "00000000",
	728 => "00000000",
	729 => "00000000",
	730 => "00000000",
	731 => "00000000",
	732 => "00000000",
	733 => "00000000",
	734 => "00000000",
	735 => "00000000",
	736 => "00000000",
	737 => "00000000",
	738 => "00000000",
	739 => "00000000",
	740 => "00000000",
	741 => "00000000",
	742 => "00000000",
	743 => "00000000",
	744 => "00000000",
	745 => "00000000",
	746 => "00000000",
	747 => "00000000",
	748 => "00000000",
	749 => "00000000",
	750 => "00000000",
	751 => "00000000",
	752 => "00000000",
	753 => "00000000",
	754 => "00000000",
	755 => "00000000",
	756 => "00000000",
	757 => "00000000",
	758 => "00000000",
	759 => "00000000",
	760 => "00000000",
	761 => "00000000",
	762 => "00000000",
	763 => "00000000",
	768 => "00000000",
	769 => "00000000",
	770 => "00000000",
	771 => "00000000",
	772 => "00000000",
	773 => "00000000",
	774 => "00000000",
	775 => "00000000",
	776 => "00000000",
	777 => "00000000",
	778 => "00000000",
	779 => "00000000",
	780 => "00000000",
	781 => "00000000",
	782 => "00000000",
	783 => "00000000",
	784 => "00000000",
	785 => "00000000",
	786 => "00000000",
	787 => "00000000",
	788 => "00000000",
	789 => "00000000",
	790 => "00000000",
	791 => "00000000",
	792 => "00000000",
	793 => "00000000",
	794 => "00000000",
	795 => "00000000",
	796 => "00000000",
	797 => "00000000",
	798 => "00000000",
	799 => "00000000",
	800 => "00000000",
	801 => "00000000",
	802 => "00000000",
	803 => "00000000",
	804 => "00000000",
	805 => "00000000",
	806 => "00000000",
	807 => "00000000",
	808 => "00000000",
	809 => "00000000",
	810 => "00000000",
	811 => "00000000",
	812 => "00000000",
	813 => "00000000",
	814 => "00000000",
	815 => "00000000",
	816 => "00000000",
	817 => "00000000",
	818 => "00000000",
	819 => "00000000",
	820 => "00000000",
	821 => "00000000",
	822 => "00000000",
	823 => "00000000",
	824 => "00000000",
	825 => "00000000",
	826 => "00000000",
	827 => "00000000",
	832 => "00000000",
	833 => "00000000",
	834 => "00000000",
	835 => "00000000",
	836 => "00000000",
	837 => "00000000",
	838 => "00000000",
	839 => "00000000",
	840 => "00000000",
	841 => "00000000",
	842 => "00000000",
	843 => "00000000",
	844 => "00000000",
	845 => "00000000",
	846 => "00000000",
	847 => "00000000",
	848 => "00000000",
	849 => "00000000",
	850 => "00000000",
	851 => "00000000",
	852 => "00000000",
	853 => "00000000",
	854 => "00000000",
	855 => "00000000",
	856 => "00000000",
	857 => "00000000",
	858 => "00000000",
	859 => "00000000",
	860 => "00000000",
	861 => "00000000",
	862 => "00000000",
	863 => "00000000",
	864 => "00000000",
	865 => "00000000",
	866 => "00000000",
	867 => "00000000",
	868 => "00000000",
	869 => "00000000",
	870 => "00000000",
	871 => "00000000",
	872 => "00000000",
	873 => "00000000",
	874 => "00000000",
	875 => "00000000",
	876 => "00000000",
	877 => "00000000",
	878 => "00000000",
	879 => "00000000",
	880 => "00000000",
	881 => "00000000",
	882 => "00000000",
	883 => "00000000",
	884 => "00000000",
	885 => "00000000",
	886 => "00000000",
	887 => "00000000",
	888 => "00000000",
	889 => "00000000",
	890 => "00000000",
	891 => "00000000",
	896 => "00000000",
	897 => "00000000",
	898 => "00000000",
	899 => "00000000",
	900 => "00000000",
	901 => "00000000",
	902 => "00000000",
	903 => "00000000",
	904 => "00000000",
	905 => "00000000",
	906 => "00000000",
	907 => "00000000",
	908 => "00000000",
	909 => "00000000",
	910 => "00000000",
	911 => "00000000",
	912 => "00000000",
	913 => "00000000",
	914 => "00000000",
	915 => "00000000",
	916 => "00000000",
	917 => "00000000",
	918 => "00000000",
	919 => "00000000",
	920 => "00000000",
	921 => "00000000",
	922 => "00000000",
	923 => "00000000",
	924 => "00000000",
	925 => "00000000",
	926 => "00000000",
	927 => "00000000",
	928 => "00000000",
	929 => "00000000",
	930 => "00000000",
	931 => "00000000",
	932 => "00000000",
	933 => "00000000",
	934 => "00000000",
	935 => "00000000",
	936 => "00000000",
	937 => "00000000",
	938 => "00000000",
	939 => "00000000",
	940 => "00000000",
	941 => "00000000",
	942 => "00000000",
	943 => "00000000",
	944 => "00000000",
	945 => "00000000",
	946 => "00000000",
	947 => "00000000",
	948 => "00000000",
	949 => "00000000",
	950 => "00000000",
	951 => "00000000",
	952 => "00000000",
	953 => "00000000",
	954 => "00000000",
	955 => "00000000",
	960 => "00000000",
	961 => "00000000",
	962 => "00000000",
	963 => "00000000",
	964 => "00000000",
	965 => "00000000",
	966 => "00000000",
	967 => "00000000",
	968 => "00000000",
	969 => "00000000",
	970 => "00000000",
	971 => "00000000",
	972 => "00000000",
	973 => "00000000",
	974 => "00000000",
	975 => "00000000",
	976 => "00000000",
	977 => "00000000",
	978 => "00000000",
	979 => "00000000",
	980 => "00000000",
	981 => "00000000",
	982 => "00000000",
	983 => "00000000",
	984 => "00000000",
	985 => "00000000",
	986 => "00000000",
	987 => "00000000",
	988 => "00000000",
	989 => "00000000",
	990 => "00000000",
	991 => "00000000",
	992 => "00000000",
	993 => "00000000",
	994 => "00000000",
	995 => "00000000",
	996 => "00000000",
	997 => "00000000",
	998 => "00000000",
	999 => "00000000",
	1000 => "00000000",
	1001 => "00000000",
	1002 => "00000000",
	1003 => "00000000",
	1004 => "00000000",
	1005 => "00000000",
	1006 => "00000000",
	1007 => "00000000",
	1008 => "00000000",
	1009 => "00000000",
	1010 => "00000000",
	1011 => "00000000",
	1012 => "00000000",
	1013 => "00000000",
	1014 => "00000000",
	1015 => "00000000",
	1016 => "00000000",
	1017 => "00000000",
	1018 => "00000000",
	1019 => "00000000",
	1024 => "00000000",
	1025 => "00000000",
	1026 => "00000000",
	1027 => "00000000",
	1028 => "00000000",
	1029 => "00000000",
	1030 => "00000000",
	1031 => "00000000",
	1032 => "00000000",
	1033 => "00000000",
	1034 => "00000000",
	1035 => "00000000",
	1036 => "00000000",
	1037 => "00000000",
	1038 => "00000000",
	1039 => "00000000",
	1040 => "00000000",
	1041 => "00000000",
	1042 => "00000000",
	1043 => "00000000",
	1044 => "00000000",
	1045 => "00000000",
	1046 => "00000000",
	1047 => "00000000",
	1048 => "00000000",
	1049 => "00000000",
	1050 => "00000000",
	1051 => "00000000",
	1052 => "00000000",
	1053 => "00000000",
	1054 => "00000000",
	1055 => "00000000",
	1056 => "00000000",
	1057 => "00000000",
	1058 => "00000000",
	1059 => "00000000",
	1060 => "00000000",
	1061 => "00000000",
	1062 => "00000000",
	1063 => "00000000",
	1064 => "00000000",
	1065 => "00000000",
	1066 => "00000000",
	1067 => "00000000",
	1068 => "00000000",
	1069 => "00000000",
	1070 => "00000000",
	1071 => "00000000",
	1072 => "00000000",
	1073 => "00000000",
	1074 => "00000000",
	1075 => "00000000",
	1076 => "00000000",
	1077 => "00000000",
	1078 => "00000000",
	1079 => "00000000",
	1080 => "00000000",
	1081 => "00000000",
	1082 => "00000000",
	1083 => "00000000",
	1088 => "00000000",
	1089 => "00000000",
	1090 => "00000000",
	1091 => "00000000",
	1092 => "00000000",
	1093 => "00000000",
	1094 => "00000000",
	1095 => "00000000",
	1096 => "00000000",
	1097 => "00000000",
	1098 => "00000000",
	1099 => "00000000",
	1100 => "00000000",
	1101 => "00000000",
	1102 => "00000000",
	1103 => "00000000",
	1104 => "00000000",
	1105 => "00000000",
	1106 => "00000000",
	1107 => "00000000",
	1108 => "00000000",
	1109 => "00000000",
	1110 => "00000000",
	1111 => "00000000",
	1112 => "00000000",
	1113 => "00000000",
	1114 => "00000000",
	1115 => "00000000",
	1116 => "00000000",
	1117 => "00000000",
	1118 => "00000000",
	1119 => "00000000",
	1120 => "00000000",
	1121 => "00000000",
	1122 => "00000000",
	1123 => "00000000",
	1124 => "00000000",
	1125 => "00000000",
	1126 => "00000000",
	1127 => "00000000",
	1128 => "00000000",
	1129 => "00000000",
	1130 => "00000000",
	1131 => "00000000",
	1132 => "00000000",
	1133 => "00000000",
	1134 => "00000000",
	1135 => "00000000",
	1136 => "00000000",
	1137 => "00000000",
	1138 => "00000000",
	1139 => "00000000",
	1140 => "00000000",
	1141 => "00000000",
	1142 => "00000000",
	1143 => "00000000",
	1144 => "00000000",
	1145 => "00000000",
	1146 => "00000000",
	1147 => "00000000",
	1152 => "00000000",
	1153 => "00000000",
	1154 => "00000000",
	1155 => "00000000",
	1156 => "00000000",
	1157 => "00000000",
	1158 => "00000000",
	1159 => "00000000",
	1160 => "00000000",
	1161 => "00000000",
	1162 => "00000000",
	1163 => "00000000",
	1164 => "00000000",
	1165 => "00000000",
	1166 => "00000000",
	1167 => "00000000",
	1168 => "00000000",
	1169 => "00000000",
	1170 => "00000000",
	1171 => "00000000",
	1172 => "00000000",
	1173 => "00000000",
	1174 => "00000000",
	1175 => "00000000",
	1176 => "00000000",
	1177 => "00000000",
	1178 => "00000000",
	1179 => "00000000",
	1180 => "00000000",
	1181 => "00000000",
	1182 => "00000000",
	1183 => "00000000",
	1184 => "00000000",
	1185 => "00000000",
	1186 => "00000000",
	1187 => "00000000",
	1188 => "00000000",
	1189 => "00000000",
	1190 => "00000000",
	1191 => "00000000",
	1192 => "00000000",
	1193 => "00000000",
	1194 => "00000000",
	1195 => "00000000",
	1196 => "00000000",
	1197 => "00000000",
	1198 => "00000000",
	1199 => "00000000",
	1200 => "00000000",
	1201 => "00000000",
	1202 => "00000000",
	1203 => "00000000",
	1204 => "00000000",
	1205 => "00000000",
	1206 => "00000000",
	1207 => "00000000",
	1208 => "00000000",
	1209 => "00000000",
	1210 => "00000000",
	1211 => "00000000",
	1216 => "00000000",
	1217 => "00000000",
	1218 => "00000000",
	1219 => "00000000",
	1220 => "00000000",
	1221 => "00000000",
	1222 => "00000000",
	1223 => "00000000",
	1224 => "00000000",
	1225 => "00000000",
	1226 => "00000000",
	1227 => "00000000",
	1228 => "00000000",
	1229 => "00000000",
	1230 => "00000000",
	1231 => "00000000",
	1232 => "00000000",
	1233 => "00000000",
	1234 => "00000000",
	1235 => "00000000",
	1236 => "00000000",
	1237 => "00000000",
	1238 => "00000000",
	1239 => "00000000",
	1240 => "00000000",
	1241 => "00000000",
	1242 => "00000000",
	1243 => "00000000",
	1244 => "00000000",
	1245 => "00000000",
	1246 => "00000000",
	1247 => "00000000",
	1248 => "00000000",
	1249 => "00000000",
	1250 => "00000000",
	1251 => "00000000",
	1252 => "00000000",
	1253 => "00000000",
	1254 => "00000000",
	1255 => "00000000",
	1256 => "00000000",
	1257 => "00000000",
	1258 => "00000000",
	1259 => "00000000",
	1260 => "00000000",
	1261 => "00000000",
	1262 => "00000000",
	1263 => "00000000",
	1264 => "00000000",
	1265 => "00000000",
	1266 => "00000000",
	1267 => "00000000",
	1268 => "00000000",
	1269 => "00000000",
	1270 => "00000000",
	1271 => "00000000",
	1272 => "00000000",
	1273 => "00000000",
	1274 => "00000000",
	1275 => "00000000",
	1280 => "00000000",
	1281 => "00000000",
	1282 => "00000000",
	1283 => "00000000",
	1284 => "00000000",
	1285 => "00000000",
	1286 => "00000000",
	1287 => "00000000",
	1288 => "00000000",
	1289 => "00000000",
	1290 => "00000000",
	1291 => "00000000",
	1292 => "00000000",
	1293 => "00000000",
	1294 => "00000000",
	1295 => "00000000",
	1296 => "00000000",
	1297 => "00000000",
	1298 => "00000000",
	1299 => "00000000",
	1300 => "00000000",
	1301 => "00000000",
	1302 => "00000000",
	1303 => "00000000",
	1304 => "00000000",
	1305 => "00000000",
	1306 => "00000000",
	1307 => "00000000",
	1308 => "00000000",
	1309 => "00000000",
	1310 => "00000000",
	1311 => "00000000",
	1312 => "00000000",
	1313 => "00000000",
	1314 => "00000000",
	1315 => "00000000",
	1316 => "00000000",
	1317 => "00000000",
	1318 => "00000000",
	1319 => "00000000",
	1320 => "00000000",
	1321 => "00000000",
	1322 => "00000000",
	1323 => "00000000",
	1324 => "00000000",
	1325 => "00000000",
	1326 => "00000000",
	1327 => "00000000",
	1328 => "00000000",
	1329 => "00000000",
	1330 => "00000000",
	1331 => "00000000",
	1332 => "00000000",
	1333 => "00000000",
	1334 => "00000000",
	1335 => "00000000",
	1336 => "00000000",
	1337 => "00000000",
	1338 => "00000000",
	1339 => "00000000",
	1344 => "00000000",
	1345 => "00000000",
	1346 => "00000000",
	1347 => "00000000",
	1348 => "00000000",
	1349 => "00000000",
	1350 => "00000000",
	1351 => "00000000",
	1352 => "00000000",
	1353 => "00000000",
	1354 => "00000000",
	1355 => "00000000",
	1356 => "00000000",
	1357 => "00000000",
	1358 => "00000000",
	1359 => "00000000",
	1360 => "00000000",
	1361 => "00000000",
	1362 => "00000000",
	1363 => "00000000",
	1364 => "00000000",
	1365 => "00000000",
	1366 => "00000000",
	1367 => "00000000",
	1368 => "00000000",
	1369 => "00000000",
	1370 => "00000000",
	1371 => "00000000",
	1372 => "00000000",
	1373 => "00000000",
	1374 => "00000000",
	1375 => "00000000",
	1376 => "00000000",
	1377 => "00000000",
	1378 => "00000000",
	1379 => "00000000",
	1380 => "00000000",
	1381 => "00000000",
	1382 => "00000000",
	1383 => "00000000",
	1384 => "00000000",
	1385 => "00000000",
	1386 => "00000000",
	1387 => "00000000",
	1388 => "00000000",
	1389 => "00000000",
	1390 => "00000000",
	1391 => "00000000",
	1392 => "00000000",
	1393 => "00000000",
	1394 => "00000000",
	1395 => "00000000",
	1396 => "00000000",
	1397 => "00000000",
	1398 => "00000000",
	1399 => "00000000",
	1400 => "00000000",
	1401 => "00000000",
	1402 => "00000000",
	1403 => "00000000",
	1408 => "00000000",
	1409 => "00000000",
	1410 => "00000000",
	1411 => "00000000",
	1412 => "00000000",
	1413 => "00000000",
	1414 => "00000000",
	1415 => "00000000",
	1416 => "00000000",
	1417 => "00000000",
	1418 => "00000000",
	1419 => "00000000",
	1420 => "00000000",
	1421 => "00000000",
	1422 => "00000000",
	1423 => "00000000",
	1424 => "00000000",
	1425 => "00000000",
	1426 => "00000000",
	1427 => "00000000",
	1428 => "00000000",
	1429 => "00000000",
	1430 => "00000000",
	1431 => "00000000",
	1432 => "00000000",
	1433 => "00000000",
	1434 => "00000000",
	1435 => "00000000",
	1436 => "00000000",
	1437 => "00000000",
	1438 => "00000000",
	1439 => "00000000",
	1440 => "00000000",
	1441 => "00000000",
	1442 => "00000000",
	1443 => "00000000",
	1444 => "00000000",
	1445 => "00000000",
	1446 => "00000000",
	1447 => "00000000",
	1448 => "00000000",
	1449 => "00000000",
	1450 => "00000000",
	1451 => "00000000",
	1452 => "00000000",
	1453 => "00000000",
	1454 => "00000000",
	1455 => "00000000",
	1456 => "00000000",
	1457 => "00000000",
	1458 => "00000000",
	1459 => "00000000",
	1460 => "00000000",
	1461 => "00000000",
	1462 => "00000000",
	1463 => "00000000",
	1464 => "00000000",
	1465 => "00000000",
	1466 => "00000000",
	1467 => "00000000",
	1472 => "00000000",
	1473 => "00000000",
	1474 => "00000000",
	1475 => "00000000",
	1476 => "00000000",
	1477 => "00000000",
	1478 => "00000000",
	1479 => "00000000",
	1480 => "00000000",
	1481 => "00000000",
	1482 => "00000000",
	1483 => "00000000",
	1484 => "00000000",
	1485 => "00000000",
	1486 => "00000000",
	1487 => "00000000",
	1488 => "00000000",
	1489 => "00000000",
	1490 => "00000000",
	1491 => "00000000",
	1492 => "00000000",
	1493 => "00000000",
	1494 => "00000000",
	1495 => "00000000",
	1496 => "00000000",
	1497 => "00000000",
	1498 => "00000000",
	1499 => "00000000",
	1500 => "00000000",
	1501 => "00000000",
	1502 => "00000000",
	1503 => "00000000",
	1504 => "00000000",
	1505 => "00000000",
	1506 => "00000000",
	1507 => "00000000",
	1508 => "00000000",
	1509 => "00000000",
	1510 => "00000000",
	1511 => "00000000",
	1512 => "00000000",
	1513 => "00000000",
	1514 => "00000000",
	1515 => "00000000",
	1516 => "00000000",
	1517 => "00000000",
	1518 => "00000000",
	1519 => "00000000",
	1520 => "00000000",
	1521 => "00000000",
	1522 => "00000000",
	1523 => "00000000",
	1524 => "00000000",
	1525 => "00000000",
	1526 => "00000000",
	1527 => "00000000",
	1528 => "00000000",
	1529 => "00000000",
	1530 => "00000000",
	1531 => "00000000",
	1536 => "00000000",
	1537 => "00000000",
	1538 => "00000000",
	1539 => "00000000",
	1540 => "00000000",
	1541 => "00000000",
	1542 => "00000000",
	1543 => "00000000",
	1544 => "00000000",
	1545 => "00000000",
	1546 => "00000000",
	1547 => "00000000",
	1548 => "00000000",
	1549 => "00000000",
	1550 => "00000000",
	1551 => "00000000",
	1552 => "00000000",
	1553 => "00000000",
	1554 => "00000000",
	1555 => "00000000",
	1556 => "00000000",
	1557 => "00000000",
	1558 => "00000000",
	1559 => "00000000",
	1560 => "00000000",
	1561 => "00000000",
	1562 => "00000000",
	1563 => "00000000",
	1564 => "00000000",
	1565 => "00000000",
	1566 => "00000000",
	1567 => "00000000",
	1568 => "00000000",
	1569 => "00000000",
	1570 => "00000000",
	1571 => "00000000",
	1572 => "00000000",
	1573 => "00000000",
	1574 => "00000000",
	1575 => "00000000",
	1576 => "00000000",
	1577 => "00000000",
	1578 => "00000000",
	1579 => "00000000",
	1580 => "00000000",
	1581 => "00000000",
	1582 => "00000000",
	1583 => "00000000",
	1584 => "00000000",
	1585 => "00000000",
	1586 => "00000000",
	1587 => "00000000",
	1588 => "00000000",
	1589 => "00000000",
	1590 => "00000000",
	1591 => "00000000",
	1592 => "00000000",
	1593 => "00000000",
	1594 => "00000000",
	1595 => "00000000",
	1600 => "00000000",
	1601 => "00000000",
	1602 => "00000000",
	1603 => "00000000",
	1604 => "00000000",
	1605 => "00000000",
	1606 => "00000000",
	1607 => "00000000",
	1608 => "00000000",
	1609 => "00000000",
	1610 => "00000000",
	1611 => "00000000",
	1612 => "00000000",
	1613 => "00000000",
	1614 => "00000000",
	1615 => "00000000",
	1616 => "00000000",
	1617 => "00000000",
	1618 => "00000000",
	1619 => "00000000",
	1620 => "00000000",
	1621 => "00000000",
	1622 => "00000000",
	1623 => "00000000",
	1624 => "00000000",
	1625 => "00000000",
	1626 => "00000000",
	1627 => "00000000",
	1628 => "00000000",
	1629 => "00000000",
	1630 => "00000000",
	1631 => "00000000",
	1632 => "00000000",
	1633 => "00000000",
	1634 => "00000000",
	1635 => "00000000",
	1636 => "00000000",
	1637 => "00000000",
	1638 => "00000000",
	1639 => "00000000",
	1640 => "00000000",
	1641 => "00000000",
	1642 => "00000000",
	1643 => "00000000",
	1644 => "00000000",
	1645 => "00000000",
	1646 => "00000000",
	1647 => "00000000",
	1648 => "00000000",
	1649 => "00000000",
	1650 => "00000000",
	1651 => "00000000",
	1652 => "00000000",
	1653 => "00000000",
	1654 => "00000000",
	1655 => "00000000",
	1656 => "00000000",
	1657 => "00000000",
	1658 => "00000000",
	1659 => "00000000",
	1664 => "00000000",
	1665 => "00000000",
	1666 => "00000000",
	1667 => "00000000",
	1668 => "00000000",
	1669 => "00000000",
	1670 => "00000000",
	1671 => "00000000",
	1672 => "00000000",
	1673 => "00000000",
	1674 => "00000000",
	1675 => "00000000",
	1676 => "00000000",
	1677 => "00000000",
	1678 => "00000000",
	1679 => "00000000",
	1680 => "00000000",
	1681 => "00000000",
	1682 => "00000000",
	1683 => "00000000",
	1684 => "00000000",
	1685 => "00000000",
	1686 => "00000000",
	1687 => "00000000",
	1688 => "00000000",
	1689 => "00000000",
	1690 => "00000000",
	1691 => "00000000",
	1692 => "00000000",
	1693 => "00000000",
	1694 => "00000000",
	1695 => "00000000",
	1696 => "00000000",
	1697 => "00000000",
	1698 => "00000000",
	1699 => "00000000",
	1700 => "00000000",
	1701 => "00000000",
	1702 => "00000000",
	1703 => "00000000",
	1704 => "00000000",
	1705 => "00000000",
	1706 => "00000000",
	1707 => "00000000",
	1708 => "00000000",
	1709 => "00000000",
	1710 => "00000000",
	1711 => "00000000",
	1712 => "00000000",
	1713 => "00000000",
	1714 => "00000000",
	1715 => "00000000",
	1716 => "00000000",
	1717 => "00000000",
	1718 => "00000000",
	1719 => "00000000",
	1720 => "00000000",
	1721 => "00000000",
	1722 => "00000000",
	1723 => "00000000",
	1728 => "00000000",
	1729 => "00000000",
	1730 => "00000000",
	1731 => "00000000",
	1732 => "00000000",
	1733 => "00000000",
	1734 => "00000000",
	1735 => "00000000",
	1736 => "00000000",
	1737 => "00000000",
	1738 => "00000000",
	1739 => "00000000",
	1740 => "00000000",
	1741 => "00000000",
	1742 => "00000000",
	1743 => "00000000",
	1744 => "00000000",
	1745 => "00000000",
	1746 => "00000000",
	1747 => "00000000",
	1748 => "00000000",
	1749 => "00000000",
	1750 => "00000000",
	1751 => "00000000",
	1752 => "00000000",
	1753 => "00000000",
	1754 => "00000000",
	1755 => "00000000",
	1756 => "00000000",
	1757 => "00000000",
	1758 => "00000000",
	1759 => "00000000",
	1760 => "00000000",
	1761 => "00000000",
	1762 => "00000000",
	1763 => "00000000",
	1764 => "00000000",
	1765 => "00000000",
	1766 => "00000000",
	1767 => "00000000",
	1768 => "00000000",
	1769 => "00000000",
	1770 => "00000000",
	1771 => "00000000",
	1772 => "00000000",
	1773 => "00000000",
	1774 => "00000000",
	1775 => "00000000",
	1776 => "00000000",
	1777 => "00000000",
	1778 => "00000000",
	1779 => "00000000",
	1780 => "00000000",
	1781 => "00000000",
	1782 => "00000000",
	1783 => "00000000",
	1784 => "00000000",
	1785 => "00000000",
	1786 => "00000000",
	1787 => "00000000",
	1792 => "00000000",
	1793 => "00000000",
	1794 => "00000000",
	1795 => "00000000",
	1796 => "00000000",
	1797 => "00000000",
	1798 => "00000000",
	1799 => "00000000",
	1800 => "00000000",
	1801 => "00000000",
	1802 => "00000000",
	1803 => "00000000",
	1804 => "00000000",
	1805 => "00000000",
	1806 => "00000000",
	1807 => "00000000",
	1808 => "00000000",
	1809 => "00000000",
	1810 => "00000000",
	1811 => "00000000",
	1812 => "00000000",
	1813 => "00000000",
	1814 => "00000000",
	1815 => "00000000",
	1816 => "00000000",
	1817 => "00000000",
	1818 => "00000000",
	1819 => "00000000",
	1820 => "00000000",
	1821 => "00000000",
	1822 => "00000000",
	1823 => "00000000",
	1824 => "00000000",
	1825 => "00000000",
	1826 => "00000000",
	1827 => "00000000",
	1828 => "00000000",
	1829 => "00000000",
	1830 => "00000000",
	1831 => "00000000",
	1832 => "00000000",
	1833 => "00000000",
	1834 => "00000000",
	1835 => "00000000",
	1836 => "00000000",
	1837 => "00000000",
	1838 => "00000000",
	1839 => "00000000",
	1840 => "00000000",
	1841 => "00000000",
	1842 => "00000000",
	1843 => "00000000",
	1844 => "00000000",
	1845 => "00000000",
	1846 => "00000000",
	1847 => "00000000",
	1848 => "00000000",
	1849 => "00000000",
	1850 => "00000000",
	1851 => "00000000",
	1856 => "00000000",
	1857 => "00000000",
	1858 => "00000000",
	1859 => "00000000",
	1860 => "00000000",
	1861 => "00000000",
	1862 => "00000000",
	1863 => "00000000",
	1864 => "00000000",
	1865 => "00000000",
	1866 => "00000000",
	1867 => "00000000",
	1868 => "00000000",
	1869 => "00000000",
	1870 => "00000000",
	1871 => "00000000",
	1872 => "00000000",
	1873 => "00000000",
	1874 => "00000000",
	1875 => "00000000",
	1876 => "00000000",
	1877 => "00000000",
	1878 => "00000000",
	1879 => "00000000",
	1880 => "00000000",
	1881 => "00000000",
	1882 => "00000000",
	1883 => "00000000",
	1884 => "00000000",
	1885 => "00000000",
	1886 => "00000000",
	1887 => "00000000",
	1888 => "00000000",
	1889 => "00000000",
	1890 => "00000000",
	1891 => "00000000",
	1892 => "00000000",
	1893 => "00000000",
	1894 => "00000000",
	1895 => "00000000",
	1896 => "00000000",
	1897 => "00000000",
	1898 => "00000000",
	1899 => "00000000",
	1900 => "00000000",
	1901 => "00000000",
	1902 => "00000000",
	1903 => "00000000",
	1904 => "00000000",
	1905 => "00000000",
	1906 => "00000000",
	1907 => "00000000",
	1908 => "00000000",
	1909 => "00000000",
	1910 => "00000000",
	1911 => "00000000",
	1912 => "00000000",
	1913 => "00000000",
	1914 => "00000000",
	1915 => "00000000",
	1920 => "00000000",
	1921 => "00000000",
	1922 => "00000000",
	1923 => "00000000",
	1924 => "00000000",
	1925 => "00000000",
	1926 => "00000000",
	1927 => "00000000",
	1928 => "00000000",
	1929 => "00000000",
	1930 => "00000000",
	1931 => "00000000",
	1932 => "00000000",
	1933 => "00000000",
	1934 => "00000000",
	1935 => "00000000",
	1936 => "00000000",
	1937 => "00000000",
	1938 => "00000000",
	1939 => "00000000",
	1940 => "00000000",
	1941 => "00000000",
	1942 => "00000000",
	1943 => "00000000",
	1944 => "00000000",
	1945 => "00000000",
	1946 => "00000000",
	1947 => "00000000",
	1948 => "00000000",
	1949 => "00000000",
	1950 => "00000000",
	1951 => "00000000",
	1952 => "00000000",
	1953 => "00000000",
	1954 => "00000000",
	1955 => "00000000",
	1956 => "00000000",
	1957 => "00000000",
	1958 => "00000000",
	1959 => "00000000",
	1960 => "00000000",
	1961 => "00000000",
	1962 => "00000000",
	1963 => "00000000",
	1964 => "00000000",
	1965 => "00000000",
	1966 => "00000000",
	1967 => "00000000",
	1968 => "00000000",
	1969 => "00000000",
	1970 => "00000000",
	1971 => "00000000",
	1972 => "00000000",
	1973 => "00000000",
	1974 => "00000000",
	1975 => "00000000",
	1976 => "00000000",
	1977 => "00000000",
	1978 => "00000000",
	1979 => "00000000",
	1984 => "00000000",
	1985 => "00000000",
	1986 => "00000000",
	1987 => "00000000",
	1988 => "00000000",
	1989 => "00000000",
	1990 => "00000000",
	1991 => "00000000",
	1992 => "00000000",
	1993 => "00000000",
	1994 => "00000000",
	1995 => "00000000",
	1996 => "00000000",
	1997 => "00000000",
	1998 => "00000000",
	1999 => "00000000",
	2000 => "00000000",
	2001 => "00000000",
	2002 => "00000000",
	2003 => "00000000",
	2004 => "00000000",
	2005 => "00000000",
	2006 => "00000000",
	2007 => "00000000",
	2008 => "00000000",
	2009 => "00000000",
	2010 => "00000000",
	2011 => "00000000",
	2012 => "00000000",
	2013 => "00000000",
	2014 => "00000000",
	2015 => "00000000",
	2016 => "00000000",
	2017 => "00000000",
	2018 => "00000000",
	2019 => "00000000",
	2020 => "00000000",
	2021 => "00000000",
	2022 => "00000000",
	2023 => "00000000",
	2024 => "00000000",
	2025 => "00000000",
	2026 => "00000000",
	2027 => "00000000",
	2028 => "00000000",
	2029 => "00000000",
	2030 => "00000000",
	2031 => "00000000",
	2032 => "00000000",
	2033 => "00000000",
	2034 => "00000000",
	2035 => "00000000",
	2036 => "00000000",
	2037 => "00000000",
	2038 => "00000000",
	2039 => "00000000",
	2040 => "00000000",
	2041 => "00000000",
	2042 => "00000000",
	2043 => "00000000",
	2048 => "00000000",
	2049 => "00000000",
	2050 => "00000000",
	2051 => "00000000",
	2052 => "00000000",
	2053 => "00000000",
	2054 => "00000000",
	2055 => "00000000",
	2056 => "00000000",
	2057 => "00000000",
	2058 => "00000000",
	2059 => "00000000",
	2060 => "00000000",
	2061 => "00000000",
	2062 => "00000000",
	2063 => "00000000",
	2064 => "00000000",
	2065 => "00000000",
	2066 => "00000000",
	2067 => "00000000",
	2068 => "00000000",
	2069 => "00000000",
	2070 => "00000000",
	2071 => "00000000",
	2072 => "00000000",
	2073 => "00000000",
	2074 => "00000000",
	2075 => "00000000",
	2076 => "00000000",
	2077 => "00000000",
	2078 => "00000000",
	2079 => "00000000",
	2080 => "00000000",
	2081 => "00000000",
	2082 => "00000000",
	2083 => "00000000",
	2084 => "00000000",
	2085 => "00000000",
	2086 => "00000000",
	2087 => "00000000",
	2088 => "00000000",
	2089 => "00000000",
	2090 => "00000000",
	2091 => "00000000",
	2092 => "00000000",
	2093 => "00000000",
	2094 => "00000000",
	2095 => "00000000",
	2096 => "00000000",
	2097 => "00000000",
	2098 => "00000000",
	2099 => "00000000",
	2100 => "00000000",
	2101 => "00000000",
	2102 => "00000000",
	2103 => "00000000",
	2104 => "00000000",
	2105 => "00000000",
	2106 => "00000000",
	2107 => "00000000",
	2112 => "00000000",
	2113 => "00000000",
	2114 => "00000000",
	2115 => "00000000",
	2116 => "00000000",
	2117 => "00000000",
	2118 => "00000000",
	2119 => "00000000",
	2120 => "00000000",
	2121 => "00000000",
	2122 => "00000000",
	2123 => "00000000",
	2124 => "00000000",
	2125 => "00000000",
	2126 => "00000000",
	2127 => "00000000",
	2128 => "00000000",
	2129 => "00000000",
	2130 => "00000000",
	2131 => "00000000",
	2132 => "00000000",
	2133 => "00000000",
	2134 => "00000000",
	2135 => "00000000",
	2136 => "00000000",
	2137 => "00000000",
	2138 => "00000000",
	2139 => "00000000",
	2140 => "00000000",
	2141 => "00000000",
	2142 => "00000000",
	2143 => "00000000",
	2144 => "00000000",
	2145 => "00000000",
	2146 => "00000000",
	2147 => "00000000",
	2148 => "00000000",
	2149 => "00000000",
	2150 => "00000000",
	2151 => "00000000",
	2152 => "00000000",
	2153 => "00000000",
	2154 => "00000000",
	2155 => "00000000",
	2156 => "00000000",
	2157 => "00000000",
	2158 => "00000000",
	2159 => "00000000",
	2160 => "00000000",
	2161 => "00000000",
	2162 => "00000000",
	2163 => "00000000",
	2164 => "00000000",
	2165 => "00000000",
	2166 => "00000000",
	2167 => "00000000",
	2168 => "00000000",
	2169 => "00000000",
	2170 => "00000000",
	2171 => "00000000",
	2176 => "00000000",
	2177 => "00000000",
	2178 => "00000000",
	2179 => "00000000",
	2180 => "00000000",
	2181 => "00000000",
	2182 => "00000000",
	2183 => "00000000",
	2184 => "00000000",
	2185 => "00000000",
	2186 => "00000000",
	2187 => "00000000",
	2188 => "00000000",
	2189 => "00000000",
	2190 => "00000000",
	2191 => "00000000",
	2192 => "00000000",
	2193 => "00000000",
	2194 => "00000000",
	2195 => "00000000",
	2196 => "00000000",
	2197 => "00000000",
	2198 => "00000000",
	2199 => "00000000",
	2200 => "00000000",
	2201 => "00000000",
	2202 => "00000000",
	2203 => "00000000",
	2204 => "00000000",
	2205 => "00000000",
	2206 => "00000000",
	2207 => "00000000",
	2208 => "00000000",
	2209 => "00000000",
	2210 => "00000000",
	2211 => "00000000",
	2212 => "00000000",
	2213 => "00000000",
	2214 => "00000000",
	2215 => "00000000",
	2216 => "00000000",
	2217 => "00000000",
	2218 => "00000000",
	2219 => "00000000",
	2220 => "00000000",
	2221 => "00000000",
	2222 => "00000000",
	2223 => "00000000",
	2224 => "00000000",
	2225 => "00000000",
	2226 => "00000000",
	2227 => "00000000",
	2228 => "00000000",
	2229 => "00000000",
	2230 => "00000000",
	2231 => "00000000",
	2232 => "00000000",
	2233 => "00000000",
	2234 => "00000000",
	2235 => "00000000",
	2240 => "00000000",
	2241 => "00000000",
	2242 => "00000000",
	2243 => "00000000",
	2244 => "00000000",
	2245 => "00000000",
	2246 => "00000000",
	2247 => "00000000",
	2248 => "00000000",
	2249 => "00000000",
	2250 => "00000000",
	2251 => "00000000",
	2252 => "00000000",
	2253 => "00000000",
	2254 => "00000000",
	2255 => "00000000",
	2256 => "00000000",
	2257 => "00000000",
	2258 => "00000000",
	2259 => "00000000",
	2260 => "00000000",
	2261 => "00000000",
	2262 => "00000000",
	2263 => "00000000",
	2264 => "00000000",
	2265 => "00000000",
	2266 => "00000000",
	2267 => "00000000",
	2268 => "00000000",
	2269 => "00000000",
	2270 => "00000000",
	2271 => "00000000",
	2272 => "00000000",
	2273 => "00000000",
	2274 => "00000000",
	2275 => "00000000",
	2276 => "00000000",
	2277 => "00000000",
	2278 => "00000000",
	2279 => "00000000",
	2280 => "00000000",
	2281 => "00000000",
	2282 => "00000000",
	2283 => "00000000",
	2284 => "00000000",
	2285 => "00000000",
	2286 => "00000000",
	2287 => "00000000",
	2288 => "00000000",
	2289 => "00000000",
	2290 => "00000000",
	2291 => "00000000",
	2292 => "00000000",
	2293 => "00000000",
	2294 => "00000000",
	2295 => "00000000",
	2296 => "00000000",
	2297 => "00000000",
	2298 => "00000000",
	2299 => "00000000",
	2304 => "00000000",
	2305 => "00000000",
	2306 => "00000000",
	2307 => "00000000",
	2308 => "00000000",
	2309 => "00000000",
	2310 => "00000000",
	2311 => "00000000",
	2312 => "00000000",
	2313 => "00000000",
	2314 => "00000000",
	2315 => "00000000",
	2316 => "00000000",
	2317 => "00000000",
	2318 => "00000000",
	2319 => "00000000",
	2320 => "00000000",
	2321 => "00000000",
	2322 => "00000000",
	2323 => "00000000",
	2324 => "00000000",
	2325 => "00000000",
	2326 => "00000000",
	2327 => "00000000",
	2328 => "00000000",
	2329 => "00000000",
	2330 => "00000000",
	2331 => "00000000",
	2332 => "00000000",
	2333 => "00000000",
	2334 => "00000000",
	2335 => "00000000",
	2336 => "00000000",
	2337 => "00000000",
	2338 => "00000000",
	2339 => "00000000",
	2340 => "00000000",
	2341 => "00000000",
	2342 => "00000000",
	2343 => "00000000",
	2344 => "00000000",
	2345 => "00000000",
	2346 => "00000000",
	2347 => "00000000",
	2348 => "00000000",
	2349 => "00000000",
	2350 => "00000000",
	2351 => "00000000",
	2352 => "00000000",
	2353 => "00000000",
	2354 => "00000000",
	2355 => "00000000",
	2356 => "00000000",
	2357 => "00000000",
	2358 => "00000000",
	2359 => "00000000",
	2360 => "00000000",
	2361 => "00000000",
	2362 => "00000000",
	2363 => "00000000",
	2368 => "00000000",
	2369 => "00000000",
	2370 => "00000000",
	2371 => "00000000",
	2372 => "00000000",
	2373 => "00000000",
	2374 => "00000000",
	2375 => "00000000",
	2376 => "00000000",
	2377 => "00000000",
	2378 => "00000000",
	2379 => "00000000",
	2380 => "00000000",
	2381 => "00000000",
	2382 => "00000000",
	2383 => "00000000",
	2384 => "00000000",
	2385 => "00000000",
	2386 => "00000000",
	2387 => "00000000",
	2388 => "00000000",
	2389 => "00000000",
	2390 => "00000000",
	2391 => "00000000",
	2392 => "00000000",
	2393 => "00000000",
	2394 => "00000000",
	2395 => "00000000",
	2396 => "00000000",
	2397 => "00000000",
	2398 => "00000000",
	2399 => "00000000",
	2400 => "00000000",
	2401 => "00000000",
	2402 => "00000000",
	2403 => "00000000",
	2404 => "00000000",
	2405 => "00000000",
	2406 => "00000000",
	2407 => "00000000",
	2408 => "00000000",
	2409 => "00000000",
	2410 => "00000000",
	2411 => "00000000",
	2412 => "00000000",
	2413 => "00000000",
	2414 => "00000000",
	2415 => "00000000",
	2416 => "00000000",
	2417 => "00000000",
	2418 => "00000000",
	2419 => "00000000",
	2420 => "00000000",
	2421 => "00000000",
	2422 => "00000000",
	2423 => "00000000",
	2424 => "00000000",
	2425 => "00000000",
	2426 => "00000000",
	2427 => "00000000",
	2432 => "00000000",
	2433 => "00000000",
	2434 => "00000000",
	2435 => "00000000",
	2436 => "00000000",
	2437 => "00000000",
	2438 => "00000000",
	2439 => "00000000",
	2440 => "00000000",
	2441 => "00000000",
	2442 => "00000000",
	2443 => "00000000",
	2444 => "00000000",
	2445 => "00000000",
	2446 => "00000000",
	2447 => "00000000",
	2448 => "00000000",
	2449 => "00000000",
	2450 => "00000000",
	2451 => "00000000",
	2452 => "00000000",
	2453 => "00000000",
	2454 => "00000000",
	2455 => "00000000",
	2456 => "00000000",
	2457 => "00000000",
	2458 => "00000000",
	2459 => "00000000",
	2460 => "00000000",
	2461 => "00000000",
	2462 => "00000000",
	2463 => "00000000",
	2464 => "00000000",
	2465 => "00000000",
	2466 => "00000000",
	2467 => "00000000",
	2468 => "00000000",
	2469 => "00000000",
	2470 => "00000000",
	2471 => "00000000",
	2472 => "00000000",
	2473 => "00000000",
	2474 => "00000000",
	2475 => "00000000",
	2476 => "00000000",
	2477 => "00000000",
	2478 => "00000000",
	2479 => "00000000",
	2480 => "00000000",
	2481 => "00000000",
	2482 => "00000000",
	2483 => "00000000",
	2484 => "00000000",
	2485 => "00000000",
	2486 => "00000000",
	2487 => "00000000",
	2488 => "00000000",
	2489 => "00000000",
	2490 => "00000000",
	2491 => "00000000",
	2496 => "00000000",
	2497 => "00000000",
	2498 => "00000000",
	2499 => "00000000",
	2500 => "00000000",
	2501 => "00000000",
	2502 => "00000000",
	2503 => "00000000",
	2504 => "00000000",
	2505 => "00000000",
	2506 => "00000000",
	2507 => "00000000",
	2508 => "00000000",
	2509 => "00000000",
	2510 => "00000000",
	2511 => "00000000",
	2512 => "00000000",
	2513 => "00000000",
	2514 => "00000000",
	2515 => "00000000",
	2516 => "00000000",
	2517 => "00000000",
	2518 => "00000000",
	2519 => "00000000",
	2520 => "00000000",
	2521 => "00000000",
	2522 => "00000000",
	2523 => "00000000",
	2524 => "00000000",
	2525 => "00000000",
	2526 => "00000000",
	2527 => "00000000",
	2528 => "00000000",
	2529 => "00000000",
	2530 => "00000000",
	2531 => "00000000",
	2532 => "00000000",
	2533 => "00000000",
	2534 => "00000000",
	2535 => "00000000",
	2536 => "00000000",
	2537 => "00000000",
	2538 => "00000000",
	2539 => "00000000",
	2540 => "00000000",
	2541 => "00000000",
	2542 => "00000000",
	2543 => "00000000",
	2544 => "00000000",
	2545 => "00000000",
	2546 => "00000000",
	2547 => "00000000",
	2548 => "00000000",
	2549 => "00000000",
	2550 => "00000000",
	2551 => "00000000",
	2552 => "00000000",
	2553 => "00000000",
	2554 => "00000000",
	2555 => "00000000",
	2560 => "00000000",
	2561 => "00000000",
	2562 => "00000000",
	2563 => "00000000",
	2564 => "00000000",
	2565 => "00000000",
	2566 => "00000000",
	2567 => "00000000",
	2568 => "00000000",
	2569 => "00000000",
	2570 => "00000000",
	2571 => "00000000",
	2572 => "00000000",
	2573 => "00000000",
	2574 => "00000000",
	2575 => "00000000",
	2576 => "00000000",
	2577 => "00000000",
	2578 => "00000000",
	2579 => "00000000",
	2580 => "00000000",
	2581 => "00000000",
	2582 => "00000000",
	2583 => "00000000",
	2584 => "00000000",
	2585 => "00000000",
	2586 => "00000000",
	2587 => "00000000",
	2588 => "00000000",
	2589 => "00000000",
	2590 => "00000000",
	2591 => "00000000",
	2592 => "00000000",
	2593 => "00000000",
	2594 => "00000000",
	2595 => "00000000",
	2596 => "00000000",
	2597 => "00000000",
	2598 => "00000000",
	2599 => "00000000",
	2600 => "00000000",
	2601 => "00000000",
	2602 => "00000000",
	2603 => "00000000",
	2604 => "00000000",
	2605 => "00000000",
	2606 => "00000000",
	2607 => "00000000",
	2608 => "00000000",
	2609 => "00000000",
	2610 => "00000000",
	2611 => "00000000",
	2612 => "00000000",
	2613 => "00000000",
	2614 => "00000000",
	2615 => "00000000",
	2616 => "00000000",
	2617 => "00000000",
	2618 => "00000000",
	2619 => "00000000",
	2624 => "00000000",
	2625 => "00000000",
	2626 => "00000000",
	2627 => "00000000",
	2628 => "00000000",
	2629 => "00000000",
	2630 => "00000000",
	2631 => "00000000",
	2632 => "00000000",
	2633 => "00000000",
	2634 => "00000000",
	2635 => "00000000",
	2636 => "00000000",
	2637 => "00000000",
	2638 => "00000000",
	2639 => "00000000",
	2640 => "00000000",
	2641 => "00000000",
	2642 => "00000000",
	2643 => "00000000",
	2644 => "00000000",
	2645 => "00000000",
	2646 => "00000000",
	2647 => "00000000",
	2648 => "00000000",
	2649 => "00000000",
	2650 => "00000000",
	2651 => "00000000",
	2652 => "00000000",
	2653 => "00000000",
	2654 => "00000000",
	2655 => "00000000",
	2656 => "00000000",
	2657 => "00000000",
	2658 => "00000000",
	2659 => "00000000",
	2660 => "00000000",
	2661 => "00000000",
	2662 => "00000000",
	2663 => "00000000",
	2664 => "00000000",
	2665 => "00000000",
	2666 => "00000000",
	2667 => "00000000",
	2668 => "00000000",
	2669 => "00000000",
	2670 => "00000000",
	2671 => "00000000",
	2672 => "00000000",
	2673 => "00000000",
	2674 => "00000000",
	2675 => "00000000",
	2676 => "00000000",
	2677 => "00000000",
	2678 => "00000000",
	2679 => "00000000",
	2680 => "00000000",
	2681 => "00000000",
	2682 => "00000000",
	2683 => "00000000",
	2688 => "00000000",
	2689 => "00000000",
	2690 => "00000000",
	2691 => "00000000",
	2692 => "00000000",
	2693 => "00000000",
	2694 => "00000000",
	2695 => "00000000",
	2696 => "00000000",
	2697 => "00000000",
	2698 => "00000000",
	2699 => "00000000",
	2700 => "00000000",
	2701 => "00000000",
	2702 => "00000000",
	2703 => "00000000",
	2704 => "00000000",
	2705 => "00000000",
	2706 => "00000000",
	2707 => "00000000",
	2708 => "00000000",
	2709 => "00000000",
	2710 => "00000000",
	2711 => "00000000",
	2712 => "00000000",
	2713 => "00000000",
	2714 => "00000000",
	2715 => "00000000",
	2716 => "00000000",
	2717 => "00000000",
	2718 => "00000000",
	2719 => "00000000",
	2720 => "00000000",
	2721 => "00000000",
	2722 => "00000000",
	2723 => "00000000",
	2724 => "00000000",
	2725 => "00000000",
	2726 => "00000000",
	2727 => "00000000",
	2728 => "00000000",
	2729 => "00000000",
	2730 => "00000000",
	2731 => "00000000",
	2732 => "00000000",
	2733 => "00000000",
	2734 => "00000000",
	2735 => "00000000",
	2736 => "00000000",
	2737 => "00000000",
	2738 => "00000000",
	2739 => "00000000",
	2740 => "00000000",
	2741 => "00000000",
	2742 => "00000000",
	2743 => "00000000",
	2744 => "00000000",
	2745 => "00000000",
	2746 => "00000000",
	2747 => "00000000",
	2752 => "00000000",
	2753 => "00000000",
	2754 => "00000000",
	2755 => "00000000",
	2756 => "00000000",
	2757 => "00000000",
	2758 => "00000000",
	2759 => "00000000",
	2760 => "00000000",
	2761 => "00000000",
	2762 => "00000000",
	2763 => "00000000",
	2764 => "00000000",
	2765 => "00000000",
	2766 => "00000000",
	2767 => "00000000",
	2768 => "00000000",
	2769 => "00000000",
	2770 => "00000000",
	2771 => "00000000",
	2772 => "00000000",
	2773 => "00000000",
	2774 => "00000000",
	2775 => "00000000",
	2776 => "00000000",
	2777 => "00000000",
	2778 => "00000000",
	2779 => "00000000",
	2780 => "00000000",
	2781 => "00000000",
	2782 => "00000000",
	2783 => "00000000",
	2784 => "00000000",
	2785 => "00000000",
	2786 => "00000000",
	2787 => "00000000",
	2788 => "00000000",
	2789 => "00000000",
	2790 => "00000000",
	2791 => "00000000",
	2792 => "00000000",
	2793 => "00000000",
	2794 => "00000000",
	2795 => "00000000",
	2796 => "00000000",
	2797 => "00000000",
	2798 => "00000000",
	2799 => "00000000",
	2800 => "00000000",
	2801 => "00000000",
	2802 => "00000000",
	2803 => "00000000",
	2804 => "00000000",
	2805 => "00000000",
	2806 => "00000000",
	2807 => "00000000",
	2808 => "00000000",
	2809 => "00000000",
	2810 => "00000000",
	2811 => "00000000",
	2816 => "00000000",
	2817 => "00000000",
	2818 => "00000000",
	2819 => "00000000",
	2820 => "00000000",
	2821 => "00000000",
	2822 => "00000000",
	2823 => "00000000",
	2824 => "00000000",
	2825 => "00000000",
	2826 => "00000000",
	2827 => "00000000",
	2828 => "00000000",
	2829 => "00000000",
	2830 => "00000000",
	2831 => "00000000",
	2832 => "00000000",
	2833 => "00000000",
	2834 => "00000000",
	2835 => "00000000",
	2836 => "00000000",
	2837 => "00000000",
	2838 => "00000000",
	2839 => "00000000",
	2840 => "00000000",
	2841 => "00000000",
	2842 => "00000000",
	2843 => "00000000",
	2844 => "00000000",
	2845 => "00000000",
	2846 => "00000000",
	2847 => "00000000",
	2848 => "00000000",
	2849 => "00000000",
	2850 => "00000000",
	2851 => "00000000",
	2852 => "00000000",
	2853 => "00000000",
	2854 => "00000000",
	2855 => "00000000",
	2856 => "00000000",
	2857 => "00000000",
	2858 => "00000000",
	2859 => "00000000",
	2860 => "00000000",
	2861 => "00000000",
	2862 => "00000000",
	2863 => "00000000",
	2864 => "00000000",
	2865 => "00000000",
	2866 => "00000000",
	2867 => "00000000",
	2868 => "00000000",
	2869 => "00000000",
	2870 => "00000000",
	2871 => "00000000",
	2872 => "00000000",
	2873 => "00000000",
	2874 => "00000000",
	2875 => "00000000",
	2880 => "00000000",
	2881 => "00000000",
	2882 => "00000000",
	2883 => "00000000",
	2884 => "00000000",
	2885 => "00000000",
	2886 => "00000000",
	2887 => "00000000",
	2888 => "00000000",
	2889 => "00000000",
	2890 => "00000000",
	2891 => "00000000",
	2892 => "00000000",
	2893 => "00000000",
	2894 => "00000000",
	2895 => "00000000",
	2896 => "00000000",
	2897 => "00000000",
	2898 => "00000000",
	2899 => "00000000",
	2900 => "00000000",
	2901 => "00000000",
	2902 => "00000000",
	2903 => "00000000",
	2904 => "00000000",
	2905 => "00000000",
	2906 => "00000000",
	2907 => "00000000",
	2908 => "00000000",
	2909 => "00000000",
	2910 => "00000000",
	2911 => "00000000",
	2912 => "00000000",
	2913 => "00000000",
	2914 => "00000000",
	2915 => "00000000",
	2916 => "00000000",
	2917 => "00000000",
	2918 => "00000000",
	2919 => "00000000",
	2920 => "00000000",
	2921 => "00000000",
	2922 => "00000000",
	2923 => "00000000",
	2924 => "00000000",
	2925 => "00000000",
	2926 => "00000000",
	2927 => "00000000",
	2928 => "00000000",
	2929 => "00000000",
	2930 => "00000000",
	2931 => "00000000",
	2932 => "00000000",
	2933 => "00000000",
	2934 => "00000000",
	2935 => "00000000",
	2936 => "00000000",
	2937 => "00000000",
	2938 => "00000000",
	2939 => "00000000",
	2944 => "00000000",
	2945 => "00000000",
	2946 => "00000000",
	2947 => "00000000",
	2948 => "00000000",
	2949 => "00000000",
	2950 => "00000000",
	2951 => "00000000",
	2952 => "00000000",
	2953 => "00000000",
	2954 => "00000000",
	2955 => "00000000",
	2956 => "00000000",
	2957 => "00000000",
	2958 => "00000000",
	2959 => "00000000",
	2960 => "00000000",
	2961 => "00000000",
	2962 => "00000000",
	2963 => "00000000",
	2964 => "00000000",
	2965 => "00000000",
	2966 => "00000000",
	2967 => "00000000",
	2968 => "00000000",
	2969 => "00000000",
	2970 => "00000000",
	2971 => "00000000",
	2972 => "00000000",
	2973 => "00000000",
	2974 => "00000000",
	2975 => "00000000",
	2976 => "00000000",
	2977 => "00000000",
	2978 => "00000000",
	2979 => "00000000",
	2980 => "00000000",
	2981 => "00000000",
	2982 => "00000000",
	2983 => "00000000",
	2984 => "00000000",
	2985 => "00000000",
	2986 => "00000000",
	2987 => "00000000",
	2988 => "00000000",
	2989 => "00000000",
	2990 => "00000000",
	2991 => "00000000",
	2992 => "00000000",
	2993 => "00000000",
	2994 => "00000000",
	2995 => "00000000",
	2996 => "00000000",
	2997 => "00000000",
	2998 => "00000000",
	2999 => "00000000",
	3000 => "00000000",
	3001 => "00000000",
	3002 => "00000000",
	3003 => "00000000",
	3008 => "00000000",
	3009 => "00000000",
	3010 => "00000000",
	3011 => "00000000",
	3012 => "00000000",
	3013 => "00000000",
	3014 => "00000000",
	3015 => "00000000",
	3016 => "00000000",
	3017 => "00000000",
	3018 => "00000000",
	3019 => "00000000",
	3020 => "00000000",
	3021 => "00000000",
	3022 => "00000000",
	3023 => "00000000",
	3024 => "00000000",
	3025 => "00000000",
	3026 => "00000000",
	3027 => "00000000",
	3028 => "00000000",
	3029 => "00000000",
	3030 => "00000000",
	3031 => "00000000",
	3032 => "00000000",
	3033 => "00000000",
	3034 => "00000000",
	3035 => "00000000",
	3036 => "00000000",
	3037 => "00000000",
	3038 => "00000000",
	3039 => "00000000",
	3040 => "00000000",
	3041 => "00000000",
	3042 => "00000000",
	3043 => "00000000",
	3044 => "00000000",
	3045 => "00000000",
	3046 => "00000000",
	3047 => "00000000",
	3048 => "00000000",
	3049 => "00000000",
	3050 => "00000000",
	3051 => "00000000",
	3052 => "00000000",
	3053 => "00000000",
	3054 => "00000000",
	3055 => "00000000",
	3056 => "00000000",
	3057 => "00000000",
	3058 => "00000000",
	3059 => "00000000",
	3060 => "00000000",
	3061 => "00000000",
	3062 => "00000000",
	3063 => "00000000",
	3064 => "00000000",
	3065 => "00000000",
	3066 => "00000000",
	3067 => "00000000",
	3072 => "00000000",
	3073 => "00000000",
	3074 => "00000000",
	3075 => "00000000",
	3076 => "00000000",
	3077 => "00000000",
	3078 => "00000000",
	3079 => "00000000",
	3080 => "00000000",
	3081 => "00000000",
	3082 => "00000000",
	3083 => "00000000",
	3084 => "00000000",
	3085 => "00000000",
	3086 => "00000000",
	3087 => "00000000",
	3088 => "00000000",
	3089 => "00000000",
	3090 => "00000000",
	3091 => "00000000",
	3092 => "00000000",
	3093 => "00000000",
	3094 => "00000000",
	3095 => "00000000",
	3096 => "00000000",
	3097 => "00000000",
	3098 => "00000000",
	3099 => "00000000",
	3100 => "00000000",
	3101 => "00000000",
	3102 => "00000000",
	3103 => "00000000",
	3104 => "00000000",
	3105 => "00000000",
	3106 => "00000000",
	3107 => "00000000",
	3108 => "00000000",
	3109 => "00000000",
	3110 => "00000000",
	3111 => "00000000",
	3112 => "00000000",
	3113 => "00000000",
	3114 => "00000000",
	3115 => "00000000",
	3116 => "00000000",
	3117 => "00000000",
	3118 => "00000000",
	3119 => "00000000",
	3120 => "00000000",
	3121 => "00000000",
	3122 => "00000000",
	3123 => "00000000",
	3124 => "00000000",
	3125 => "00000000",
	3126 => "00000000",
	3127 => "00000000",
	3128 => "00000000",
	3129 => "00000000",
	3130 => "00000000",
	3131 => "00000000",
	3136 => "00000000",
	3137 => "00000000",
	3138 => "00000000",
	3139 => "00000000",
	3140 => "00000000",
	3141 => "00000000",
	3142 => "00000000",
	3143 => "00000000",
	3144 => "00000000",
	3145 => "00000000",
	3146 => "00000000",
	3147 => "00000000",
	3148 => "00000000",
	3149 => "00000000",
	3150 => "00000000",
	3151 => "00000000",
	3152 => "00000000",
	3153 => "00000000",
	3154 => "00000000",
	3155 => "00000000",
	3156 => "00000000",
	3157 => "00000000",
	3158 => "00000000",
	3159 => "00000000",
	3160 => "00000000",
	3161 => "00000000",
	3162 => "00000000",
	3163 => "00000000",
	3164 => "00000000",
	3165 => "00000000",
	3166 => "00000000",
	3167 => "00000000",
	3168 => "00000000",
	3169 => "00000000",
	3170 => "00000000",
	3171 => "00000000",
	3172 => "00000000",
	3173 => "00000000",
	3174 => "00000000",
	3175 => "00000000",
	3176 => "00000000",
	3177 => "00000000",
	3178 => "00000000",
	3179 => "00000000",
	3180 => "00000000",
	3181 => "00000000",
	3182 => "00000000",
	3183 => "00000000",
	3184 => "00000000",
	3185 => "00000000",
	3186 => "00000000",
	3187 => "00000000",
	3188 => "00000000",
	3189 => "00000000",
	3190 => "00000000",
	3191 => "00000000",
	3192 => "00000000",
	3193 => "00000000",
	3194 => "00000000",
	3195 => "00000000",
	3200 => "00000000",
	3201 => "00000000",
	3202 => "00000000",
	3203 => "00000000",
	3204 => "00000000",
	3205 => "00000000",
	3206 => "00000000",
	3207 => "00000000",
	3208 => "00000000",
	3209 => "00000000",
	3210 => "00000000",
	3211 => "00000000",
	3212 => "00000000",
	3213 => "00000000",
	3214 => "00000000",
	3215 => "00000000",
	3216 => "00000000",
	3217 => "00000000",
	3218 => "00000000",
	3219 => "00000000",
	3220 => "00000000",
	3221 => "00000000",
	3222 => "00000000",
	3223 => "00000000",
	3224 => "00000000",
	3225 => "00000000",
	3226 => "00000000",
	3227 => "00000000",
	3228 => "00000000",
	3229 => "00000000",
	3230 => "00000000",
	3231 => "00000000",
	3232 => "00000000",
	3233 => "00000000",
	3234 => "00000000",
	3235 => "00000000",
	3236 => "00000000",
	3237 => "00000000",
	3238 => "00000000",
	3239 => "00000000",
	3240 => "00000000",
	3241 => "00000000",
	3242 => "00000000",
	3243 => "00000000",
	3244 => "00000000",
	3245 => "00000000",
	3246 => "00000000",
	3247 => "00000000",
	3248 => "00000000",
	3249 => "00000000",
	3250 => "00000000",
	3251 => "00000000",
	3252 => "00000000",
	3253 => "00000000",
	3254 => "00000000",
	3255 => "00000000",
	3256 => "00000000",
	3257 => "00000000",
	3258 => "00000000",
	3259 => "00000000",
	3264 => "00000000",
	3265 => "00000000",
	3266 => "00000000",
	3267 => "00000000",
	3268 => "00000000",
	3269 => "00000000",
	3270 => "00000000",
	3271 => "00000000",
	3272 => "00000000",
	3273 => "00000000",
	3274 => "00000000",
	3275 => "00000000",
	3276 => "00000000",
	3277 => "00000000",
	3278 => "00000000",
	3279 => "00000000",
	3280 => "00000000",
	3281 => "00000000",
	3282 => "00000000",
	3283 => "00000000",
	3284 => "00000000",
	3285 => "00000000",
	3286 => "00000000",
	3287 => "00000000",
	3288 => "00000000",
	3289 => "00000000",
	3290 => "00000000",
	3291 => "00000000",
	3292 => "00000000",
	3293 => "00000000",
	3294 => "00000000",
	3295 => "00000000",
	3296 => "00000000",
	3297 => "00000000",
	3298 => "00000000",
	3299 => "00000000",
	3300 => "00000000",
	3301 => "00000000",
	3302 => "00000000",
	3303 => "00000000",
	3304 => "00000000",
	3305 => "00000000",
	3306 => "00000000",
	3307 => "00000000",
	3308 => "00000000",
	3309 => "00000000",
	3310 => "00000000",
	3311 => "00000000",
	3312 => "00000000",
	3313 => "00000000",
	3314 => "00000000",
	3315 => "00000000",
	3316 => "00000000",
	3317 => "00000000",
	3318 => "00000000",
	3319 => "00000000",
	3320 => "00000000",
	3321 => "00000000",
	3322 => "00000000",
	3323 => "00000000",
	3328 => "00000000",
	3329 => "00000000",
	3330 => "00000000",
	3331 => "00000000",
	3332 => "00000000",
	3333 => "00000000",
	3334 => "00000000",
	3335 => "00000000",
	3336 => "00000000",
	3337 => "00000000",
	3338 => "00000000",
	3339 => "00000000",
	3340 => "00000000",
	3341 => "00000000",
	3342 => "00000000",
	3343 => "00000000",
	3344 => "00000000",
	3345 => "00000000",
	3346 => "00000000",
	3347 => "00000000",
	3348 => "00000000",
	3349 => "00000000",
	3350 => "00000000",
	3351 => "00000000",
	3352 => "00000000",
	3353 => "00000000",
	3354 => "00000000",
	3355 => "00000000",
	3356 => "00000000",
	3357 => "00000000",
	3358 => "00000000",
	3359 => "00000000",
	3360 => "00000000",
	3361 => "00000000",
	3362 => "00000000",
	3363 => "00000000",
	3364 => "00000000",
	3365 => "00000000",
	3366 => "00000000",
	3367 => "00000000",
	3368 => "00000000",
	3369 => "00000000",
	3370 => "00000000",
	3371 => "00000000",
	3372 => "00000000",
	3373 => "00000000",
	3374 => "00000000",
	3375 => "00000000",
	3376 => "00000000",
	3377 => "00000000",
	3378 => "00000000",
	3379 => "00000000",
	3380 => "00000000",
	3381 => "00000000",
	3382 => "00000000",
	3383 => "00000000",
	3384 => "00000000",
	3385 => "00000000",
	3386 => "00000000",
	3387 => "00000000",
	3392 => "00000000",
	3393 => "00000000",
	3394 => "00000000",
	3395 => "00000000",
	3396 => "00000000",
	3397 => "00000000",
	3398 => "00000000",
	3399 => "00000000",
	3400 => "00000000",
	3401 => "00000000",
	3402 => "00000000",
	3403 => "00000000",
	3404 => "00000000",
	3405 => "00000000",
	3406 => "00000000",
	3407 => "00000000",
	3408 => "00000000",
	3409 => "00000000",
	3410 => "00000000",
	3411 => "00000000",
	3412 => "00000000",
	3413 => "00000000",
	3414 => "00000000",
	3415 => "00000000",
	3416 => "00000000",
	3417 => "00000000",
	3418 => "00000000",
	3419 => "00000000",
	3420 => "00000000",
	3421 => "00000000",
	3422 => "00000000",
	3423 => "00000000",
	3424 => "00000000",
	3425 => "00000000",
	3426 => "00000000",
	3427 => "00000000",
	3428 => "00000000",
	3429 => "00000000",
	3430 => "00000000",
	3431 => "00000000",
	3432 => "00000000",
	3433 => "00000000",
	3434 => "00000000",
	3435 => "00000000",
	3436 => "00000000",
	3437 => "00000000",
	3438 => "00000000",
	3439 => "00000000",
	3440 => "00000000",
	3441 => "00000000",
	3442 => "00000000",
	3443 => "00000000",
	3444 => "00000000",
	3445 => "00000000",
	3446 => "00000000",
	3447 => "00000000",
	3448 => "00000000",
	3449 => "00000000",
	3450 => "00000000",
	3451 => "00000000",
	3456 => "00000000",
	3457 => "00000000",
	3458 => "00000000",
	3459 => "00000000",
	3460 => "00000000",
	3461 => "00000000",
	3462 => "00000000",
	3463 => "00000000",
	3464 => "00000000",
	3465 => "00000000",
	3466 => "00000000",
	3467 => "00000000",
	3468 => "00000000",
	3469 => "00000000",
	3470 => "00000000",
	3471 => "00000000",
	3472 => "00000000",
	3473 => "00000000",
	3474 => "00000000",
	3475 => "00000000",
	3476 => "00000000",
	3477 => "00000000",
	3478 => "00000000",
	3479 => "00000000",
	3480 => "00000000",
	3481 => "00000000",
	3482 => "00000000",
	3483 => "00000000",
	3484 => "00000000",
	3485 => "00000000",
	3486 => "00000000",
	3487 => "00000000",
	3488 => "00000000",
	3489 => "00000000",
	3490 => "00000000",
	3491 => "00000000",
	3492 => "00000000",
	3493 => "00000000",
	3494 => "00000000",
	3495 => "00000000",
	3496 => "00000000",
	3497 => "00000000",
	3498 => "00000000",
	3499 => "00000000",
	3500 => "00000000",
	3501 => "00000000",
	3502 => "00000000",
	3503 => "00000000",
	3504 => "00000000",
	3505 => "00000000",
	3506 => "00000000",
	3507 => "00000000",
	3508 => "00000000",
	3509 => "00000000",
	3510 => "00000000",
	3511 => "00000000",
	3512 => "00000000",
	3513 => "00000000",
	3514 => "00000000",
	3515 => "00000000",
	3520 => "00000000",
	3521 => "00000000",
	3522 => "00000000",
	3523 => "00000000",
	3524 => "00000000",
	3525 => "00000000",
	3526 => "00000000",
	3527 => "00000000",
	3528 => "00000000",
	3529 => "00000000",
	3530 => "00000000",
	3531 => "00000000",
	3532 => "00000000",
	3533 => "00000000",
	3534 => "00000000",
	3535 => "00000000",
	3536 => "00000000",
	3537 => "00000000",
	3538 => "00000000",
	3539 => "00000000",
	3540 => "00000000",
	3541 => "00000000",
	3542 => "00000000",
	3543 => "00000000",
	3544 => "00000000",
	3545 => "00000000",
	3546 => "00000000",
	3547 => "00000000",
	3548 => "00000000",
	3549 => "00000000",
	3550 => "00000000",
	3551 => "00000000",
	3552 => "00000000",
	3553 => "00000000",
	3554 => "00000000",
	3555 => "00000000",
	3556 => "00000000",
	3557 => "00000000",
	3558 => "00000000",
	3559 => "00000000",
	3560 => "00000000",
	3561 => "00000000",
	3562 => "00000000",
	3563 => "00000000",
	3564 => "00000000",
	3565 => "00000000",
	3566 => "00000000",
	3567 => "00000000",
	3568 => "00000000",
	3569 => "00000000",
	3570 => "00000000",
	3571 => "00000000",
	3572 => "00000000",
	3573 => "00000000",
	3574 => "00000000",
	3575 => "00000000",
	3576 => "00000000",
	3577 => "00000000",
	3578 => "00000000",
	3579 => "00000000",
	3584 => "00000000",
	3585 => "00000000",
	3586 => "00000000",
	3587 => "00000000",
	3588 => "00000000",
	3589 => "00000000",
	3590 => "00000000",
	3591 => "00000000",
	3592 => "00000000",
	3593 => "00000000",
	3594 => "00000000",
	3595 => "00000000",
	3596 => "00000000",
	3597 => "00000000",
	3598 => "00000000",
	3599 => "00000000",
	3600 => "00000000",
	3601 => "00000000",
	3602 => "00000000",
	3603 => "00000000",
	3604 => "00000000",
	3605 => "00000000",
	3606 => "00000000",
	3607 => "00000000",
	3608 => "00000000",
	3609 => "00000000",
	3610 => "00000000",
	3611 => "00000000",
	3612 => "00000000",
	3613 => "00000000",
	3614 => "00000000",
	3615 => "00000000",
	3616 => "00000000",
	3617 => "00000000",
	3618 => "00000000",
	3619 => "00000000",
	3620 => "00000000",
	3621 => "00000000",
	3622 => "00000000",
	3623 => "00000000",
	3624 => "00000000",
	3625 => "00000000",
	3626 => "00000000",
	3627 => "00000000",
	3628 => "00000000",
	3629 => "00000000",
	3630 => "00000000",
	3631 => "00000000",
	3632 => "00000000",
	3633 => "00000000",
	3634 => "00000000",
	3635 => "00000000",
	3636 => "00000000",
	3637 => "00000000",
	3638 => "00000000",
	3639 => "00000000",
	3640 => "00000000",
	3641 => "00000000",
	3642 => "00000000",
	3643 => "00000000",
	3648 => "00000000",
	3649 => "00000000",
	3650 => "00000000",
	3651 => "00000000",
	3652 => "00000000",
	3653 => "00000000",
	3654 => "00000000",
	3655 => "00000000",
	3656 => "00000000",
	3657 => "00000000",
	3658 => "00000000",
	3659 => "00000000",
	3660 => "00000000",
	3661 => "00000000",
	3662 => "00000000",
	3663 => "00000000",
	3664 => "00000000",
	3665 => "00000000",
	3666 => "00000000",
	3667 => "00000000",
	3668 => "00000000",
	3669 => "00000000",
	3670 => "00000000",
	3671 => "00000000",
	3672 => "00000000",
	3673 => "00000000",
	3674 => "00000000",
	3675 => "00000000",
	3676 => "00000000",
	3677 => "00000000",
	3678 => "00000000",
	3679 => "00000000",
	3680 => "00000000",
	3681 => "00000000",
	3682 => "00000000",
	3683 => "00000000",
	3684 => "00000000",
	3685 => "00000000",
	3686 => "00000000",
	3687 => "00000000",
	3688 => "00000000",
	3689 => "00000000",
	3690 => "00000000",
	3691 => "00000000",
	3692 => "00000000",
	3693 => "00000000",
	3694 => "00000000",
	3695 => "00000000",
	3696 => "00000000",
	3697 => "00000000",
	3698 => "00000000",
	3699 => "00000000",
	3700 => "00000000",
	3701 => "00000000",
	3702 => "00000000",
	3703 => "00000000",
	3704 => "00000000",
	3705 => "00000000",
	3706 => "00000000",
	3707 => "00000000",
	3712 => "00000000",
	3713 => "00000000",
	3714 => "00000000",
	3715 => "00000000",
	3716 => "00000000",
	3717 => "00000000",
	3718 => "00000000",
	3719 => "00000000",
	3720 => "00000000",
	3721 => "00000000",
	3722 => "00000000",
	3723 => "00000000",
	3724 => "00000000",
	3725 => "00000000",
	3726 => "00000000",
	3727 => "00000000",
	3728 => "00000000",
	3729 => "00000000",
	3730 => "00000000",
	3731 => "00000000",
	3732 => "00000000",
	3733 => "00000000",
	3734 => "00000000",
	3735 => "00000000",
	3736 => "00000000",
	3737 => "00000000",
	3738 => "00000000",
	3739 => "00000000",
	3740 => "00000000",
	3741 => "00000000",
	3742 => "00000000",
	3743 => "00000000",
	3744 => "00000000",
	3745 => "00000000",
	3746 => "00000000",
	3747 => "00000000",
	3748 => "00000000",
	3749 => "00000000",
	3750 => "00000000",
	3751 => "00000000",
	3752 => "00000000",
	3753 => "00000000",
	3754 => "00000000",
	3755 => "00000000",
	3756 => "00000000",
	3757 => "00000000",
	3758 => "00000000",
	3759 => "00000000",
	3760 => "00000000",
	3761 => "00000000",
	3762 => "00000000",
	3763 => "00000000",
	3764 => "00000000",
	3765 => "00000000",
	3766 => "00000000",
	3767 => "00000000",
	3768 => "00000000",
	3769 => "00000000",
	3770 => "00000000",
	3771 => "00000000",
	3776 => "00000000",
	3777 => "00000000",
	3778 => "00000000",
	3779 => "00000000",
	3780 => "00000000",
	3781 => "00000000",
	3782 => "00000000",
	3783 => "00000000",
	3784 => "00000000",
	3785 => "00000000",
	3786 => "00000000",
	3787 => "00000000",
	3788 => "00000000",
	3789 => "00000000",
	3790 => "00000000",
	3791 => "00000000",
	3792 => "00000000",
	3793 => "00000000",
	3794 => "00000000",
	3795 => "00000000",
	3796 => "00000000",
	3797 => "00000000",
	3798 => "00000000",
	3799 => "00000000",
	3800 => "00000000",
	3801 => "00000000",
	3802 => "00000000",
	3803 => "00000000",
	3804 => "00000000",
	3805 => "00000000",
	3806 => "00000000",
	3807 => "00000000",
	3808 => "00000000",
	3809 => "00000000",
	3810 => "00000000",
	3811 => "00000000",
	3812 => "00000000",
	3813 => "00000000",
	3814 => "00000000",
	3815 => "00000000",
	3816 => "00000000",
	3817 => "00000000",
	3818 => "00000000",
	3819 => "00000000",
	3820 => "00000000",
	3821 => "00000000",
	3822 => "00000000",
	3823 => "00000000",
	3824 => "00000000",
	3825 => "00000000",
	3826 => "00000000",
	3827 => "00000000",
	3828 => "00000000",
	3829 => "00000000",
	3830 => "00000000",
	3831 => "00000000",
	3832 => "00000000",
	3833 => "00000000",
	3834 => "00000000",
	3835 => "00000000",

	others => (others => '0')
);

begin
	
	-- process ROM
	process (CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (EN = '1') then
				DATA <= ROM(conv_integer(ADDR));
			end if;
		end if;
	end process;
	
end Behavioral;

