		49280 to 49659 => '1',
		50304 to 50683 => '1',
		51328 to 51707 => '1',
		52352 to 52731 => '1',
		53376 to 53755 => '1',
		54400 to 54529 => '1',
		54650 to 54654 => '1',
		54775 to 54779 => '1',
		55424 to 55553 => '1',
		55674 to 55678 => '1',
		55799 to 55803 => '1',
		56448 to 56577 => '1',
		56698 to 56702 => '1',
		56823 to 56827 => '1',
		57472 to 57601 => '1',
		57722 to 57726 => '1',
		57847 to 57851 => '1',
		58496 to 58625 => '1',
		58746 to 58750 => '1',
		58871 to 58875 => '1',
		59520 to 59649 => '1',
		59770 to 59774 => '1',
		59895 to 59899 => '1',
		60544 to 60673 => '1',
		60794 to 60798 => '1',
		60919 to 60923 => '1',
		61568 to 61697 => '1',
		61818 to 61822 => '1',
		61943 to 61947 => '1',
		62592 to 62721 => '1',
		62842 to 62846 => '1',
		62967 to 62971 => '1',
		63616 to 63745 => '1',
		63866 to 63870 => '1',
		63991 to 63995 => '1',
		64640 to 64769 => '1',
		64890 to 64894 => '1',
		65015 to 65019 => '1',
		65664 to 65793 => '1',
		65914 to 65918 => '1',
		66039 to 66043 => '1',
		66688 to 66817 => '1',
		66938 to 66942 => '1',
		67063 to 67067 => '1',
		67712 to 67841 => '1',
		67962 to 67966 => '1',
		68087 to 68091 => '1',
		68736 to 68865 => '1',
		68986 to 68990 => '1',
		69111 to 69115 => '1',
		69760 to 69889 => '1',
		70010 to 70014 => '1',
		70135 to 70139 => '1',
		70784 to 70913 => '1',
		71034 to 71038 => '1',
		71159 to 71163 => '1',
		71808 to 71937 => '1',
		72058 to 72062 => '1',
		72183 to 72187 => '1',
		72832 to 72961 => '1',
		73082 to 73086 => '1',
		73207 to 73211 => '1',
		73856 to 73985 => '1',
		74106 to 74110 => '1',
		74231 to 74235 => '1',
		74880 to 75009 => '1',
		75130 to 75134 => '1',
		75255 to 75259 => '1',
		75904 to 76033 => '1',
		76154 to 76158 => '1',
		76279 to 76283 => '1',
		76928 to 77057 => '1',
		77178 to 77182 => '1',
		77303 to 77307 => '1',
		77952 to 78081 => '1',
		78202 to 78206 => '1',
		78327 to 78331 => '1',
		78976 to 79105 => '1',
		79226 to 79230 => '1',
		79351 to 79355 => '1',
		80000 to 80129 => '1',
		80250 to 80254 => '1',
		80375 to 80379 => '1',
		81024 to 81153 => '1',
		81274 to 81278 => '1',
		81399 to 81403 => '1',
		82048 to 82177 => '1',
		82298 to 82302 => '1',
		82423 to 82427 => '1',
		83072 to 83201 => '1',
		83322 to 83326 => '1',
		83447 to 83451 => '1',
		84096 to 84225 => '1',
		84346 to 84350 => '1',
		84471 to 84475 => '1',
		85120 to 85249 => '1',
		85370 to 85374 => '1',
		85495 to 85499 => '1',
		86144 to 86273 => '1',
		86394 to 86398 => '1',
		86519 to 86523 => '1',
		87168 to 87297 => '1',
		87418 to 87422 => '1',
		87543 to 87547 => '1',
		88192 to 88321 => '1',
		88442 to 88446 => '1',
		88567 to 88571 => '1',
		89216 to 89345 => '1',
		89466 to 89470 => '1',
		89591 to 89595 => '1',
		90240 to 90369 => '1',
		90490 to 90494 => '1',
		90615 to 90619 => '1',
		91264 to 91393 => '1',
		91514 to 91518 => '1',
		91639 to 91643 => '1',
		92288 to 92417 => '1',
		92538 to 92542 => '1',
		92663 to 92667 => '1',
		93312 to 93441 => '1',
		93562 to 93566 => '1',
		93687 to 93691 => '1',
		94336 to 94465 => '1',
		94586 to 94590 => '1',
		94711 to 94715 => '1',
		95360 to 95489 => '1',
		95610 to 95614 => '1',
		95735 to 95739 => '1',
		96384 to 96513 => '1',
		96634 to 96638 => '1',
		96759 to 96763 => '1',
		97408 to 97537 => '1',
		97658 to 97662 => '1',
		97783 to 97787 => '1',
		98432 to 98561 => '1',
		98682 to 98686 => '1',
		98807 to 98811 => '1',
		99456 to 99585 => '1',
		99706 to 99710 => '1',
		99831 to 99835 => '1',
		100480 to 100609 => '1',
		100730 to 100734 => '1',
		100855 to 100859 => '1',
		101504 to 101633 => '1',
		101754 to 101758 => '1',
		101879 to 101883 => '1',
		102528 to 102657 => '1',
		102778 to 102782 => '1',
		102903 to 102907 => '1',
		103552 to 103681 => '1',
		103802 to 103806 => '1',
		103927 to 103931 => '1',
		104576 to 104705 => '1',
		104826 to 104830 => '1',
		104951 to 104955 => '1',
		105600 to 105729 => '1',
		105850 to 105854 => '1',
		105975 to 105979 => '1',
		106624 to 106753 => '1',
		106874 to 106878 => '1',
		106999 to 107003 => '1',
		107648 to 107777 => '1',
		107898 to 107902 => '1',
		108023 to 108027 => '1',
		108672 to 108801 => '1',
		108922 to 108926 => '1',
		109047 to 109051 => '1',
		109696 to 109825 => '1',
		109946 to 109950 => '1',
		110071 to 110075 => '1',
		110720 to 110849 => '1',
		110970 to 110974 => '1',
		111095 to 111099 => '1',
		111744 to 111873 => '1',
		111994 to 111998 => '1',
		112119 to 112123 => '1',
		112768 to 112897 => '1',
		113018 to 113022 => '1',
		113143 to 113147 => '1',
		113792 to 113921 => '1',
		114042 to 114046 => '1',
		114167 to 114171 => '1',
		114816 to 114945 => '1',
		115066 to 115070 => '1',
		115191 to 115195 => '1',
		115840 to 115969 => '1',
		116090 to 116094 => '1',
		116215 to 116219 => '1',
		116864 to 116993 => '1',
		117114 to 117118 => '1',
		117239 to 117243 => '1',
		117888 to 118017 => '1',
		118138 to 118142 => '1',
		118263 to 118267 => '1',
		118912 to 119041 => '1',
		119162 to 119166 => '1',
		119287 to 119291 => '1',
		119936 to 120065 => '1',
		120186 to 120190 => '1',
		120311 to 120315 => '1',
		120960 to 121089 => '1',
		121210 to 121214 => '1',
		121335 to 121339 => '1',
		121984 to 122113 => '1',
		122234 to 122238 => '1',
		122359 to 122363 => '1',
		123008 to 123137 => '1',
		123258 to 123262 => '1',
		123383 to 123387 => '1',
		124032 to 124161 => '1',
		124282 to 124286 => '1',
		124407 to 124411 => '1',
		125056 to 125185 => '1',
		125306 to 125310 => '1',
		125431 to 125435 => '1',
		126080 to 126209 => '1',
		126330 to 126334 => '1',
		126455 to 126459 => '1',
		127104 to 127233 => '1',
		127354 to 127358 => '1',
		127479 to 127483 => '1',
		128128 to 128257 => '1',
		128378 to 128382 => '1',
		128503 to 128507 => '1',
		129152 to 129281 => '1',
		129402 to 129406 => '1',
		129527 to 129531 => '1',
		130176 to 130305 => '1',
		130426 to 130430 => '1',
		130551 to 130555 => '1',
		131200 to 131329 => '1',
		131450 to 131454 => '1',
		131575 to 131579 => '1',
		132224 to 132353 => '1',
		132474 to 132478 => '1',
		132599 to 132603 => '1',
		133248 to 133377 => '1',
		133498 to 133502 => '1',
		133623 to 133627 => '1',
		134272 to 134401 => '1',
		134522 to 134526 => '1',
		134647 to 134651 => '1',
		135296 to 135425 => '1',
		135546 to 135550 => '1',
		135671 to 135675 => '1',
		136320 to 136449 => '1',
		136570 to 136574 => '1',
		136695 to 136699 => '1',
		137344 to 137473 => '1',
		137594 to 137598 => '1',
		137719 to 137723 => '1',
		138368 to 138497 => '1',
		138618 to 138622 => '1',
		138743 to 138747 => '1',
		139392 to 139521 => '1',
		139642 to 139646 => '1',
		139767 to 139771 => '1',
		140416 to 140545 => '1',
		140666 to 140670 => '1',
		140791 to 140795 => '1',
		141440 to 141569 => '1',
		141690 to 141694 => '1',
		141815 to 141819 => '1',
		142464 to 142593 => '1',
		142714 to 142718 => '1',
		142839 to 142843 => '1',
		143488 to 143617 => '1',
		143738 to 143742 => '1',
		143863 to 143867 => '1',
		144512 to 144641 => '1',
		144762 to 144766 => '1',
		144887 to 144891 => '1',
		145536 to 145665 => '1',
		145786 to 145790 => '1',
		145911 to 145915 => '1',
		146560 to 146689 => '1',
		146810 to 146814 => '1',
		146935 to 146939 => '1',
		147584 to 147713 => '1',
		147834 to 147838 => '1',
		147959 to 147963 => '1',
		148608 to 148737 => '1',
		148858 to 148862 => '1',
		148983 to 148987 => '1',
		149632 to 149761 => '1',
		149882 to 149886 => '1',
		150007 to 150011 => '1',
		150656 to 150785 => '1',
		150906 to 150910 => '1',
		151031 to 151035 => '1',
		151680 to 151809 => '1',
		151930 to 151934 => '1',
		152055 to 152059 => '1',
		152704 to 152833 => '1',
		152954 to 152958 => '1',
		153079 to 153083 => '1',
		153728 to 153857 => '1',
		153978 to 153982 => '1',
		154103 to 154107 => '1',
		154752 to 154881 => '1',
		155002 to 155006 => '1',
		155127 to 155131 => '1',
		155776 to 155905 => '1',
		156026 to 156030 => '1',
		156151 to 156155 => '1',
		156800 to 156929 => '1',
		157050 to 157054 => '1',
		157175 to 157179 => '1',
		157824 to 157953 => '1',
		158074 to 158078 => '1',
		158199 to 158203 => '1',
		158848 to 158977 => '1',
		159098 to 159102 => '1',
		159223 to 159227 => '1',
		159872 to 160001 => '1',
		160122 to 160126 => '1',
		160247 to 160251 => '1',
		160896 to 161025 => '1',
		161146 to 161150 => '1',
		161271 to 161275 => '1',
		161920 to 162049 => '1',
		162170 to 162174 => '1',
		162295 to 162299 => '1',
		162944 to 163073 => '1',
		163194 to 163198 => '1',
		163319 to 163323 => '1',
		163968 to 164097 => '1',
		164218 to 164222 => '1',
		164343 to 164347 => '1',
		164992 to 165121 => '1',
		165242 to 165246 => '1',
		165367 to 165371 => '1',
		166016 to 166145 => '1',
		166266 to 166270 => '1',
		166391 to 166395 => '1',
		167040 to 167169 => '1',
		167290 to 167294 => '1',
		167415 to 167419 => '1',
		168064 to 168193 => '1',
		168314 to 168318 => '1',
		168439 to 168443 => '1',
		169088 to 169217 => '1',
		169338 to 169342 => '1',
		169463 to 169467 => '1',
		170112 to 170241 => '1',
		170362 to 170366 => '1',
		170487 to 170491 => '1',
		171136 to 171265 => '1',
		171386 to 171390 => '1',
		171511 to 171515 => '1',
		172160 to 172289 => '1',
		172410 to 172414 => '1',
		172535 to 172539 => '1',
		173184 to 173313 => '1',
		173434 to 173438 => '1',
		173559 to 173563 => '1',
		174208 to 174337 => '1',
		174458 to 174462 => '1',
		174583 to 174587 => '1',
		175232 to 175361 => '1',
		175482 to 175486 => '1',
		175607 to 175611 => '1',
		176256 to 176385 => '1',
		176506 to 176510 => '1',
		176631 to 176635 => '1',
		177280 to 177659 => '1',
		178304 to 178683 => '1',
		179328 to 179707 => '1',
		180352 to 180731 => '1',
		181376 to 181755 => '1',
		182400 to 182404 => '1',
		182525 to 182529 => '1',
		182650 to 182654 => '1',
		182775 to 182779 => '1',
		183424 to 183428 => '1',
		183549 to 183553 => '1',
		183674 to 183678 => '1',
		183799 to 183803 => '1',
		184448 to 184452 => '1',
		184573 to 184577 => '1',
		184698 to 184702 => '1',
		184823 to 184827 => '1',
		185472 to 185476 => '1',
		185597 to 185601 => '1',
		185722 to 185726 => '1',
		185847 to 185851 => '1',
		186496 to 186500 => '1',
		186621 to 186625 => '1',
		186746 to 186750 => '1',
		186871 to 186875 => '1',
		187520 to 187524 => '1',
		187645 to 187649 => '1',
		187770 to 187774 => '1',
		187895 to 187899 => '1',
		188544 to 188548 => '1',
		188669 to 188673 => '1',
		188794 to 188798 => '1',
		188919 to 188923 => '1',
		189568 to 189572 => '1',
		189693 to 189697 => '1',
		189818 to 189822 => '1',
		189943 to 189947 => '1',
		190592 to 190596 => '1',
		190717 to 190721 => '1',
		190842 to 190846 => '1',
		190967 to 190971 => '1',
		191616 to 191620 => '1',
		191741 to 191745 => '1',
		191866 to 191870 => '1',
		191991 to 191995 => '1',
		192640 to 192644 => '1',
		192765 to 192769 => '1',
		192890 to 192894 => '1',
		193015 to 193019 => '1',
		193664 to 193668 => '1',
		193789 to 193793 => '1',
		193914 to 193918 => '1',
		194039 to 194043 => '1',
		194688 to 194692 => '1',
		194813 to 194817 => '1',
		194938 to 194942 => '1',
		195063 to 195067 => '1',
		195712 to 195716 => '1',
		195837 to 195841 => '1',
		195962 to 195966 => '1',
		196087 to 196091 => '1',
		196736 to 196740 => '1',
		196861 to 196865 => '1',
		196986 to 196990 => '1',
		197111 to 197115 => '1',
		197760 to 197764 => '1',
		197885 to 197889 => '1',
		198010 to 198014 => '1',
		198135 to 198139 => '1',
		198784 to 198788 => '1',
		198909 to 198913 => '1',
		199034 to 199038 => '1',
		199159 to 199163 => '1',
		199808 to 199812 => '1',
		199933 to 199937 => '1',
		200058 to 200062 => '1',
		200183 to 200187 => '1',
		200832 to 200836 => '1',
		200957 to 200961 => '1',
		201082 to 201086 => '1',
		201207 to 201211 => '1',
		201856 to 201860 => '1',
		201981 to 201985 => '1',
		202106 to 202110 => '1',
		202231 to 202235 => '1',
		202880 to 202884 => '1',
		203005 to 203009 => '1',
		203130 to 203134 => '1',
		203255 to 203259 => '1',
		203904 to 203908 => '1',
		204029 to 204033 => '1',
		204154 to 204158 => '1',
		204279 to 204283 => '1',
		204928 to 204932 => '1',
		205053 to 205057 => '1',
		205178 to 205182 => '1',
		205303 to 205307 => '1',
		205952 to 205956 => '1',
		206077 to 206081 => '1',
		206202 to 206206 => '1',
		206327 to 206331 => '1',
		206976 to 206980 => '1',
		207101 to 207105 => '1',
		207226 to 207230 => '1',
		207351 to 207355 => '1',
		208000 to 208004 => '1',
		208125 to 208129 => '1',
		208250 to 208254 => '1',
		208375 to 208379 => '1',
		209024 to 209028 => '1',
		209149 to 209153 => '1',
		209274 to 209278 => '1',
		209399 to 209403 => '1',
		210048 to 210052 => '1',
		210173 to 210177 => '1',
		210298 to 210302 => '1',
		210423 to 210427 => '1',
		211072 to 211076 => '1',
		211197 to 211201 => '1',
		211322 to 211326 => '1',
		211447 to 211451 => '1',
		212096 to 212100 => '1',
		212221 to 212225 => '1',
		212346 to 212350 => '1',
		212471 to 212475 => '1',
		213120 to 213124 => '1',
		213245 to 213249 => '1',
		213370 to 213374 => '1',
		213495 to 213499 => '1',
		214144 to 214148 => '1',
		214269 to 214273 => '1',
		214394 to 214398 => '1',
		214519 to 214523 => '1',
		215168 to 215172 => '1',
		215293 to 215297 => '1',
		215418 to 215422 => '1',
		215543 to 215547 => '1',
		216192 to 216196 => '1',
		216317 to 216321 => '1',
		216442 to 216446 => '1',
		216567 to 216571 => '1',
		217216 to 217220 => '1',
		217341 to 217345 => '1',
		217466 to 217470 => '1',
		217591 to 217595 => '1',
		218240 to 218244 => '1',
		218365 to 218369 => '1',
		218490 to 218494 => '1',
		218615 to 218619 => '1',
		219264 to 219268 => '1',
		219389 to 219393 => '1',
		219514 to 219518 => '1',
		219639 to 219643 => '1',
		220288 to 220292 => '1',
		220413 to 220417 => '1',
		220538 to 220542 => '1',
		220663 to 220667 => '1',
		221312 to 221316 => '1',
		221437 to 221441 => '1',
		221562 to 221566 => '1',
		221687 to 221691 => '1',
		222336 to 222340 => '1',
		222461 to 222465 => '1',
		222586 to 222590 => '1',
		222711 to 222715 => '1',
		223360 to 223364 => '1',
		223485 to 223489 => '1',
		223610 to 223614 => '1',
		223735 to 223739 => '1',
		224384 to 224388 => '1',
		224509 to 224513 => '1',
		224634 to 224638 => '1',
		224759 to 224763 => '1',
		225408 to 225412 => '1',
		225533 to 225537 => '1',
		225658 to 225662 => '1',
		225783 to 225787 => '1',
		226432 to 226436 => '1',
		226557 to 226561 => '1',
		226682 to 226686 => '1',
		226807 to 226811 => '1',
		227456 to 227460 => '1',
		227581 to 227585 => '1',
		227706 to 227710 => '1',
		227831 to 227835 => '1',
		228480 to 228484 => '1',
		228605 to 228609 => '1',
		228730 to 228734 => '1',
		228855 to 228859 => '1',
		229504 to 229508 => '1',
		229629 to 229633 => '1',
		229754 to 229758 => '1',
		229879 to 229883 => '1',
		230528 to 230532 => '1',
		230653 to 230657 => '1',
		230778 to 230782 => '1',
		230903 to 230907 => '1',
		231552 to 231556 => '1',
		231677 to 231681 => '1',
		231802 to 231806 => '1',
		231927 to 231931 => '1',
		232576 to 232580 => '1',
		232701 to 232705 => '1',
		232826 to 232830 => '1',
		232951 to 232955 => '1',
		233600 to 233604 => '1',
		233725 to 233729 => '1',
		233850 to 233854 => '1',
		233975 to 233979 => '1',
		234624 to 234628 => '1',
		234749 to 234753 => '1',
		234874 to 234878 => '1',
		234999 to 235003 => '1',
		235648 to 235652 => '1',
		235773 to 235777 => '1',
		235898 to 235902 => '1',
		236023 to 236027 => '1',
		236672 to 236676 => '1',
		236797 to 236801 => '1',
		236922 to 236926 => '1',
		237047 to 237051 => '1',
		237696 to 237700 => '1',
		237821 to 237825 => '1',
		237946 to 237950 => '1',
		238071 to 238075 => '1',
		238720 to 238724 => '1',
		238845 to 238849 => '1',
		238970 to 238974 => '1',
		239095 to 239099 => '1',
		239744 to 239748 => '1',
		239869 to 239873 => '1',
		239994 to 239998 => '1',
		240119 to 240123 => '1',
		240768 to 240772 => '1',
		240893 to 240897 => '1',
		241018 to 241022 => '1',
		241143 to 241147 => '1',
		241792 to 241796 => '1',
		241917 to 241921 => '1',
		242042 to 242046 => '1',
		242167 to 242171 => '1',
		242816 to 242820 => '1',
		242941 to 242945 => '1',
		243066 to 243070 => '1',
		243191 to 243195 => '1',
		243840 to 243844 => '1',
		243965 to 243969 => '1',
		244090 to 244094 => '1',
		244215 to 244219 => '1',
		244864 to 244868 => '1',
		244989 to 244993 => '1',
		245114 to 245118 => '1',
		245239 to 245243 => '1',
		245888 to 245892 => '1',
		246013 to 246017 => '1',
		246138 to 246142 => '1',
		246263 to 246267 => '1',
		246912 to 246916 => '1',
		247037 to 247041 => '1',
		247162 to 247166 => '1',
		247287 to 247291 => '1',
		247936 to 247940 => '1',
		248061 to 248065 => '1',
		248186 to 248190 => '1',
		248311 to 248315 => '1',
		248960 to 248964 => '1',
		249085 to 249089 => '1',
		249210 to 249214 => '1',
		249335 to 249339 => '1',
		249984 to 249988 => '1',
		250109 to 250113 => '1',
		250234 to 250238 => '1',
		250359 to 250363 => '1',
		251008 to 251012 => '1',
		251133 to 251137 => '1',
		251258 to 251262 => '1',
		251383 to 251387 => '1',
		252032 to 252036 => '1',
		252157 to 252161 => '1',
		252282 to 252286 => '1',
		252407 to 252411 => '1',
		253056 to 253060 => '1',
		253181 to 253185 => '1',
		253306 to 253310 => '1',
		253431 to 253435 => '1',
		254080 to 254084 => '1',
		254205 to 254209 => '1',
		254330 to 254334 => '1',
		254455 to 254459 => '1',
		255104 to 255108 => '1',
		255229 to 255233 => '1',
		255354 to 255358 => '1',
		255479 to 255483 => '1',
		256128 to 256132 => '1',
		256253 to 256257 => '1',
		256378 to 256382 => '1',
		256503 to 256507 => '1',
		257152 to 257156 => '1',
		257277 to 257281 => '1',
		257402 to 257406 => '1',
		257527 to 257531 => '1',
		258176 to 258180 => '1',
		258301 to 258305 => '1',
		258426 to 258430 => '1',
		258551 to 258555 => '1',
		259200 to 259204 => '1',
		259325 to 259329 => '1',
		259450 to 259454 => '1',
		259575 to 259579 => '1',
		260224 to 260228 => '1',
		260349 to 260353 => '1',
		260474 to 260478 => '1',
		260599 to 260603 => '1',
		261248 to 261252 => '1',
		261373 to 261377 => '1',
		261498 to 261502 => '1',
		261623 to 261627 => '1',
		262272 to 262276 => '1',
		262397 to 262401 => '1',
		262522 to 262526 => '1',
		262647 to 262651 => '1',
		263296 to 263300 => '1',
		263421 to 263425 => '1',
		263546 to 263550 => '1',
		263671 to 263675 => '1',
		264320 to 264324 => '1',
		264445 to 264449 => '1',
		264570 to 264574 => '1',
		264695 to 264699 => '1',
		265344 to 265348 => '1',
		265469 to 265473 => '1',
		265594 to 265598 => '1',
		265719 to 265723 => '1',
		266368 to 266372 => '1',
		266493 to 266497 => '1',
		266618 to 266622 => '1',
		266743 to 266747 => '1',
		267392 to 267396 => '1',
		267517 to 267521 => '1',
		267642 to 267646 => '1',
		267767 to 267771 => '1',
		268416 to 268420 => '1',
		268541 to 268545 => '1',
		268666 to 268670 => '1',
		268791 to 268795 => '1',
		269440 to 269444 => '1',
		269565 to 269569 => '1',
		269690 to 269694 => '1',
		269815 to 269819 => '1',
		270464 to 270468 => '1',
		270589 to 270593 => '1',
		270714 to 270718 => '1',
		270839 to 270843 => '1',
		271488 to 271492 => '1',
		271613 to 271617 => '1',
		271738 to 271742 => '1',
		271863 to 271867 => '1',
		272512 to 272516 => '1',
		272637 to 272641 => '1',
		272762 to 272766 => '1',
		272887 to 272891 => '1',
		273536 to 273540 => '1',
		273661 to 273665 => '1',
		273786 to 273790 => '1',
		273911 to 273915 => '1',
		274560 to 274564 => '1',
		274685 to 274689 => '1',
		274810 to 274814 => '1',
		274935 to 274939 => '1',
		275584 to 275588 => '1',
		275709 to 275713 => '1',
		275834 to 275838 => '1',
		275959 to 275963 => '1',
		276608 to 276612 => '1',
		276733 to 276737 => '1',
		276858 to 276862 => '1',
		276983 to 276987 => '1',
		277632 to 277636 => '1',
		277757 to 277761 => '1',
		277882 to 277886 => '1',
		278007 to 278011 => '1',
		278656 to 278660 => '1',
		278781 to 278785 => '1',
		278906 to 278910 => '1',
		279031 to 279035 => '1',
		279680 to 279684 => '1',
		279805 to 279809 => '1',
		279930 to 279934 => '1',
		280055 to 280059 => '1',
		280704 to 280708 => '1',
		280829 to 280833 => '1',
		280954 to 280958 => '1',
		281079 to 281083 => '1',
		281728 to 281732 => '1',
		281853 to 281857 => '1',
		281978 to 281982 => '1',
		282103 to 282107 => '1',
		282752 to 282756 => '1',
		282877 to 282881 => '1',
		283002 to 283006 => '1',
		283127 to 283131 => '1',
		283776 to 283780 => '1',
		283901 to 283905 => '1',
		284026 to 284030 => '1',
		284151 to 284155 => '1',
		284800 to 284804 => '1',
		284925 to 284929 => '1',
		285050 to 285054 => '1',
		285175 to 285179 => '1',
		285824 to 285828 => '1',
		285949 to 285953 => '1',
		286074 to 286078 => '1',
		286199 to 286203 => '1',
		286848 to 286852 => '1',
		286973 to 286977 => '1',
		287098 to 287102 => '1',
		287223 to 287227 => '1',
		287872 to 287876 => '1',
		287997 to 288001 => '1',
		288122 to 288126 => '1',
		288247 to 288251 => '1',
		288896 to 288900 => '1',
		289021 to 289025 => '1',
		289146 to 289150 => '1',
		289271 to 289275 => '1',
		289920 to 289924 => '1',
		290045 to 290049 => '1',
		290170 to 290174 => '1',
		290295 to 290299 => '1',
		290944 to 290948 => '1',
		291069 to 291073 => '1',
		291194 to 291198 => '1',
		291319 to 291323 => '1',
		291968 to 291972 => '1',
		292093 to 292097 => '1',
		292218 to 292222 => '1',
		292343 to 292347 => '1',
		292992 to 292996 => '1',
		293117 to 293121 => '1',
		293242 to 293246 => '1',
		293367 to 293371 => '1',
		294016 to 294020 => '1',
		294141 to 294145 => '1',
		294266 to 294270 => '1',
		294391 to 294395 => '1',
		295040 to 295044 => '1',
		295165 to 295169 => '1',
		295290 to 295294 => '1',
		295415 to 295419 => '1',
		296064 to 296068 => '1',
		296189 to 296193 => '1',
		296314 to 296318 => '1',
		296439 to 296443 => '1',
		297088 to 297092 => '1',
		297213 to 297217 => '1',
		297338 to 297342 => '1',
		297463 to 297467 => '1',
		298112 to 298116 => '1',
		298237 to 298241 => '1',
		298362 to 298366 => '1',
		298487 to 298491 => '1',
		299136 to 299140 => '1',
		299261 to 299265 => '1',
		299386 to 299390 => '1',
		299511 to 299515 => '1',
		300160 to 300164 => '1',
		300285 to 300289 => '1',
		300410 to 300414 => '1',
		300535 to 300539 => '1',
		301184 to 301188 => '1',
		301309 to 301313 => '1',
		301434 to 301438 => '1',
		301559 to 301563 => '1',
		302208 to 302212 => '1',
		302333 to 302337 => '1',
		302458 to 302462 => '1',
		302583 to 302587 => '1',
		303232 to 303236 => '1',
		303357 to 303361 => '1',
		303482 to 303486 => '1',
		303607 to 303611 => '1',
		304256 to 304260 => '1',
		304381 to 304385 => '1',
		304506 to 304510 => '1',
		304631 to 304635 => '1',
		305280 to 305659 => '1',
		306304 to 306683 => '1',
		307328 to 307707 => '1',
		308352 to 308731 => '1',
		309376 to 309755 => '1',
		310400 to 310404 => '1',
		310525 to 310529 => '1',
		310650 to 310654 => '1',
		310775 to 310779 => '1',
		311424 to 311428 => '1',
		311549 to 311553 => '1',
		311674 to 311678 => '1',
		311799 to 311803 => '1',
		312448 to 312452 => '1',
		312573 to 312577 => '1',
		312698 to 312702 => '1',
		312823 to 312827 => '1',
		313472 to 313476 => '1',
		313597 to 313601 => '1',
		313722 to 313726 => '1',
		313847 to 313851 => '1',
		314496 to 314500 => '1',
		314621 to 314625 => '1',
		314746 to 314750 => '1',
		314871 to 314875 => '1',
		315520 to 315524 => '1',
		315645 to 315649 => '1',
		315770 to 315774 => '1',
		315895 to 315899 => '1',
		316544 to 316548 => '1',
		316669 to 316673 => '1',
		316794 to 316798 => '1',
		316919 to 316923 => '1',
		317568 to 317572 => '1',
		317693 to 317697 => '1',
		317818 to 317822 => '1',
		317943 to 317947 => '1',
		318592 to 318596 => '1',
		318717 to 318721 => '1',
		318842 to 318846 => '1',
		318967 to 318971 => '1',
		319616 to 319620 => '1',
		319741 to 319745 => '1',
		319866 to 319870 => '1',
		319991 to 319995 => '1',
		320640 to 320644 => '1',
		320765 to 320769 => '1',
		320890 to 320894 => '1',
		321015 to 321019 => '1',
		321664 to 321668 => '1',
		321789 to 321793 => '1',
		321914 to 321918 => '1',
		322039 to 322043 => '1',
		322688 to 322692 => '1',
		322813 to 322817 => '1',
		322938 to 322942 => '1',
		323063 to 323067 => '1',
		323712 to 323716 => '1',
		323837 to 323841 => '1',
		323962 to 323966 => '1',
		324087 to 324091 => '1',
		324736 to 324740 => '1',
		324861 to 324865 => '1',
		324986 to 324990 => '1',
		325111 to 325115 => '1',
		325760 to 325764 => '1',
		325885 to 325889 => '1',
		326010 to 326014 => '1',
		326135 to 326139 => '1',
		326784 to 326788 => '1',
		326909 to 326913 => '1',
		327034 to 327038 => '1',
		327159 to 327163 => '1',
		327808 to 327812 => '1',
		327933 to 327937 => '1',
		328058 to 328062 => '1',
		328183 to 328187 => '1',
		328832 to 328836 => '1',
		328957 to 328961 => '1',
		329082 to 329086 => '1',
		329207 to 329211 => '1',
		329856 to 329860 => '1',
		329981 to 329985 => '1',
		330106 to 330110 => '1',
		330231 to 330235 => '1',
		330880 to 330884 => '1',
		331005 to 331009 => '1',
		331130 to 331134 => '1',
		331255 to 331259 => '1',
		331904 to 331908 => '1',
		332029 to 332033 => '1',
		332154 to 332158 => '1',
		332279 to 332283 => '1',
		332928 to 332932 => '1',
		333053 to 333057 => '1',
		333178 to 333182 => '1',
		333303 to 333307 => '1',
		333952 to 333956 => '1',
		334077 to 334081 => '1',
		334202 to 334206 => '1',
		334327 to 334331 => '1',
		334976 to 334980 => '1',
		335101 to 335105 => '1',
		335226 to 335230 => '1',
		335351 to 335355 => '1',
		336000 to 336004 => '1',
		336125 to 336129 => '1',
		336250 to 336254 => '1',
		336375 to 336379 => '1',
		337024 to 337028 => '1',
		337149 to 337153 => '1',
		337274 to 337278 => '1',
		337399 to 337403 => '1',
		338048 to 338052 => '1',
		338173 to 338177 => '1',
		338298 to 338302 => '1',
		338423 to 338427 => '1',
		339072 to 339076 => '1',
		339197 to 339201 => '1',
		339322 to 339326 => '1',
		339447 to 339451 => '1',
		340096 to 340100 => '1',
		340221 to 340225 => '1',
		340346 to 340350 => '1',
		340471 to 340475 => '1',
		341120 to 341124 => '1',
		341245 to 341249 => '1',
		341370 to 341374 => '1',
		341495 to 341499 => '1',
		342144 to 342148 => '1',
		342269 to 342273 => '1',
		342394 to 342398 => '1',
		342519 to 342523 => '1',
		343168 to 343172 => '1',
		343293 to 343297 => '1',
		343418 to 343422 => '1',
		343543 to 343547 => '1',
		344192 to 344196 => '1',
		344317 to 344321 => '1',
		344442 to 344446 => '1',
		344567 to 344571 => '1',
		345216 to 345220 => '1',
		345341 to 345345 => '1',
		345466 to 345470 => '1',
		345591 to 345595 => '1',
		346240 to 346244 => '1',
		346365 to 346369 => '1',
		346490 to 346494 => '1',
		346615 to 346619 => '1',
		347264 to 347268 => '1',
		347389 to 347393 => '1',
		347514 to 347518 => '1',
		347639 to 347643 => '1',
		348288 to 348292 => '1',
		348413 to 348417 => '1',
		348538 to 348542 => '1',
		348663 to 348667 => '1',
		349312 to 349316 => '1',
		349437 to 349441 => '1',
		349562 to 349566 => '1',
		349687 to 349691 => '1',
		350336 to 350340 => '1',
		350461 to 350465 => '1',
		350586 to 350590 => '1',
		350711 to 350715 => '1',
		351360 to 351364 => '1',
		351485 to 351489 => '1',
		351610 to 351614 => '1',
		351735 to 351739 => '1',
		352384 to 352388 => '1',
		352509 to 352513 => '1',
		352634 to 352638 => '1',
		352759 to 352763 => '1',
		353408 to 353412 => '1',
		353533 to 353537 => '1',
		353658 to 353662 => '1',
		353783 to 353787 => '1',
		354432 to 354436 => '1',
		354557 to 354561 => '1',
		354682 to 354686 => '1',
		354807 to 354811 => '1',
		355456 to 355460 => '1',
		355581 to 355585 => '1',
		355706 to 355710 => '1',
		355831 to 355835 => '1',
		356480 to 356484 => '1',
		356605 to 356609 => '1',
		356730 to 356734 => '1',
		356855 to 356859 => '1',
		357504 to 357508 => '1',
		357629 to 357633 => '1',
		357754 to 357758 => '1',
		357879 to 357883 => '1',
		358528 to 358532 => '1',
		358653 to 358657 => '1',
		358778 to 358782 => '1',
		358903 to 358907 => '1',
		359552 to 359556 => '1',
		359677 to 359681 => '1',
		359802 to 359806 => '1',
		359927 to 359931 => '1',
		360576 to 360580 => '1',
		360701 to 360705 => '1',
		360826 to 360830 => '1',
		360951 to 360955 => '1',
		361600 to 361604 => '1',
		361725 to 361729 => '1',
		361850 to 361854 => '1',
		361975 to 361979 => '1',
		362624 to 362628 => '1',
		362749 to 362753 => '1',
		362874 to 362878 => '1',
		362999 to 363003 => '1',
		363648 to 363652 => '1',
		363773 to 363777 => '1',
		363898 to 363902 => '1',
		364023 to 364027 => '1',
		364672 to 364676 => '1',
		364797 to 364801 => '1',
		364922 to 364926 => '1',
		365047 to 365051 => '1',
		365696 to 365700 => '1',
		365821 to 365825 => '1',
		365946 to 365950 => '1',
		366071 to 366075 => '1',
		366720 to 366724 => '1',
		366845 to 366849 => '1',
		366970 to 366974 => '1',
		367095 to 367099 => '1',
		367744 to 367748 => '1',
		367869 to 367873 => '1',
		367994 to 367998 => '1',
		368119 to 368123 => '1',
		368768 to 368772 => '1',
		368893 to 368897 => '1',
		369018 to 369022 => '1',
		369143 to 369147 => '1',
		369792 to 369796 => '1',
		369917 to 369921 => '1',
		370042 to 370046 => '1',
		370167 to 370171 => '1',
		370816 to 370820 => '1',
		370941 to 370945 => '1',
		371066 to 371070 => '1',
		371191 to 371195 => '1',
		371840 to 371844 => '1',
		371965 to 371969 => '1',
		372090 to 372094 => '1',
		372215 to 372219 => '1',
		372864 to 372868 => '1',
		372989 to 372993 => '1',
		373114 to 373118 => '1',
		373239 to 373243 => '1',
		373888 to 373892 => '1',
		374013 to 374017 => '1',
		374138 to 374142 => '1',
		374263 to 374267 => '1',
		374912 to 374916 => '1',
		375037 to 375041 => '1',
		375162 to 375166 => '1',
		375287 to 375291 => '1',
		375936 to 375940 => '1',
		376061 to 376065 => '1',
		376186 to 376190 => '1',
		376311 to 376315 => '1',
		376960 to 376964 => '1',
		377085 to 377089 => '1',
		377210 to 377214 => '1',
		377335 to 377339 => '1',
		377984 to 377988 => '1',
		378109 to 378113 => '1',
		378234 to 378238 => '1',
		378359 to 378363 => '1',
		379008 to 379012 => '1',
		379133 to 379137 => '1',
		379258 to 379262 => '1',
		379383 to 379387 => '1',
		380032 to 380036 => '1',
		380157 to 380161 => '1',
		380282 to 380286 => '1',
		380407 to 380411 => '1',
		381056 to 381060 => '1',
		381181 to 381185 => '1',
		381306 to 381310 => '1',
		381431 to 381435 => '1',
		382080 to 382084 => '1',
		382205 to 382209 => '1',
		382330 to 382334 => '1',
		382455 to 382459 => '1',
		383104 to 383108 => '1',
		383229 to 383233 => '1',
		383354 to 383358 => '1',
		383479 to 383483 => '1',
		384128 to 384132 => '1',
		384253 to 384257 => '1',
		384378 to 384382 => '1',
		384503 to 384507 => '1',
		385152 to 385156 => '1',
		385277 to 385281 => '1',
		385402 to 385406 => '1',
		385527 to 385531 => '1',
		386176 to 386180 => '1',
		386301 to 386305 => '1',
		386426 to 386430 => '1',
		386551 to 386555 => '1',
		387200 to 387204 => '1',
		387325 to 387329 => '1',
		387450 to 387454 => '1',
		387575 to 387579 => '1',
		388224 to 388228 => '1',
		388349 to 388353 => '1',
		388474 to 388478 => '1',
		388599 to 388603 => '1',
		389248 to 389252 => '1',
		389373 to 389377 => '1',
		389498 to 389502 => '1',
		389623 to 389627 => '1',
		390272 to 390276 => '1',
		390397 to 390401 => '1',
		390522 to 390526 => '1',
		390647 to 390651 => '1',
		391296 to 391300 => '1',
		391421 to 391425 => '1',
		391546 to 391550 => '1',
		391671 to 391675 => '1',
		392320 to 392324 => '1',
		392445 to 392449 => '1',
		392570 to 392574 => '1',
		392695 to 392699 => '1',
		393344 to 393348 => '1',
		393469 to 393473 => '1',
		393594 to 393598 => '1',
		393719 to 393723 => '1',
		394368 to 394372 => '1',
		394493 to 394497 => '1',
		394618 to 394622 => '1',
		394743 to 394747 => '1',
		395392 to 395396 => '1',
		395517 to 395521 => '1',
		395642 to 395646 => '1',
		395767 to 395771 => '1',
		396416 to 396420 => '1',
		396541 to 396545 => '1',
		396666 to 396670 => '1',
		396791 to 396795 => '1',
		397440 to 397444 => '1',
		397565 to 397569 => '1',
		397690 to 397694 => '1',
		397815 to 397819 => '1',
		398464 to 398468 => '1',
		398589 to 398593 => '1',
		398714 to 398718 => '1',
		398839 to 398843 => '1',
		399488 to 399492 => '1',
		399613 to 399617 => '1',
		399738 to 399742 => '1',
		399863 to 399867 => '1',
		400512 to 400516 => '1',
		400637 to 400641 => '1',
		400762 to 400766 => '1',
		400887 to 400891 => '1',
		401536 to 401540 => '1',
		401661 to 401665 => '1',
		401786 to 401790 => '1',
		401911 to 401915 => '1',
		402560 to 402564 => '1',
		402685 to 402689 => '1',
		402810 to 402814 => '1',
		402935 to 402939 => '1',
		403584 to 403588 => '1',
		403709 to 403713 => '1',
		403834 to 403838 => '1',
		403959 to 403963 => '1',
		404608 to 404612 => '1',
		404733 to 404737 => '1',
		404858 to 404862 => '1',
		404983 to 404987 => '1',
		405632 to 405636 => '1',
		405757 to 405761 => '1',
		405882 to 405886 => '1',
		406007 to 406011 => '1',
		406656 to 406660 => '1',
		406781 to 406785 => '1',
		406906 to 406910 => '1',
		407031 to 407035 => '1',
		407680 to 407684 => '1',
		407805 to 407809 => '1',
		407930 to 407934 => '1',
		408055 to 408059 => '1',
		408704 to 408708 => '1',
		408829 to 408833 => '1',
		408954 to 408958 => '1',
		409079 to 409083 => '1',
		409728 to 409732 => '1',
		409853 to 409857 => '1',
		409978 to 409982 => '1',
		410103 to 410107 => '1',
		410752 to 410756 => '1',
		410877 to 410881 => '1',
		411002 to 411006 => '1',
		411127 to 411131 => '1',
		411776 to 411780 => '1',
		411901 to 411905 => '1',
		412026 to 412030 => '1',
		412151 to 412155 => '1',
		412800 to 412804 => '1',
		412925 to 412929 => '1',
		413050 to 413054 => '1',
		413175 to 413179 => '1',
		413824 to 413828 => '1',
		413949 to 413953 => '1',
		414074 to 414078 => '1',
		414199 to 414203 => '1',
		414848 to 414852 => '1',
		414973 to 414977 => '1',
		415098 to 415102 => '1',
		415223 to 415227 => '1',
		415872 to 415876 => '1',
		415997 to 416001 => '1',
		416122 to 416126 => '1',
		416247 to 416251 => '1',
		416896 to 416900 => '1',
		417021 to 417025 => '1',
		417146 to 417150 => '1',
		417271 to 417275 => '1',
		417920 to 417924 => '1',
		418045 to 418049 => '1',
		418170 to 418174 => '1',
		418295 to 418299 => '1',
		418944 to 418948 => '1',
		419069 to 419073 => '1',
		419194 to 419198 => '1',
		419319 to 419323 => '1',
		419968 to 419972 => '1',
		420093 to 420097 => '1',
		420218 to 420222 => '1',
		420343 to 420347 => '1',
		420992 to 420996 => '1',
		421117 to 421121 => '1',
		421242 to 421246 => '1',
		421367 to 421371 => '1',
		422016 to 422020 => '1',
		422141 to 422145 => '1',
		422266 to 422270 => '1',
		422391 to 422395 => '1',
		423040 to 423044 => '1',
		423165 to 423169 => '1',
		423290 to 423294 => '1',
		423415 to 423419 => '1',
		424064 to 424068 => '1',
		424189 to 424193 => '1',
		424314 to 424318 => '1',
		424439 to 424443 => '1',
		425088 to 425092 => '1',
		425213 to 425217 => '1',
		425338 to 425342 => '1',
		425463 to 425467 => '1',
		426112 to 426116 => '1',
		426237 to 426241 => '1',
		426362 to 426366 => '1',
		426487 to 426491 => '1',
		427136 to 427140 => '1',
		427261 to 427265 => '1',
		427386 to 427390 => '1',
		427511 to 427515 => '1',
		428160 to 428164 => '1',
		428285 to 428289 => '1',
		428410 to 428414 => '1',
		428535 to 428539 => '1',
		429184 to 429188 => '1',
		429309 to 429313 => '1',
		429434 to 429438 => '1',
		429559 to 429563 => '1',
		430208 to 430212 => '1',
		430333 to 430337 => '1',
		430458 to 430462 => '1',
		430583 to 430587 => '1',
		431232 to 431236 => '1',
		431357 to 431361 => '1',
		431482 to 431486 => '1',
		431607 to 431611 => '1',
		432256 to 432260 => '1',
		432381 to 432385 => '1',
		432506 to 432510 => '1',
		432631 to 432635 => '1',
		433280 to 433659 => '1',
		434304 to 434683 => '1',
		435328 to 435707 => '1',
		436352 to 436731 => '1',
		437376 to 437755 => '1',
