library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;

entity ROM_O is
	port (CLK : in std_logic;
		  EN : in std_logic;
		  ADDR : in std_logic_vector(13 downto 0);
		  DATA : out std_logic);
end ROM_O;

architecture Behavioral of ROM_O is

type zone_memoire is array ((2**14)-1 downto 0) of std_logic;
constant ROM: zone_memoire := (
		0 => '0',
		1 => '0',
		2 => '0',
		3 => '0',
		4 => '0',
		5 => '0',
		6 => '0',
		7 => '0',
		8 => '0',
		9 => '0',
		10 => '0',
		11 => '0',
		12 => '0',
		13 => '0',
		14 => '0',
		15 => '0',
		16 => '0',
		17 => '0',
		18 => '0',
		19 => '0',
		20 => '0',
		21 => '0',
		22 => '0',
		23 => '0',
		24 => '0',
		25 => '0',
		26 => '0',
		27 => '0',
		28 => '0',
		29 => '0',
		30 => '0',
		31 => '0',
		32 => '0',
		33 => '0',
		34 => '0',
		35 => '0',
		36 => '0',
		37 => '0',
		38 => '0',
		39 => '0',
		40 => '0',
		41 => '0',
		42 => '0',
		43 => '0',
		44 => '0',
		45 => '0',
		46 => '0',
		47 => '0',
		48 => '0',
		49 => '0',
		50 => '0',
		51 => '0',
		52 => '0',
		53 => '0',
		54 => '0',
		55 => '0',
		56 => '0',
		57 => '0',
		58 => '0',
		59 => '0',
		60 => '0',
		61 => '0',
		62 => '0',
		63 => '0',
		64 => '0',
		65 => '0',
		66 => '0',
		67 => '0',
		68 => '0',
		69 => '0',
		70 => '0',
		71 => '0',
		72 => '0',
		73 => '0',
		74 => '0',
		75 => '0',
		76 => '0',
		77 => '0',
		78 => '0',
		79 => '0',
		80 => '0',
		81 => '0',
		82 => '0',
		83 => '0',
		84 => '0',
		85 => '0',
		86 => '0',
		87 => '0',
		88 => '0',
		89 => '0',
		90 => '0',
		91 => '0',
		92 => '0',
		93 => '0',
		94 => '0',
		95 => '0',
		96 => '0',
		97 => '0',
		98 => '0',
		99 => '0',
		100 => '0',
		101 => '0',
		102 => '0',
		103 => '0',
		104 => '0',
		105 => '0',
		106 => '0',
		107 => '0',
		108 => '0',
		109 => '0',
		110 => '0',
		111 => '0',
		112 => '0',
		113 => '0',
		114 => '0',
		115 => '0',
		116 => '0',
		117 => '0',
		118 => '0',
		119 => '0',
		128 => '0',
		129 => '0',
		130 => '0',
		131 => '0',
		132 => '0',
		133 => '0',
		134 => '0',
		135 => '0',
		136 => '0',
		137 => '0',
		138 => '0',
		139 => '0',
		140 => '0',
		141 => '0',
		142 => '0',
		143 => '0',
		144 => '0',
		145 => '0',
		146 => '0',
		147 => '0',
		148 => '0',
		149 => '0',
		150 => '0',
		151 => '0',
		152 => '0',
		153 => '0',
		154 => '0',
		155 => '0',
		156 => '0',
		157 => '0',
		158 => '0',
		159 => '0',
		160 => '0',
		161 => '0',
		162 => '0',
		163 => '0',
		164 => '0',
		165 => '0',
		166 => '0',
		167 => '0',
		168 => '0',
		169 => '0',
		170 => '0',
		171 => '0',
		172 => '0',
		173 => '0',
		174 => '0',
		175 => '0',
		176 => '0',
		177 => '0',
		178 => '0',
		179 => '0',
		180 => '0',
		181 => '0',
		182 => '0',
		183 => '0',
		184 => '0',
		185 => '0',
		186 => '0',
		187 => '0',
		188 => '0',
		189 => '0',
		190 => '0',
		191 => '0',
		192 => '0',
		193 => '0',
		194 => '0',
		195 => '0',
		196 => '0',
		197 => '0',
		198 => '0',
		199 => '0',
		200 => '0',
		201 => '0',
		202 => '0',
		203 => '0',
		204 => '0',
		205 => '0',
		206 => '0',
		207 => '0',
		208 => '0',
		209 => '0',
		210 => '0',
		211 => '0',
		212 => '0',
		213 => '0',
		214 => '0',
		215 => '0',
		216 => '0',
		217 => '0',
		218 => '0',
		219 => '0',
		220 => '0',
		221 => '0',
		222 => '0',
		223 => '0',
		224 => '0',
		225 => '0',
		226 => '0',
		227 => '0',
		228 => '0',
		229 => '0',
		230 => '0',
		231 => '0',
		232 => '0',
		233 => '0',
		234 => '0',
		235 => '0',
		236 => '0',
		237 => '0',
		238 => '0',
		239 => '0',
		240 => '0',
		241 => '0',
		242 => '0',
		243 => '0',
		244 => '0',
		245 => '0',
		246 => '0',
		247 => '0',
		256 => '0',
		257 => '0',
		258 => '0',
		259 => '0',
		260 => '0',
		261 => '0',
		262 => '0',
		263 => '0',
		264 => '0',
		265 => '0',
		266 => '0',
		267 => '0',
		268 => '0',
		269 => '0',
		270 => '0',
		271 => '0',
		272 => '0',
		273 => '0',
		274 => '0',
		275 => '0',
		276 => '0',
		277 => '0',
		278 => '0',
		279 => '0',
		280 => '0',
		281 => '0',
		282 => '0',
		283 => '0',
		284 => '0',
		285 => '0',
		286 => '0',
		287 => '0',
		288 => '0',
		289 => '0',
		290 => '0',
		291 => '0',
		292 => '0',
		293 => '0',
		294 => '0',
		295 => '0',
		296 => '0',
		297 => '0',
		298 => '0',
		299 => '0',
		300 => '0',
		301 => '0',
		302 => '0',
		303 => '0',
		304 => '0',
		305 => '0',
		306 => '0',
		307 => '0',
		308 => '0',
		309 => '0',
		310 => '0',
		311 => '0',
		312 => '0',
		313 => '0',
		314 => '0',
		315 => '0',
		316 => '0',
		317 => '0',
		318 => '0',
		319 => '0',
		320 => '0',
		321 => '0',
		322 => '0',
		323 => '0',
		324 => '0',
		325 => '0',
		326 => '0',
		327 => '0',
		328 => '0',
		329 => '0',
		330 => '0',
		331 => '0',
		332 => '0',
		333 => '0',
		334 => '0',
		335 => '0',
		336 => '0',
		337 => '0',
		338 => '0',
		339 => '0',
		340 => '0',
		341 => '0',
		342 => '0',
		343 => '0',
		344 => '0',
		345 => '0',
		346 => '0',
		347 => '0',
		348 => '0',
		349 => '0',
		350 => '0',
		351 => '0',
		352 => '0',
		353 => '0',
		354 => '0',
		355 => '0',
		356 => '0',
		357 => '0',
		358 => '0',
		359 => '0',
		360 => '0',
		361 => '0',
		362 => '0',
		363 => '0',
		364 => '0',
		365 => '0',
		366 => '0',
		367 => '0',
		368 => '0',
		369 => '0',
		370 => '0',
		371 => '0',
		372 => '0',
		373 => '0',
		374 => '0',
		375 => '0',
		384 => '0',
		385 => '0',
		386 => '0',
		387 => '0',
		388 => '0',
		389 => '0',
		390 => '0',
		391 => '0',
		392 => '0',
		393 => '0',
		394 => '0',
		395 => '0',
		396 => '0',
		397 => '0',
		398 => '0',
		399 => '0',
		400 => '0',
		401 => '0',
		402 => '0',
		403 => '0',
		404 => '0',
		405 => '0',
		406 => '0',
		407 => '0',
		408 => '0',
		409 => '0',
		410 => '0',
		411 => '0',
		412 => '0',
		413 => '0',
		414 => '0',
		415 => '0',
		416 => '0',
		417 => '0',
		418 => '0',
		419 => '0',
		420 => '0',
		421 => '0',
		422 => '0',
		423 => '0',
		424 => '0',
		425 => '0',
		426 => '0',
		427 => '0',
		428 => '0',
		429 => '0',
		430 => '0',
		431 => '0',
		432 => '0',
		433 => '0',
		434 => '0',
		435 => '0',
		436 => '0',
		437 => '0',
		438 => '0',
		439 => '0',
		440 => '0',
		441 => '0',
		442 => '0',
		443 => '0',
		444 => '0',
		445 => '0',
		446 => '0',
		447 => '0',
		448 => '0',
		449 => '0',
		450 => '0',
		451 => '0',
		452 => '0',
		453 => '0',
		454 => '0',
		455 => '0',
		456 => '0',
		457 => '0',
		458 => '0',
		459 => '0',
		460 => '0',
		461 => '0',
		462 => '0',
		463 => '0',
		464 => '0',
		465 => '0',
		466 => '0',
		467 => '0',
		468 => '0',
		469 => '0',
		470 => '0',
		471 => '0',
		472 => '0',
		473 => '0',
		474 => '0',
		475 => '0',
		476 => '0',
		477 => '0',
		478 => '0',
		479 => '0',
		480 => '0',
		481 => '0',
		482 => '0',
		483 => '0',
		484 => '0',
		485 => '0',
		486 => '0',
		487 => '0',
		488 => '0',
		489 => '0',
		490 => '0',
		491 => '0',
		492 => '0',
		493 => '0',
		494 => '0',
		495 => '0',
		496 => '0',
		497 => '0',
		498 => '0',
		499 => '0',
		500 => '0',
		501 => '0',
		502 => '0',
		503 => '0',
		512 => '0',
		513 => '0',
		514 => '0',
		515 => '0',
		516 => '0',
		517 => '0',
		518 => '0',
		519 => '0',
		520 => '0',
		521 => '0',
		522 => '0',
		523 => '0',
		524 => '0',
		525 => '0',
		526 => '0',
		527 => '0',
		528 => '0',
		529 => '0',
		530 => '0',
		531 => '0',
		532 => '0',
		533 => '0',
		534 => '0',
		535 => '0',
		536 => '0',
		537 => '0',
		538 => '0',
		539 => '0',
		540 => '0',
		541 => '0',
		542 => '0',
		543 => '0',
		544 => '0',
		545 => '0',
		546 => '0',
		547 => '0',
		548 => '0',
		549 => '0',
		550 => '0',
		551 => '0',
		552 => '0',
		553 => '0',
		554 => '0',
		555 => '0',
		556 => '0',
		557 => '0',
		558 => '0',
		559 => '0',
		560 => '0',
		561 => '0',
		562 => '0',
		563 => '0',
		564 => '0',
		565 => '0',
		566 => '0',
		567 => '0',
		568 => '0',
		569 => '0',
		570 => '0',
		571 => '0',
		572 => '0',
		573 => '0',
		574 => '0',
		575 => '0',
		576 => '0',
		577 => '0',
		578 => '0',
		579 => '0',
		580 => '0',
		581 => '0',
		582 => '0',
		583 => '0',
		584 => '0',
		585 => '0',
		586 => '0',
		587 => '0',
		588 => '0',
		589 => '0',
		590 => '0',
		591 => '0',
		592 => '0',
		593 => '0',
		594 => '0',
		595 => '0',
		596 => '0',
		597 => '0',
		598 => '0',
		599 => '0',
		600 => '0',
		601 => '0',
		602 => '0',
		603 => '0',
		604 => '0',
		605 => '0',
		606 => '0',
		607 => '0',
		608 => '0',
		609 => '0',
		610 => '0',
		611 => '0',
		612 => '0',
		613 => '0',
		614 => '0',
		615 => '0',
		616 => '0',
		617 => '0',
		618 => '0',
		619 => '0',
		620 => '0',
		621 => '0',
		622 => '0',
		623 => '0',
		624 => '0',
		625 => '0',
		626 => '0',
		627 => '0',
		628 => '0',
		629 => '0',
		630 => '0',
		631 => '0',
		640 => '0',
		641 => '0',
		642 => '0',
		643 => '0',
		644 => '0',
		645 => '0',
		646 => '0',
		647 => '0',
		648 => '0',
		649 => '0',
		650 => '0',
		651 => '0',
		652 => '0',
		653 => '0',
		654 => '0',
		655 => '0',
		656 => '0',
		657 => '0',
		658 => '0',
		659 => '0',
		660 => '0',
		661 => '0',
		662 => '0',
		663 => '0',
		664 => '0',
		665 => '0',
		666 => '0',
		667 => '0',
		668 => '0',
		669 => '0',
		670 => '0',
		671 => '0',
		672 => '0',
		673 => '0',
		674 => '0',
		675 => '0',
		676 => '0',
		677 => '0',
		678 => '0',
		679 => '0',
		680 => '0',
		681 => '0',
		682 => '0',
		683 => '0',
		684 => '0',
		685 => '0',
		686 => '0',
		687 => '0',
		688 => '0',
		689 => '0',
		690 => '0',
		691 => '0',
		692 => '0',
		693 => '0',
		694 => '0',
		695 => '0',
		696 => '0',
		697 => '0',
		698 => '0',
		699 => '0',
		700 => '0',
		701 => '0',
		702 => '0',
		703 => '0',
		704 => '0',
		705 => '0',
		706 => '0',
		707 => '0',
		708 => '0',
		709 => '0',
		710 => '0',
		711 => '0',
		712 => '0',
		713 => '0',
		714 => '0',
		715 => '0',
		716 => '0',
		717 => '0',
		718 => '0',
		719 => '0',
		720 => '0',
		721 => '0',
		722 => '0',
		723 => '0',
		724 => '0',
		725 => '0',
		726 => '0',
		727 => '0',
		728 => '0',
		729 => '0',
		730 => '0',
		731 => '0',
		732 => '0',
		733 => '0',
		734 => '0',
		735 => '0',
		736 => '0',
		737 => '0',
		738 => '0',
		739 => '0',
		740 => '0',
		741 => '0',
		742 => '0',
		743 => '0',
		744 => '0',
		745 => '0',
		746 => '0',
		747 => '0',
		748 => '0',
		749 => '0',
		750 => '0',
		751 => '0',
		752 => '0',
		753 => '0',
		754 => '0',
		755 => '0',
		756 => '0',
		757 => '0',
		758 => '0',
		759 => '0',
		768 => '0',
		769 => '0',
		770 => '0',
		771 => '0',
		772 => '0',
		773 => '0',
		774 => '0',
		775 => '0',
		776 => '0',
		777 => '0',
		778 => '0',
		779 => '0',
		780 => '0',
		781 => '0',
		782 => '0',
		783 => '0',
		784 => '0',
		785 => '0',
		786 => '0',
		787 => '0',
		788 => '0',
		789 => '0',
		790 => '0',
		791 => '0',
		792 => '0',
		793 => '0',
		794 => '0',
		795 => '0',
		796 => '0',
		797 => '0',
		798 => '0',
		799 => '0',
		800 => '0',
		801 => '0',
		802 => '0',
		803 => '0',
		804 => '0',
		805 => '0',
		806 => '0',
		807 => '0',
		808 => '0',
		809 => '0',
		810 => '0',
		811 => '0',
		812 => '0',
		813 => '0',
		814 => '0',
		815 => '0',
		816 => '0',
		817 => '0',
		818 => '0',
		819 => '0',
		820 => '0',
		821 => '0',
		822 => '0',
		823 => '0',
		824 => '0',
		825 => '0',
		826 => '0',
		827 => '0',
		828 => '0',
		829 => '0',
		830 => '0',
		831 => '0',
		832 => '0',
		833 => '0',
		834 => '0',
		835 => '0',
		836 => '0',
		837 => '0',
		838 => '0',
		839 => '0',
		840 => '0',
		841 => '0',
		842 => '0',
		843 => '0',
		844 => '0',
		845 => '0',
		846 => '0',
		847 => '0',
		848 => '0',
		849 => '0',
		850 => '0',
		851 => '0',
		852 => '0',
		853 => '0',
		854 => '0',
		855 => '0',
		856 => '0',
		857 => '0',
		858 => '0',
		859 => '0',
		860 => '0',
		861 => '0',
		862 => '0',
		863 => '0',
		864 => '0',
		865 => '0',
		866 => '0',
		867 => '0',
		868 => '0',
		869 => '0',
		870 => '0',
		871 => '0',
		872 => '0',
		873 => '0',
		874 => '0',
		875 => '0',
		876 => '0',
		877 => '0',
		878 => '0',
		879 => '0',
		880 => '0',
		881 => '0',
		882 => '0',
		883 => '0',
		884 => '0',
		885 => '0',
		886 => '0',
		887 => '0',
		896 => '0',
		897 => '0',
		898 => '0',
		899 => '0',
		900 => '0',
		901 => '0',
		902 => '0',
		903 => '0',
		904 => '0',
		905 => '0',
		906 => '0',
		907 => '0',
		908 => '0',
		909 => '0',
		910 => '0',
		911 => '0',
		912 => '0',
		913 => '0',
		914 => '0',
		915 => '0',
		916 => '0',
		917 => '0',
		918 => '0',
		919 => '0',
		920 => '0',
		921 => '0',
		922 => '0',
		923 => '0',
		924 => '0',
		925 => '0',
		926 => '0',
		927 => '0',
		928 => '0',
		929 => '0',
		930 => '0',
		931 => '0',
		932 => '0',
		933 => '0',
		934 => '0',
		935 => '0',
		936 => '0',
		937 => '0',
		938 => '0',
		939 => '0',
		940 => '0',
		941 => '0',
		942 => '0',
		943 => '0',
		944 => '0',
		945 => '0',
		946 => '0',
		947 => '0',
		948 => '0',
		949 => '0',
		950 => '0',
		951 => '0',
		952 => '0',
		953 => '0',
		954 => '0',
		955 => '0',
		956 => '0',
		957 => '0',
		958 => '0',
		959 => '0',
		960 => '0',
		961 => '0',
		962 => '0',
		963 => '0',
		964 => '0',
		965 => '0',
		966 => '0',
		967 => '0',
		968 => '0',
		969 => '0',
		970 => '0',
		971 => '0',
		972 => '0',
		973 => '0',
		974 => '0',
		975 => '0',
		976 => '0',
		977 => '0',
		978 => '0',
		979 => '0',
		980 => '0',
		981 => '0',
		982 => '0',
		983 => '0',
		984 => '0',
		985 => '0',
		986 => '0',
		987 => '0',
		988 => '0',
		989 => '0',
		990 => '0',
		991 => '0',
		992 => '0',
		993 => '0',
		994 => '0',
		995 => '0',
		996 => '0',
		997 => '0',
		998 => '0',
		999 => '0',
		1000 => '0',
		1001 => '0',
		1002 => '0',
		1003 => '0',
		1004 => '0',
		1005 => '0',
		1006 => '0',
		1007 => '0',
		1008 => '0',
		1009 => '0',
		1010 => '0',
		1011 => '0',
		1012 => '0',
		1013 => '0',
		1014 => '0',
		1015 => '0',
		1024 => '0',
		1025 => '0',
		1026 => '0',
		1027 => '0',
		1028 => '0',
		1029 => '0',
		1030 => '0',
		1031 => '0',
		1032 => '0',
		1033 => '0',
		1034 => '0',
		1035 => '0',
		1036 => '0',
		1037 => '0',
		1038 => '0',
		1039 => '0',
		1040 => '0',
		1041 => '0',
		1042 => '0',
		1043 => '0',
		1044 => '0',
		1045 => '0',
		1046 => '0',
		1047 => '0',
		1048 => '0',
		1049 => '0',
		1050 => '0',
		1051 => '0',
		1052 => '0',
		1053 => '0',
		1054 => '0',
		1055 => '0',
		1056 => '0',
		1057 => '0',
		1058 => '0',
		1059 => '0',
		1060 => '0',
		1061 => '0',
		1062 => '0',
		1063 => '0',
		1064 => '0',
		1065 => '0',
		1066 => '0',
		1067 => '0',
		1068 => '0',
		1069 => '0',
		1070 => '0',
		1071 => '0',
		1072 => '0',
		1073 => '0',
		1074 => '0',
		1075 => '0',
		1076 => '0',
		1077 => '0',
		1078 => '0',
		1079 => '0',
		1080 => '0',
		1081 => '0',
		1082 => '0',
		1083 => '0',
		1084 => '0',
		1085 => '0',
		1086 => '0',
		1087 => '0',
		1088 => '0',
		1089 => '0',
		1090 => '0',
		1091 => '0',
		1092 => '0',
		1093 => '0',
		1094 => '0',
		1095 => '0',
		1096 => '0',
		1097 => '0',
		1098 => '0',
		1099 => '0',
		1100 => '0',
		1101 => '0',
		1102 => '0',
		1103 => '0',
		1104 => '0',
		1105 => '0',
		1106 => '0',
		1107 => '0',
		1108 => '0',
		1109 => '0',
		1110 => '0',
		1111 => '0',
		1112 => '0',
		1113 => '0',
		1114 => '0',
		1115 => '0',
		1116 => '0',
		1117 => '0',
		1118 => '0',
		1119 => '0',
		1120 => '0',
		1121 => '0',
		1122 => '0',
		1123 => '0',
		1124 => '0',
		1125 => '0',
		1126 => '0',
		1127 => '0',
		1128 => '0',
		1129 => '0',
		1130 => '0',
		1131 => '0',
		1132 => '0',
		1133 => '0',
		1134 => '0',
		1135 => '0',
		1136 => '0',
		1137 => '0',
		1138 => '0',
		1139 => '0',
		1140 => '0',
		1141 => '0',
		1142 => '0',
		1143 => '0',
		1152 => '0',
		1153 => '0',
		1154 => '0',
		1155 => '0',
		1156 => '0',
		1157 => '0',
		1158 => '0',
		1159 => '0',
		1160 => '0',
		1161 => '0',
		1162 => '0',
		1163 => '0',
		1164 => '0',
		1165 => '0',
		1166 => '0',
		1167 => '0',
		1168 => '0',
		1169 => '0',
		1170 => '0',
		1171 => '0',
		1172 => '0',
		1173 => '0',
		1174 => '0',
		1175 => '0',
		1176 => '0',
		1177 => '0',
		1178 => '0',
		1179 => '0',
		1180 => '0',
		1181 => '0',
		1182 => '0',
		1183 => '0',
		1184 => '0',
		1185 => '0',
		1186 => '0',
		1187 => '0',
		1188 => '0',
		1189 => '0',
		1190 => '0',
		1191 => '0',
		1192 => '0',
		1193 => '0',
		1194 => '0',
		1195 => '0',
		1196 => '0',
		1197 => '0',
		1198 => '0',
		1199 => '0',
		1200 => '0',
		1201 => '0',
		1202 => '0',
		1203 => '0',
		1204 => '0',
		1205 => '0',
		1206 => '0',
		1207 => '0',
		1208 => '0',
		1209 => '0',
		1210 => '0',
		1211 => '0',
		1212 => '0',
		1213 => '0',
		1214 => '0',
		1215 => '0',
		1216 => '0',
		1217 => '0',
		1218 => '0',
		1219 => '0',
		1220 => '0',
		1221 => '0',
		1222 => '0',
		1223 => '0',
		1224 => '0',
		1225 => '0',
		1226 => '0',
		1227 => '0',
		1228 => '0',
		1229 => '0',
		1230 => '0',
		1231 => '0',
		1232 => '0',
		1233 => '0',
		1234 => '0',
		1235 => '0',
		1236 => '0',
		1237 => '0',
		1238 => '0',
		1239 => '0',
		1240 => '0',
		1241 => '0',
		1242 => '0',
		1243 => '0',
		1244 => '0',
		1245 => '0',
		1246 => '0',
		1247 => '0',
		1248 => '0',
		1249 => '0',
		1250 => '0',
		1251 => '0',
		1252 => '0',
		1253 => '0',
		1254 => '0',
		1255 => '0',
		1256 => '0',
		1257 => '0',
		1258 => '0',
		1259 => '0',
		1260 => '0',
		1261 => '0',
		1262 => '0',
		1263 => '0',
		1264 => '0',
		1265 => '0',
		1266 => '0',
		1267 => '0',
		1268 => '0',
		1269 => '0',
		1270 => '0',
		1271 => '0',
		1280 => '0',
		1281 => '0',
		1282 => '0',
		1283 => '0',
		1284 => '0',
		1285 => '0',
		1286 => '0',
		1287 => '0',
		1288 => '0',
		1289 => '0',
		1290 => '0',
		1291 => '0',
		1292 => '0',
		1293 => '0',
		1294 => '0',
		1295 => '0',
		1296 => '0',
		1297 => '0',
		1298 => '0',
		1299 => '0',
		1300 => '0',
		1301 => '0',
		1302 => '0',
		1303 => '0',
		1304 => '0',
		1305 => '0',
		1306 => '0',
		1307 => '0',
		1308 => '0',
		1309 => '0',
		1310 => '0',
		1311 => '0',
		1312 => '0',
		1313 => '0',
		1314 => '0',
		1315 => '0',
		1316 => '0',
		1317 => '0',
		1318 => '0',
		1319 => '0',
		1320 => '0',
		1321 => '0',
		1322 => '0',
		1323 => '0',
		1324 => '0',
		1325 => '0',
		1326 => '0',
		1327 => '0',
		1328 => '0',
		1329 => '0',
		1330 => '0',
		1331 => '0',
		1332 => '0',
		1333 => '0',
		1334 => '0',
		1335 => '0',
		1336 => '0',
		1337 => '0',
		1338 => '0',
		1339 => '0',
		1340 => '0',
		1341 => '0',
		1342 => '0',
		1343 => '0',
		1344 => '0',
		1345 => '0',
		1346 => '0',
		1347 => '0',
		1348 => '0',
		1349 => '0',
		1350 => '0',
		1351 => '0',
		1352 => '0',
		1353 => '0',
		1354 => '0',
		1355 => '0',
		1356 => '0',
		1357 => '0',
		1358 => '0',
		1359 => '0',
		1360 => '0',
		1361 => '0',
		1362 => '0',
		1363 => '0',
		1364 => '0',
		1365 => '0',
		1366 => '0',
		1367 => '0',
		1368 => '0',
		1369 => '0',
		1370 => '0',
		1371 => '0',
		1372 => '0',
		1373 => '0',
		1374 => '0',
		1375 => '0',
		1376 => '0',
		1377 => '0',
		1378 => '0',
		1379 => '0',
		1380 => '0',
		1381 => '0',
		1382 => '0',
		1383 => '0',
		1384 => '0',
		1385 => '0',
		1386 => '0',
		1387 => '0',
		1388 => '0',
		1389 => '0',
		1390 => '0',
		1391 => '0',
		1392 => '0',
		1393 => '0',
		1394 => '0',
		1395 => '0',
		1396 => '0',
		1397 => '0',
		1398 => '0',
		1399 => '0',
		1408 => '0',
		1409 => '0',
		1410 => '0',
		1411 => '0',
		1412 => '0',
		1413 => '0',
		1414 => '0',
		1415 => '0',
		1416 => '0',
		1417 => '0',
		1418 => '0',
		1419 => '0',
		1420 => '0',
		1421 => '0',
		1422 => '0',
		1423 => '0',
		1424 => '0',
		1425 => '0',
		1426 => '0',
		1427 => '0',
		1428 => '0',
		1429 => '0',
		1430 => '0',
		1431 => '0',
		1432 => '0',
		1433 => '0',
		1434 => '0',
		1435 => '0',
		1436 => '0',
		1437 => '0',
		1438 => '0',
		1439 => '0',
		1440 => '0',
		1441 => '0',
		1442 => '0',
		1443 => '0',
		1444 => '0',
		1445 => '0',
		1446 => '0',
		1447 => '0',
		1448 => '0',
		1449 => '0',
		1450 => '0',
		1451 => '0',
		1452 => '0',
		1453 => '0',
		1454 => '0',
		1455 => '0',
		1456 => '0',
		1457 => '0',
		1458 => '0',
		1459 => '0',
		1460 => '0',
		1461 => '0',
		1462 => '0',
		1463 => '0',
		1464 => '0',
		1465 => '0',
		1466 => '0',
		1467 => '0',
		1468 => '0',
		1469 => '0',
		1470 => '0',
		1471 => '0',
		1472 => '0',
		1473 => '0',
		1474 => '0',
		1475 => '0',
		1476 => '0',
		1477 => '0',
		1478 => '0',
		1479 => '0',
		1480 => '0',
		1481 => '0',
		1482 => '0',
		1483 => '0',
		1484 => '0',
		1485 => '0',
		1486 => '0',
		1487 => '0',
		1488 => '0',
		1489 => '0',
		1490 => '0',
		1491 => '0',
		1492 => '0',
		1493 => '0',
		1494 => '0',
		1495 => '0',
		1496 => '0',
		1497 => '0',
		1498 => '0',
		1499 => '0',
		1500 => '0',
		1501 => '0',
		1502 => '0',
		1503 => '0',
		1504 => '0',
		1505 => '0',
		1506 => '0',
		1507 => '0',
		1508 => '0',
		1509 => '0',
		1510 => '0',
		1511 => '0',
		1512 => '0',
		1513 => '0',
		1514 => '0',
		1515 => '0',
		1516 => '0',
		1517 => '0',
		1518 => '0',
		1519 => '0',
		1520 => '0',
		1521 => '0',
		1522 => '0',
		1523 => '0',
		1524 => '0',
		1525 => '0',
		1526 => '0',
		1527 => '0',
		1536 => '0',
		1537 => '0',
		1538 => '0',
		1539 => '0',
		1540 => '0',
		1541 => '0',
		1542 => '0',
		1543 => '0',
		1544 => '0',
		1545 => '0',
		1546 => '0',
		1547 => '0',
		1548 => '0',
		1549 => '0',
		1550 => '0',
		1551 => '0',
		1552 => '0',
		1553 => '0',
		1554 => '0',
		1555 => '0',
		1556 => '0',
		1557 => '0',
		1558 => '0',
		1559 => '0',
		1560 => '0',
		1561 => '0',
		1562 => '0',
		1563 => '0',
		1564 => '0',
		1565 => '0',
		1566 => '0',
		1567 => '0',
		1568 => '0',
		1569 => '0',
		1570 => '0',
		1571 => '0',
		1572 => '0',
		1573 => '0',
		1574 => '0',
		1575 => '0',
		1576 => '0',
		1577 => '0',
		1578 => '0',
		1579 => '0',
		1580 => '0',
		1581 => '0',
		1582 => '0',
		1583 => '0',
		1584 => '0',
		1585 => '0',
		1586 => '0',
		1587 => '0',
		1588 => '0',
		1589 => '0',
		1590 => '0',
		1591 => '0',
		1592 => '0',
		1593 => '0',
		1594 => '0',
		1595 => '0',
		1596 => '0',
		1597 => '0',
		1598 => '0',
		1599 => '0',
		1600 => '0',
		1601 => '0',
		1602 => '0',
		1603 => '0',
		1604 => '0',
		1605 => '0',
		1606 => '0',
		1607 => '0',
		1608 => '0',
		1609 => '0',
		1610 => '0',
		1611 => '0',
		1612 => '0',
		1613 => '0',
		1614 => '0',
		1615 => '0',
		1616 => '0',
		1617 => '0',
		1618 => '0',
		1619 => '0',
		1620 => '0',
		1621 => '0',
		1622 => '0',
		1623 => '0',
		1624 => '0',
		1625 => '0',
		1626 => '0',
		1627 => '0',
		1628 => '0',
		1629 => '0',
		1630 => '0',
		1631 => '0',
		1632 => '0',
		1633 => '0',
		1634 => '0',
		1635 => '0',
		1636 => '0',
		1637 => '0',
		1638 => '0',
		1639 => '0',
		1640 => '0',
		1641 => '0',
		1642 => '0',
		1643 => '0',
		1644 => '0',
		1645 => '0',
		1646 => '0',
		1647 => '0',
		1648 => '0',
		1649 => '0',
		1650 => '0',
		1651 => '0',
		1652 => '0',
		1653 => '0',
		1654 => '0',
		1655 => '0',
		1664 => '0',
		1665 => '0',
		1666 => '0',
		1667 => '0',
		1668 => '0',
		1669 => '0',
		1670 => '0',
		1671 => '0',
		1672 => '0',
		1673 => '0',
		1674 => '0',
		1675 => '0',
		1676 => '0',
		1677 => '0',
		1678 => '0',
		1679 => '0',
		1680 => '0',
		1681 => '0',
		1682 => '0',
		1683 => '0',
		1684 => '0',
		1685 => '0',
		1686 => '0',
		1687 => '0',
		1688 => '0',
		1689 => '0',
		1690 => '0',
		1691 => '0',
		1692 => '0',
		1693 => '0',
		1694 => '0',
		1695 => '0',
		1696 => '0',
		1697 => '0',
		1698 => '0',
		1699 => '0',
		1700 => '0',
		1701 => '0',
		1702 => '0',
		1703 => '0',
		1704 => '0',
		1705 => '0',
		1706 => '0',
		1707 => '0',
		1708 => '0',
		1709 => '0',
		1710 => '0',
		1711 => '0',
		1712 => '0',
		1713 => '0',
		1714 => '0',
		1715 => '0',
		1716 => '0',
		1717 => '0',
		1718 => '0',
		1719 => '0',
		1720 => '0',
		1721 => '0',
		1722 => '0',
		1723 => '0',
		1724 => '0',
		1725 => '0',
		1726 => '0',
		1727 => '0',
		1728 => '0',
		1729 => '0',
		1730 => '0',
		1731 => '0',
		1732 => '0',
		1733 => '0',
		1734 => '0',
		1735 => '0',
		1736 => '0',
		1737 => '0',
		1738 => '0',
		1739 => '0',
		1740 => '0',
		1741 => '0',
		1742 => '0',
		1743 => '0',
		1744 => '0',
		1745 => '0',
		1746 => '0',
		1747 => '0',
		1748 => '0',
		1749 => '0',
		1750 => '0',
		1751 => '0',
		1752 => '0',
		1753 => '0',
		1754 => '0',
		1755 => '0',
		1756 => '0',
		1757 => '0',
		1758 => '0',
		1759 => '0',
		1760 => '0',
		1761 => '0',
		1762 => '0',
		1763 => '0',
		1764 => '0',
		1765 => '0',
		1766 => '0',
		1767 => '0',
		1768 => '0',
		1769 => '0',
		1770 => '0',
		1771 => '0',
		1772 => '0',
		1773 => '0',
		1774 => '0',
		1775 => '0',
		1776 => '0',
		1777 => '0',
		1778 => '0',
		1779 => '0',
		1780 => '0',
		1781 => '0',
		1782 => '0',
		1783 => '0',
		1792 => '0',
		1793 => '0',
		1794 => '0',
		1795 => '0',
		1796 => '0',
		1797 => '0',
		1798 => '0',
		1799 => '0',
		1800 => '0',
		1801 => '0',
		1802 => '0',
		1803 => '0',
		1804 => '0',
		1805 => '0',
		1806 => '0',
		1807 => '0',
		1808 => '0',
		1809 => '0',
		1810 => '0',
		1811 => '0',
		1812 => '0',
		1813 => '0',
		1814 => '0',
		1815 => '0',
		1816 => '0',
		1817 => '0',
		1818 => '0',
		1819 => '0',
		1820 => '0',
		1821 => '0',
		1822 => '0',
		1823 => '0',
		1824 => '0',
		1825 => '0',
		1826 => '0',
		1827 => '0',
		1828 => '0',
		1829 => '0',
		1830 => '0',
		1831 => '0',
		1832 => '0',
		1833 => '0',
		1834 => '0',
		1835 => '0',
		1836 => '0',
		1837 => '0',
		1838 => '0',
		1839 => '0',
		1840 => '0',
		1841 => '0',
		1842 => '0',
		1843 => '0',
		1844 => '1',
		1845 => '1',
		1846 => '1',
		1847 => '1',
		1848 => '1',
		1849 => '1',
		1850 => '1',
		1851 => '1',
		1852 => '1',
		1853 => '1',
		1854 => '1',
		1855 => '1',
		1856 => '1',
		1857 => '1',
		1858 => '1',
		1859 => '1',
		1860 => '0',
		1861 => '0',
		1862 => '0',
		1863 => '0',
		1864 => '0',
		1865 => '0',
		1866 => '0',
		1867 => '0',
		1868 => '0',
		1869 => '0',
		1870 => '0',
		1871 => '0',
		1872 => '0',
		1873 => '0',
		1874 => '0',
		1875 => '0',
		1876 => '0',
		1877 => '0',
		1878 => '0',
		1879 => '0',
		1880 => '0',
		1881 => '0',
		1882 => '0',
		1883 => '0',
		1884 => '0',
		1885 => '0',
		1886 => '0',
		1887 => '0',
		1888 => '0',
		1889 => '0',
		1890 => '0',
		1891 => '0',
		1892 => '0',
		1893 => '0',
		1894 => '0',
		1895 => '0',
		1896 => '0',
		1897 => '0',
		1898 => '0',
		1899 => '0',
		1900 => '0',
		1901 => '0',
		1902 => '0',
		1903 => '0',
		1904 => '0',
		1905 => '0',
		1906 => '0',
		1907 => '0',
		1908 => '0',
		1909 => '0',
		1910 => '0',
		1911 => '0',
		1920 => '0',
		1921 => '0',
		1922 => '0',
		1923 => '0',
		1924 => '0',
		1925 => '0',
		1926 => '0',
		1927 => '0',
		1928 => '0',
		1929 => '0',
		1930 => '0',
		1931 => '0',
		1932 => '0',
		1933 => '0',
		1934 => '0',
		1935 => '0',
		1936 => '0',
		1937 => '0',
		1938 => '0',
		1939 => '0',
		1940 => '0',
		1941 => '0',
		1942 => '0',
		1943 => '0',
		1944 => '0',
		1945 => '0',
		1946 => '0',
		1947 => '0',
		1948 => '0',
		1949 => '0',
		1950 => '0',
		1951 => '0',
		1952 => '0',
		1953 => '0',
		1954 => '0',
		1955 => '0',
		1956 => '0',
		1957 => '0',
		1958 => '0',
		1959 => '0',
		1960 => '0',
		1961 => '0',
		1962 => '0',
		1963 => '0',
		1964 => '0',
		1965 => '0',
		1966 => '0',
		1967 => '1',
		1968 => '1',
		1969 => '1',
		1970 => '1',
		1971 => '1',
		1972 => '1',
		1973 => '1',
		1974 => '1',
		1975 => '1',
		1976 => '1',
		1977 => '1',
		1978 => '1',
		1979 => '1',
		1980 => '1',
		1981 => '1',
		1982 => '1',
		1983 => '1',
		1984 => '1',
		1985 => '1',
		1986 => '1',
		1987 => '1',
		1988 => '1',
		1989 => '1',
		1990 => '1',
		1991 => '1',
		1992 => '1',
		1993 => '0',
		1994 => '0',
		1995 => '0',
		1996 => '0',
		1997 => '0',
		1998 => '0',
		1999 => '0',
		2000 => '0',
		2001 => '0',
		2002 => '0',
		2003 => '0',
		2004 => '0',
		2005 => '0',
		2006 => '0',
		2007 => '0',
		2008 => '0',
		2009 => '0',
		2010 => '0',
		2011 => '0',
		2012 => '0',
		2013 => '0',
		2014 => '0',
		2015 => '0',
		2016 => '0',
		2017 => '0',
		2018 => '0',
		2019 => '0',
		2020 => '0',
		2021 => '0',
		2022 => '0',
		2023 => '0',
		2024 => '0',
		2025 => '0',
		2026 => '0',
		2027 => '0',
		2028 => '0',
		2029 => '0',
		2030 => '0',
		2031 => '0',
		2032 => '0',
		2033 => '0',
		2034 => '0',
		2035 => '0',
		2036 => '0',
		2037 => '0',
		2038 => '0',
		2039 => '0',
		2048 => '0',
		2049 => '0',
		2050 => '0',
		2051 => '0',
		2052 => '0',
		2053 => '0',
		2054 => '0',
		2055 => '0',
		2056 => '0',
		2057 => '0',
		2058 => '0',
		2059 => '0',
		2060 => '0',
		2061 => '0',
		2062 => '0',
		2063 => '0',
		2064 => '0',
		2065 => '0',
		2066 => '0',
		2067 => '0',
		2068 => '0',
		2069 => '0',
		2070 => '0',
		2071 => '0',
		2072 => '0',
		2073 => '0',
		2074 => '0',
		2075 => '0',
		2076 => '0',
		2077 => '0',
		2078 => '0',
		2079 => '0',
		2080 => '0',
		2081 => '0',
		2082 => '0',
		2083 => '0',
		2084 => '0',
		2085 => '0',
		2086 => '0',
		2087 => '0',
		2088 => '0',
		2089 => '0',
		2090 => '0',
		2091 => '0',
		2092 => '1',
		2093 => '1',
		2094 => '1',
		2095 => '1',
		2096 => '1',
		2097 => '1',
		2098 => '1',
		2099 => '1',
		2100 => '1',
		2101 => '1',
		2102 => '1',
		2103 => '1',
		2104 => '1',
		2105 => '1',
		2106 => '1',
		2107 => '1',
		2108 => '1',
		2109 => '1',
		2110 => '1',
		2111 => '1',
		2112 => '1',
		2113 => '1',
		2114 => '1',
		2115 => '1',
		2116 => '1',
		2117 => '1',
		2118 => '1',
		2119 => '1',
		2120 => '1',
		2121 => '1',
		2122 => '1',
		2123 => '1',
		2124 => '0',
		2125 => '0',
		2126 => '0',
		2127 => '0',
		2128 => '0',
		2129 => '0',
		2130 => '0',
		2131 => '0',
		2132 => '0',
		2133 => '0',
		2134 => '0',
		2135 => '0',
		2136 => '0',
		2137 => '0',
		2138 => '0',
		2139 => '0',
		2140 => '0',
		2141 => '0',
		2142 => '0',
		2143 => '0',
		2144 => '0',
		2145 => '0',
		2146 => '0',
		2147 => '0',
		2148 => '0',
		2149 => '0',
		2150 => '0',
		2151 => '0',
		2152 => '0',
		2153 => '0',
		2154 => '0',
		2155 => '0',
		2156 => '0',
		2157 => '0',
		2158 => '0',
		2159 => '0',
		2160 => '0',
		2161 => '0',
		2162 => '0',
		2163 => '0',
		2164 => '0',
		2165 => '0',
		2166 => '0',
		2167 => '0',
		2176 => '0',
		2177 => '0',
		2178 => '0',
		2179 => '0',
		2180 => '0',
		2181 => '0',
		2182 => '0',
		2183 => '0',
		2184 => '0',
		2185 => '0',
		2186 => '0',
		2187 => '0',
		2188 => '0',
		2189 => '0',
		2190 => '0',
		2191 => '0',
		2192 => '0',
		2193 => '0',
		2194 => '0',
		2195 => '0',
		2196 => '0',
		2197 => '0',
		2198 => '0',
		2199 => '0',
		2200 => '0',
		2201 => '0',
		2202 => '0',
		2203 => '0',
		2204 => '0',
		2205 => '0',
		2206 => '0',
		2207 => '0',
		2208 => '0',
		2209 => '0',
		2210 => '0',
		2211 => '0',
		2212 => '0',
		2213 => '0',
		2214 => '0',
		2215 => '0',
		2216 => '0',
		2217 => '0',
		2218 => '1',
		2219 => '1',
		2220 => '1',
		2221 => '1',
		2222 => '1',
		2223 => '1',
		2224 => '1',
		2225 => '1',
		2226 => '1',
		2227 => '1',
		2228 => '1',
		2229 => '1',
		2230 => '1',
		2231 => '1',
		2232 => '1',
		2233 => '1',
		2234 => '1',
		2235 => '1',
		2236 => '1',
		2237 => '1',
		2238 => '1',
		2239 => '1',
		2240 => '1',
		2241 => '1',
		2242 => '1',
		2243 => '1',
		2244 => '1',
		2245 => '1',
		2246 => '1',
		2247 => '1',
		2248 => '1',
		2249 => '1',
		2250 => '1',
		2251 => '1',
		2252 => '1',
		2253 => '1',
		2254 => '0',
		2255 => '0',
		2256 => '0',
		2257 => '0',
		2258 => '0',
		2259 => '0',
		2260 => '0',
		2261 => '0',
		2262 => '0',
		2263 => '0',
		2264 => '0',
		2265 => '0',
		2266 => '0',
		2267 => '0',
		2268 => '0',
		2269 => '0',
		2270 => '0',
		2271 => '0',
		2272 => '0',
		2273 => '0',
		2274 => '0',
		2275 => '0',
		2276 => '0',
		2277 => '0',
		2278 => '0',
		2279 => '0',
		2280 => '0',
		2281 => '0',
		2282 => '0',
		2283 => '0',
		2284 => '0',
		2285 => '0',
		2286 => '0',
		2287 => '0',
		2288 => '0',
		2289 => '0',
		2290 => '0',
		2291 => '0',
		2292 => '0',
		2293 => '0',
		2294 => '0',
		2295 => '0',
		2304 => '0',
		2305 => '0',
		2306 => '0',
		2307 => '0',
		2308 => '0',
		2309 => '0',
		2310 => '0',
		2311 => '0',
		2312 => '0',
		2313 => '0',
		2314 => '0',
		2315 => '0',
		2316 => '0',
		2317 => '0',
		2318 => '0',
		2319 => '0',
		2320 => '0',
		2321 => '0',
		2322 => '0',
		2323 => '0',
		2324 => '0',
		2325 => '0',
		2326 => '0',
		2327 => '0',
		2328 => '0',
		2329 => '0',
		2330 => '0',
		2331 => '0',
		2332 => '0',
		2333 => '0',
		2334 => '0',
		2335 => '0',
		2336 => '0',
		2337 => '0',
		2338 => '0',
		2339 => '0',
		2340 => '0',
		2341 => '0',
		2342 => '0',
		2343 => '0',
		2344 => '1',
		2345 => '1',
		2346 => '1',
		2347 => '1',
		2348 => '1',
		2349 => '1',
		2350 => '1',
		2351 => '1',
		2352 => '1',
		2353 => '1',
		2354 => '1',
		2355 => '1',
		2356 => '1',
		2357 => '1',
		2358 => '1',
		2359 => '1',
		2360 => '1',
		2361 => '1',
		2362 => '1',
		2363 => '1',
		2364 => '1',
		2365 => '1',
		2366 => '1',
		2367 => '1',
		2368 => '1',
		2369 => '1',
		2370 => '1',
		2371 => '1',
		2372 => '1',
		2373 => '1',
		2374 => '1',
		2375 => '1',
		2376 => '1',
		2377 => '1',
		2378 => '1',
		2379 => '1',
		2380 => '1',
		2381 => '1',
		2382 => '1',
		2383 => '1',
		2384 => '0',
		2385 => '0',
		2386 => '0',
		2387 => '0',
		2388 => '0',
		2389 => '0',
		2390 => '0',
		2391 => '0',
		2392 => '0',
		2393 => '0',
		2394 => '0',
		2395 => '0',
		2396 => '0',
		2397 => '0',
		2398 => '0',
		2399 => '0',
		2400 => '0',
		2401 => '0',
		2402 => '0',
		2403 => '0',
		2404 => '0',
		2405 => '0',
		2406 => '0',
		2407 => '0',
		2408 => '0',
		2409 => '0',
		2410 => '0',
		2411 => '0',
		2412 => '0',
		2413 => '0',
		2414 => '0',
		2415 => '0',
		2416 => '0',
		2417 => '0',
		2418 => '0',
		2419 => '0',
		2420 => '0',
		2421 => '0',
		2422 => '0',
		2423 => '0',
		2432 => '0',
		2433 => '0',
		2434 => '0',
		2435 => '0',
		2436 => '0',
		2437 => '0',
		2438 => '0',
		2439 => '0',
		2440 => '0',
		2441 => '0',
		2442 => '0',
		2443 => '0',
		2444 => '0',
		2445 => '0',
		2446 => '0',
		2447 => '0',
		2448 => '0',
		2449 => '0',
		2450 => '0',
		2451 => '0',
		2452 => '0',
		2453 => '0',
		2454 => '0',
		2455 => '0',
		2456 => '0',
		2457 => '0',
		2458 => '0',
		2459 => '0',
		2460 => '0',
		2461 => '0',
		2462 => '0',
		2463 => '0',
		2464 => '0',
		2465 => '0',
		2466 => '0',
		2467 => '0',
		2468 => '0',
		2469 => '0',
		2470 => '1',
		2471 => '1',
		2472 => '1',
		2473 => '1',
		2474 => '1',
		2475 => '1',
		2476 => '1',
		2477 => '1',
		2478 => '1',
		2479 => '1',
		2480 => '1',
		2481 => '1',
		2482 => '1',
		2483 => '1',
		2484 => '1',
		2485 => '1',
		2486 => '1',
		2487 => '1',
		2488 => '1',
		2489 => '1',
		2490 => '1',
		2491 => '1',
		2492 => '1',
		2493 => '1',
		2494 => '1',
		2495 => '1',
		2496 => '1',
		2497 => '1',
		2498 => '1',
		2499 => '1',
		2500 => '1',
		2501 => '1',
		2502 => '1',
		2503 => '1',
		2504 => '1',
		2505 => '1',
		2506 => '1',
		2507 => '1',
		2508 => '1',
		2509 => '1',
		2510 => '1',
		2511 => '1',
		2512 => '1',
		2513 => '1',
		2514 => '0',
		2515 => '0',
		2516 => '0',
		2517 => '0',
		2518 => '0',
		2519 => '0',
		2520 => '0',
		2521 => '0',
		2522 => '0',
		2523 => '0',
		2524 => '0',
		2525 => '0',
		2526 => '0',
		2527 => '0',
		2528 => '0',
		2529 => '0',
		2530 => '0',
		2531 => '0',
		2532 => '0',
		2533 => '0',
		2534 => '0',
		2535 => '0',
		2536 => '0',
		2537 => '0',
		2538 => '0',
		2539 => '0',
		2540 => '0',
		2541 => '0',
		2542 => '0',
		2543 => '0',
		2544 => '0',
		2545 => '0',
		2546 => '0',
		2547 => '0',
		2548 => '0',
		2549 => '0',
		2550 => '0',
		2551 => '0',
		2560 => '0',
		2561 => '0',
		2562 => '0',
		2563 => '0',
		2564 => '0',
		2565 => '0',
		2566 => '0',
		2567 => '0',
		2568 => '0',
		2569 => '0',
		2570 => '0',
		2571 => '0',
		2572 => '0',
		2573 => '0',
		2574 => '0',
		2575 => '0',
		2576 => '0',
		2577 => '0',
		2578 => '0',
		2579 => '0',
		2580 => '0',
		2581 => '0',
		2582 => '0',
		2583 => '0',
		2584 => '0',
		2585 => '0',
		2586 => '0',
		2587 => '0',
		2588 => '0',
		2589 => '0',
		2590 => '0',
		2591 => '0',
		2592 => '0',
		2593 => '0',
		2594 => '0',
		2595 => '0',
		2596 => '1',
		2597 => '1',
		2598 => '1',
		2599 => '1',
		2600 => '1',
		2601 => '1',
		2602 => '1',
		2603 => '1',
		2604 => '1',
		2605 => '1',
		2606 => '1',
		2607 => '1',
		2608 => '1',
		2609 => '1',
		2610 => '1',
		2611 => '1',
		2612 => '1',
		2613 => '1',
		2614 => '0',
		2615 => '0',
		2616 => '0',
		2617 => '0',
		2618 => '0',
		2619 => '0',
		2620 => '0',
		2621 => '0',
		2622 => '0',
		2623 => '0',
		2624 => '0',
		2625 => '0',
		2626 => '1',
		2627 => '1',
		2628 => '1',
		2629 => '1',
		2630 => '1',
		2631 => '1',
		2632 => '1',
		2633 => '1',
		2634 => '1',
		2635 => '1',
		2636 => '1',
		2637 => '1',
		2638 => '1',
		2639 => '1',
		2640 => '1',
		2641 => '1',
		2642 => '1',
		2643 => '1',
		2644 => '0',
		2645 => '0',
		2646 => '0',
		2647 => '0',
		2648 => '0',
		2649 => '0',
		2650 => '0',
		2651 => '0',
		2652 => '0',
		2653 => '0',
		2654 => '0',
		2655 => '0',
		2656 => '0',
		2657 => '0',
		2658 => '0',
		2659 => '0',
		2660 => '0',
		2661 => '0',
		2662 => '0',
		2663 => '0',
		2664 => '0',
		2665 => '0',
		2666 => '0',
		2667 => '0',
		2668 => '0',
		2669 => '0',
		2670 => '0',
		2671 => '0',
		2672 => '0',
		2673 => '0',
		2674 => '0',
		2675 => '0',
		2676 => '0',
		2677 => '0',
		2678 => '0',
		2679 => '0',
		2688 => '0',
		2689 => '0',
		2690 => '0',
		2691 => '0',
		2692 => '0',
		2693 => '0',
		2694 => '0',
		2695 => '0',
		2696 => '0',
		2697 => '0',
		2698 => '0',
		2699 => '0',
		2700 => '0',
		2701 => '0',
		2702 => '0',
		2703 => '0',
		2704 => '0',
		2705 => '0',
		2706 => '0',
		2707 => '0',
		2708 => '0',
		2709 => '0',
		2710 => '0',
		2711 => '0',
		2712 => '0',
		2713 => '0',
		2714 => '0',
		2715 => '0',
		2716 => '0',
		2717 => '0',
		2718 => '0',
		2719 => '0',
		2720 => '0',
		2721 => '0',
		2722 => '1',
		2723 => '1',
		2724 => '1',
		2725 => '1',
		2726 => '1',
		2727 => '1',
		2728 => '1',
		2729 => '1',
		2730 => '1',
		2731 => '1',
		2732 => '1',
		2733 => '1',
		2734 => '1',
		2735 => '1',
		2736 => '1',
		2737 => '0',
		2738 => '0',
		2739 => '0',
		2740 => '0',
		2741 => '0',
		2742 => '0',
		2743 => '0',
		2744 => '0',
		2745 => '0',
		2746 => '0',
		2747 => '0',
		2748 => '0',
		2749 => '0',
		2750 => '0',
		2751 => '0',
		2752 => '0',
		2753 => '0',
		2754 => '0',
		2755 => '0',
		2756 => '0',
		2757 => '0',
		2758 => '0',
		2759 => '1',
		2760 => '1',
		2761 => '1',
		2762 => '1',
		2763 => '1',
		2764 => '1',
		2765 => '1',
		2766 => '1',
		2767 => '1',
		2768 => '1',
		2769 => '1',
		2770 => '1',
		2771 => '1',
		2772 => '1',
		2773 => '1',
		2774 => '0',
		2775 => '0',
		2776 => '0',
		2777 => '0',
		2778 => '0',
		2779 => '0',
		2780 => '0',
		2781 => '0',
		2782 => '0',
		2783 => '0',
		2784 => '0',
		2785 => '0',
		2786 => '0',
		2787 => '0',
		2788 => '0',
		2789 => '0',
		2790 => '0',
		2791 => '0',
		2792 => '0',
		2793 => '0',
		2794 => '0',
		2795 => '0',
		2796 => '0',
		2797 => '0',
		2798 => '0',
		2799 => '0',
		2800 => '0',
		2801 => '0',
		2802 => '0',
		2803 => '0',
		2804 => '0',
		2805 => '0',
		2806 => '0',
		2807 => '0',
		2816 => '0',
		2817 => '0',
		2818 => '0',
		2819 => '0',
		2820 => '0',
		2821 => '0',
		2822 => '0',
		2823 => '0',
		2824 => '0',
		2825 => '0',
		2826 => '0',
		2827 => '0',
		2828 => '0',
		2829 => '0',
		2830 => '0',
		2831 => '0',
		2832 => '0',
		2833 => '0',
		2834 => '0',
		2835 => '0',
		2836 => '0',
		2837 => '0',
		2838 => '0',
		2839 => '0',
		2840 => '0',
		2841 => '0',
		2842 => '0',
		2843 => '0',
		2844 => '0',
		2845 => '0',
		2846 => '0',
		2847 => '0',
		2848 => '0',
		2849 => '1',
		2850 => '1',
		2851 => '1',
		2852 => '1',
		2853 => '1',
		2854 => '1',
		2855 => '1',
		2856 => '1',
		2857 => '1',
		2858 => '1',
		2859 => '1',
		2860 => '1',
		2861 => '1',
		2862 => '0',
		2863 => '0',
		2864 => '0',
		2865 => '0',
		2866 => '0',
		2867 => '0',
		2868 => '0',
		2869 => '0',
		2870 => '0',
		2871 => '1',
		2872 => '1',
		2873 => '1',
		2874 => '1',
		2875 => '1',
		2876 => '1',
		2877 => '1',
		2878 => '1',
		2879 => '1',
		2880 => '1',
		2881 => '1',
		2882 => '1',
		2883 => '0',
		2884 => '0',
		2885 => '0',
		2886 => '0',
		2887 => '0',
		2888 => '0',
		2889 => '0',
		2890 => '1',
		2891 => '1',
		2892 => '1',
		2893 => '1',
		2894 => '1',
		2895 => '1',
		2896 => '1',
		2897 => '1',
		2898 => '1',
		2899 => '1',
		2900 => '1',
		2901 => '1',
		2902 => '1',
		2903 => '0',
		2904 => '0',
		2905 => '0',
		2906 => '0',
		2907 => '0',
		2908 => '0',
		2909 => '0',
		2910 => '0',
		2911 => '0',
		2912 => '0',
		2913 => '0',
		2914 => '0',
		2915 => '0',
		2916 => '0',
		2917 => '0',
		2918 => '0',
		2919 => '0',
		2920 => '0',
		2921 => '0',
		2922 => '0',
		2923 => '0',
		2924 => '0',
		2925 => '0',
		2926 => '0',
		2927 => '0',
		2928 => '0',
		2929 => '0',
		2930 => '0',
		2931 => '0',
		2932 => '0',
		2933 => '0',
		2934 => '0',
		2935 => '0',
		2944 => '0',
		2945 => '0',
		2946 => '0',
		2947 => '0',
		2948 => '0',
		2949 => '0',
		2950 => '0',
		2951 => '0',
		2952 => '0',
		2953 => '0',
		2954 => '0',
		2955 => '0',
		2956 => '0',
		2957 => '0',
		2958 => '0',
		2959 => '0',
		2960 => '0',
		2961 => '0',
		2962 => '0',
		2963 => '0',
		2964 => '0',
		2965 => '0',
		2966 => '0',
		2967 => '0',
		2968 => '0',
		2969 => '0',
		2970 => '0',
		2971 => '0',
		2972 => '0',
		2973 => '0',
		2974 => '0',
		2975 => '1',
		2976 => '1',
		2977 => '1',
		2978 => '1',
		2979 => '1',
		2980 => '1',
		2981 => '1',
		2982 => '1',
		2983 => '1',
		2984 => '1',
		2985 => '1',
		2986 => '1',
		2987 => '1',
		2988 => '0',
		2989 => '0',
		2990 => '0',
		2991 => '0',
		2992 => '0',
		2993 => '0',
		2994 => '1',
		2995 => '1',
		2996 => '1',
		2997 => '1',
		2998 => '1',
		2999 => '1',
		3000 => '1',
		3001 => '1',
		3002 => '1',
		3003 => '1',
		3004 => '1',
		3005 => '1',
		3006 => '1',
		3007 => '1',
		3008 => '1',
		3009 => '1',
		3010 => '1',
		3011 => '1',
		3012 => '1',
		3013 => '1',
		3014 => '1',
		3015 => '1',
		3016 => '0',
		3017 => '0',
		3018 => '0',
		3019 => '0',
		3020 => '1',
		3021 => '1',
		3022 => '1',
		3023 => '1',
		3024 => '1',
		3025 => '1',
		3026 => '1',
		3027 => '1',
		3028 => '1',
		3029 => '1',
		3030 => '1',
		3031 => '1',
		3032 => '1',
		3033 => '0',
		3034 => '0',
		3035 => '0',
		3036 => '0',
		3037 => '0',
		3038 => '0',
		3039 => '0',
		3040 => '0',
		3041 => '0',
		3042 => '0',
		3043 => '0',
		3044 => '0',
		3045 => '0',
		3046 => '0',
		3047 => '0',
		3048 => '0',
		3049 => '0',
		3050 => '0',
		3051 => '0',
		3052 => '0',
		3053 => '0',
		3054 => '0',
		3055 => '0',
		3056 => '0',
		3057 => '0',
		3058 => '0',
		3059 => '0',
		3060 => '0',
		3061 => '0',
		3062 => '0',
		3063 => '0',
		3072 => '0',
		3073 => '0',
		3074 => '0',
		3075 => '0',
		3076 => '0',
		3077 => '0',
		3078 => '0',
		3079 => '0',
		3080 => '0',
		3081 => '0',
		3082 => '0',
		3083 => '0',
		3084 => '0',
		3085 => '0',
		3086 => '0',
		3087 => '0',
		3088 => '0',
		3089 => '0',
		3090 => '0',
		3091 => '0',
		3092 => '0',
		3093 => '0',
		3094 => '0',
		3095 => '0',
		3096 => '0',
		3097 => '0',
		3098 => '0',
		3099 => '0',
		3100 => '0',
		3101 => '0',
		3102 => '1',
		3103 => '1',
		3104 => '1',
		3105 => '1',
		3106 => '1',
		3107 => '1',
		3108 => '1',
		3109 => '1',
		3110 => '1',
		3111 => '1',
		3112 => '1',
		3113 => '1',
		3114 => '0',
		3115 => '0',
		3116 => '0',
		3117 => '0',
		3118 => '0',
		3119 => '1',
		3120 => '1',
		3121 => '1',
		3122 => '1',
		3123 => '1',
		3124 => '1',
		3125 => '1',
		3126 => '1',
		3127 => '1',
		3128 => '0',
		3129 => '0',
		3130 => '0',
		3131 => '0',
		3132 => '0',
		3133 => '0',
		3134 => '0',
		3135 => '0',
		3136 => '0',
		3137 => '0',
		3138 => '0',
		3139 => '0',
		3140 => '1',
		3141 => '1',
		3142 => '1',
		3143 => '1',
		3144 => '1',
		3145 => '1',
		3146 => '1',
		3147 => '0',
		3148 => '0',
		3149 => '0',
		3150 => '1',
		3151 => '1',
		3152 => '1',
		3153 => '1',
		3154 => '1',
		3155 => '1',
		3156 => '1',
		3157 => '1',
		3158 => '1',
		3159 => '1',
		3160 => '1',
		3161 => '1',
		3162 => '0',
		3163 => '0',
		3164 => '0',
		3165 => '0',
		3166 => '0',
		3167 => '0',
		3168 => '0',
		3169 => '0',
		3170 => '0',
		3171 => '0',
		3172 => '0',
		3173 => '0',
		3174 => '0',
		3175 => '0',
		3176 => '0',
		3177 => '0',
		3178 => '0',
		3179 => '0',
		3180 => '0',
		3181 => '0',
		3182 => '0',
		3183 => '0',
		3184 => '0',
		3185 => '0',
		3186 => '0',
		3187 => '0',
		3188 => '0',
		3189 => '0',
		3190 => '0',
		3191 => '0',
		3200 => '0',
		3201 => '0',
		3202 => '0',
		3203 => '0',
		3204 => '0',
		3205 => '0',
		3206 => '0',
		3207 => '0',
		3208 => '0',
		3209 => '0',
		3210 => '0',
		3211 => '0',
		3212 => '0',
		3213 => '0',
		3214 => '0',
		3215 => '0',
		3216 => '0',
		3217 => '0',
		3218 => '0',
		3219 => '0',
		3220 => '0',
		3221 => '0',
		3222 => '0',
		3223 => '0',
		3224 => '0',
		3225 => '0',
		3226 => '0',
		3227 => '0',
		3228 => '0',
		3229 => '1',
		3230 => '1',
		3231 => '1',
		3232 => '1',
		3233 => '1',
		3234 => '1',
		3235 => '1',
		3236 => '1',
		3237 => '1',
		3238 => '1',
		3239 => '1',
		3240 => '0',
		3241 => '0',
		3242 => '0',
		3243 => '0',
		3244 => '0',
		3245 => '1',
		3246 => '1',
		3247 => '1',
		3248 => '1',
		3249 => '1',
		3250 => '1',
		3251 => '0',
		3252 => '0',
		3253 => '0',
		3254 => '0',
		3255 => '0',
		3256 => '0',
		3257 => '0',
		3258 => '0',
		3259 => '0',
		3260 => '0',
		3261 => '0',
		3262 => '0',
		3263 => '0',
		3264 => '0',
		3265 => '0',
		3266 => '0',
		3267 => '0',
		3268 => '0',
		3269 => '0',
		3270 => '0',
		3271 => '0',
		3272 => '0',
		3273 => '1',
		3274 => '1',
		3275 => '1',
		3276 => '1',
		3277 => '0',
		3278 => '0',
		3279 => '0',
		3280 => '1',
		3281 => '1',
		3282 => '1',
		3283 => '1',
		3284 => '1',
		3285 => '1',
		3286 => '1',
		3287 => '1',
		3288 => '1',
		3289 => '1',
		3290 => '1',
		3291 => '0',
		3292 => '0',
		3293 => '0',
		3294 => '0',
		3295 => '0',
		3296 => '0',
		3297 => '0',
		3298 => '0',
		3299 => '0',
		3300 => '0',
		3301 => '0',
		3302 => '0',
		3303 => '0',
		3304 => '0',
		3305 => '0',
		3306 => '0',
		3307 => '0',
		3308 => '0',
		3309 => '0',
		3310 => '0',
		3311 => '0',
		3312 => '0',
		3313 => '0',
		3314 => '0',
		3315 => '0',
		3316 => '0',
		3317 => '0',
		3318 => '0',
		3319 => '0',
		3328 => '0',
		3329 => '0',
		3330 => '0',
		3331 => '0',
		3332 => '0',
		3333 => '0',
		3334 => '0',
		3335 => '0',
		3336 => '0',
		3337 => '0',
		3338 => '0',
		3339 => '0',
		3340 => '0',
		3341 => '0',
		3342 => '0',
		3343 => '0',
		3344 => '0',
		3345 => '0',
		3346 => '0',
		3347 => '0',
		3348 => '0',
		3349 => '0',
		3350 => '0',
		3351 => '0',
		3352 => '0',
		3353 => '0',
		3354 => '0',
		3355 => '0',
		3356 => '1',
		3357 => '1',
		3358 => '1',
		3359 => '1',
		3360 => '1',
		3361 => '1',
		3362 => '1',
		3363 => '1',
		3364 => '1',
		3365 => '1',
		3366 => '0',
		3367 => '0',
		3368 => '0',
		3369 => '0',
		3370 => '0',
		3371 => '1',
		3372 => '1',
		3373 => '1',
		3374 => '1',
		3375 => '1',
		3376 => '0',
		3377 => '0',
		3378 => '0',
		3379 => '0',
		3380 => '0',
		3381 => '0',
		3382 => '0',
		3383 => '0',
		3384 => '0',
		3385 => '1',
		3386 => '1',
		3387 => '1',
		3388 => '1',
		3389 => '1',
		3390 => '1',
		3391 => '1',
		3392 => '1',
		3393 => '1',
		3394 => '1',
		3395 => '1',
		3396 => '1',
		3397 => '0',
		3398 => '0',
		3399 => '0',
		3400 => '0',
		3401 => '0',
		3402 => '0',
		3403 => '0',
		3404 => '1',
		3405 => '1',
		3406 => '1',
		3407 => '0',
		3408 => '0',
		3409 => '0',
		3410 => '1',
		3411 => '1',
		3412 => '1',
		3413 => '1',
		3414 => '1',
		3415 => '1',
		3416 => '1',
		3417 => '1',
		3418 => '1',
		3419 => '1',
		3420 => '0',
		3421 => '0',
		3422 => '0',
		3423 => '0',
		3424 => '0',
		3425 => '0',
		3426 => '0',
		3427 => '0',
		3428 => '0',
		3429 => '0',
		3430 => '0',
		3431 => '0',
		3432 => '0',
		3433 => '0',
		3434 => '0',
		3435 => '0',
		3436 => '0',
		3437 => '0',
		3438 => '0',
		3439 => '0',
		3440 => '0',
		3441 => '0',
		3442 => '0',
		3443 => '0',
		3444 => '0',
		3445 => '0',
		3446 => '0',
		3447 => '0',
		3456 => '0',
		3457 => '0',
		3458 => '0',
		3459 => '0',
		3460 => '0',
		3461 => '0',
		3462 => '0',
		3463 => '0',
		3464 => '0',
		3465 => '0',
		3466 => '0',
		3467 => '0',
		3468 => '0',
		3469 => '0',
		3470 => '0',
		3471 => '0',
		3472 => '0',
		3473 => '0',
		3474 => '0',
		3475 => '0',
		3476 => '0',
		3477 => '0',
		3478 => '0',
		3479 => '0',
		3480 => '0',
		3481 => '0',
		3482 => '0',
		3483 => '1',
		3484 => '1',
		3485 => '1',
		3486 => '1',
		3487 => '1',
		3488 => '1',
		3489 => '1',
		3490 => '1',
		3491 => '1',
		3492 => '1',
		3493 => '0',
		3494 => '0',
		3495 => '0',
		3496 => '0',
		3497 => '1',
		3498 => '1',
		3499 => '1',
		3500 => '1',
		3501 => '1',
		3502 => '0',
		3503 => '0',
		3504 => '0',
		3505 => '0',
		3506 => '0',
		3507 => '0',
		3508 => '1',
		3509 => '1',
		3510 => '1',
		3511 => '1',
		3512 => '1',
		3513 => '1',
		3514 => '0',
		3515 => '0',
		3516 => '0',
		3517 => '0',
		3518 => '0',
		3519 => '0',
		3520 => '0',
		3521 => '0',
		3522 => '0',
		3523 => '0',
		3524 => '0',
		3525 => '0',
		3526 => '1',
		3527 => '1',
		3528 => '1',
		3529 => '1',
		3530 => '0',
		3531 => '0',
		3532 => '0',
		3533 => '0',
		3534 => '1',
		3535 => '1',
		3536 => '1',
		3537 => '0',
		3538 => '0',
		3539 => '1',
		3540 => '1',
		3541 => '1',
		3542 => '1',
		3543 => '1',
		3544 => '1',
		3545 => '1',
		3546 => '1',
		3547 => '1',
		3548 => '1',
		3549 => '0',
		3550 => '0',
		3551 => '0',
		3552 => '0',
		3553 => '0',
		3554 => '0',
		3555 => '0',
		3556 => '0',
		3557 => '0',
		3558 => '0',
		3559 => '0',
		3560 => '0',
		3561 => '0',
		3562 => '0',
		3563 => '0',
		3564 => '0',
		3565 => '0',
		3566 => '0',
		3567 => '0',
		3568 => '0',
		3569 => '0',
		3570 => '0',
		3571 => '0',
		3572 => '0',
		3573 => '0',
		3574 => '0',
		3575 => '0',
		3584 => '0',
		3585 => '0',
		3586 => '0',
		3587 => '0',
		3588 => '0',
		3589 => '0',
		3590 => '0',
		3591 => '0',
		3592 => '0',
		3593 => '0',
		3594 => '0',
		3595 => '0',
		3596 => '0',
		3597 => '0',
		3598 => '0',
		3599 => '0',
		3600 => '0',
		3601 => '0',
		3602 => '0',
		3603 => '0',
		3604 => '0',
		3605 => '0',
		3606 => '0',
		3607 => '0',
		3608 => '0',
		3609 => '0',
		3610 => '1',
		3611 => '1',
		3612 => '1',
		3613 => '1',
		3614 => '1',
		3615 => '1',
		3616 => '1',
		3617 => '1',
		3618 => '1',
		3619 => '0',
		3620 => '0',
		3621 => '0',
		3622 => '0',
		3623 => '1',
		3624 => '1',
		3625 => '1',
		3626 => '1',
		3627 => '1',
		3628 => '0',
		3629 => '0',
		3630 => '0',
		3631 => '0',
		3632 => '0',
		3633 => '1',
		3634 => '1',
		3635 => '1',
		3636 => '1',
		3637 => '0',
		3638 => '0',
		3639 => '0',
		3640 => '0',
		3641 => '0',
		3642 => '0',
		3643 => '0',
		3644 => '0',
		3645 => '0',
		3646 => '0',
		3647 => '0',
		3648 => '0',
		3649 => '0',
		3650 => '0',
		3651 => '0',
		3652 => '0',
		3653 => '0',
		3654 => '0',
		3655 => '0',
		3656 => '0',
		3657 => '0',
		3658 => '0',
		3659 => '1',
		3660 => '1',
		3661 => '0',
		3662 => '0',
		3663 => '0',
		3664 => '1',
		3665 => '1',
		3666 => '1',
		3667 => '0',
		3668 => '0',
		3669 => '1',
		3670 => '1',
		3671 => '1',
		3672 => '1',
		3673 => '1',
		3674 => '1',
		3675 => '1',
		3676 => '1',
		3677 => '1',
		3678 => '0',
		3679 => '0',
		3680 => '0',
		3681 => '0',
		3682 => '0',
		3683 => '0',
		3684 => '0',
		3685 => '0',
		3686 => '0',
		3687 => '0',
		3688 => '0',
		3689 => '0',
		3690 => '0',
		3691 => '0',
		3692 => '0',
		3693 => '0',
		3694 => '0',
		3695 => '0',
		3696 => '0',
		3697 => '0',
		3698 => '0',
		3699 => '0',
		3700 => '0',
		3701 => '0',
		3702 => '0',
		3703 => '0',
		3712 => '0',
		3713 => '0',
		3714 => '0',
		3715 => '0',
		3716 => '0',
		3717 => '0',
		3718 => '0',
		3719 => '0',
		3720 => '0',
		3721 => '0',
		3722 => '0',
		3723 => '0',
		3724 => '0',
		3725 => '0',
		3726 => '0',
		3727 => '0',
		3728 => '0',
		3729 => '0',
		3730 => '0',
		3731 => '0',
		3732 => '0',
		3733 => '0',
		3734 => '0',
		3735 => '0',
		3736 => '0',
		3737 => '1',
		3738 => '1',
		3739 => '1',
		3740 => '1',
		3741 => '1',
		3742 => '1',
		3743 => '1',
		3744 => '1',
		3745 => '1',
		3746 => '0',
		3747 => '0',
		3748 => '0',
		3749 => '0',
		3750 => '1',
		3751 => '1',
		3752 => '1',
		3753 => '1',
		3754 => '0',
		3755 => '0',
		3756 => '0',
		3757 => '0',
		3758 => '0',
		3759 => '1',
		3760 => '1',
		3761 => '1',
		3762 => '0',
		3763 => '0',
		3764 => '0',
		3765 => '0',
		3766 => '0',
		3767 => '0',
		3768 => '0',
		3769 => '0',
		3770 => '0',
		3771 => '0',
		3772 => '0',
		3773 => '0',
		3774 => '0',
		3775 => '0',
		3776 => '0',
		3777 => '0',
		3778 => '0',
		3779 => '0',
		3780 => '0',
		3781 => '0',
		3782 => '0',
		3783 => '0',
		3784 => '0',
		3785 => '0',
		3786 => '0',
		3787 => '0',
		3788 => '0',
		3789 => '0',
		3790 => '1',
		3791 => '0',
		3792 => '0',
		3793 => '0',
		3794 => '1',
		3795 => '1',
		3796 => '0',
		3797 => '0',
		3798 => '1',
		3799 => '1',
		3800 => '1',
		3801 => '1',
		3802 => '1',
		3803 => '1',
		3804 => '1',
		3805 => '1',
		3806 => '1',
		3807 => '0',
		3808 => '0',
		3809 => '0',
		3810 => '0',
		3811 => '0',
		3812 => '0',
		3813 => '0',
		3814 => '0',
		3815 => '0',
		3816 => '0',
		3817 => '0',
		3818 => '0',
		3819 => '0',
		3820 => '0',
		3821 => '0',
		3822 => '0',
		3823 => '0',
		3824 => '0',
		3825 => '0',
		3826 => '0',
		3827 => '0',
		3828 => '0',
		3829 => '0',
		3830 => '0',
		3831 => '0',
		3840 => '0',
		3841 => '0',
		3842 => '0',
		3843 => '0',
		3844 => '0',
		3845 => '0',
		3846 => '0',
		3847 => '0',
		3848 => '0',
		3849 => '0',
		3850 => '0',
		3851 => '0',
		3852 => '0',
		3853 => '0',
		3854 => '0',
		3855 => '0',
		3856 => '0',
		3857 => '0',
		3858 => '0',
		3859 => '0',
		3860 => '0',
		3861 => '0',
		3862 => '0',
		3863 => '0',
		3864 => '1',
		3865 => '1',
		3866 => '1',
		3867 => '1',
		3868 => '1',
		3869 => '1',
		3870 => '1',
		3871 => '1',
		3872 => '1',
		3873 => '0',
		3874 => '0',
		3875 => '0',
		3876 => '1',
		3877 => '1',
		3878 => '1',
		3879 => '1',
		3880 => '0',
		3881 => '0',
		3882 => '0',
		3883 => '0',
		3884 => '0',
		3885 => '1',
		3886 => '1',
		3887 => '1',
		3888 => '0',
		3889 => '0',
		3890 => '0',
		3891 => '0',
		3892 => '0',
		3893 => '0',
		3894 => '0',
		3895 => '0',
		3896 => '0',
		3897 => '0',
		3898 => '0',
		3899 => '0',
		3900 => '0',
		3901 => '0',
		3902 => '0',
		3903 => '0',
		3904 => '0',
		3905 => '0',
		3906 => '0',
		3907 => '0',
		3908 => '0',
		3909 => '0',
		3910 => '0',
		3911 => '0',
		3912 => '0',
		3913 => '0',
		3914 => '0',
		3915 => '0',
		3916 => '0',
		3917 => '0',
		3918 => '0',
		3919 => '0',
		3920 => '1',
		3921 => '0',
		3922 => '0',
		3923 => '0',
		3924 => '1',
		3925 => '1',
		3926 => '0',
		3927 => '1',
		3928 => '1',
		3929 => '1',
		3930 => '1',
		3931 => '1',
		3932 => '1',
		3933 => '1',
		3934 => '1',
		3935 => '1',
		3936 => '0',
		3937 => '0',
		3938 => '0',
		3939 => '0',
		3940 => '0',
		3941 => '0',
		3942 => '0',
		3943 => '0',
		3944 => '0',
		3945 => '0',
		3946 => '0',
		3947 => '0',
		3948 => '0',
		3949 => '0',
		3950 => '0',
		3951 => '0',
		3952 => '0',
		3953 => '0',
		3954 => '0',
		3955 => '0',
		3956 => '0',
		3957 => '0',
		3958 => '0',
		3959 => '0',
		3968 => '0',
		3969 => '0',
		3970 => '0',
		3971 => '0',
		3972 => '0',
		3973 => '0',
		3974 => '0',
		3975 => '0',
		3976 => '0',
		3977 => '0',
		3978 => '0',
		3979 => '0',
		3980 => '0',
		3981 => '0',
		3982 => '0',
		3983 => '0',
		3984 => '0',
		3985 => '0',
		3986 => '0',
		3987 => '0',
		3988 => '0',
		3989 => '0',
		3990 => '0',
		3991 => '1',
		3992 => '1',
		3993 => '1',
		3994 => '1',
		3995 => '1',
		3996 => '1',
		3997 => '1',
		3998 => '1',
		3999 => '1',
		4000 => '0',
		4001 => '0',
		4002 => '0',
		4003 => '1',
		4004 => '1',
		4005 => '1',
		4006 => '1',
		4007 => '0',
		4008 => '0',
		4009 => '0',
		4010 => '0',
		4011 => '1',
		4012 => '1',
		4013 => '1',
		4014 => '0',
		4015 => '0',
		4016 => '0',
		4017 => '0',
		4018 => '0',
		4019 => '0',
		4020 => '0',
		4021 => '0',
		4022 => '0',
		4023 => '0',
		4024 => '0',
		4025 => '0',
		4026 => '0',
		4027 => '0',
		4028 => '0',
		4029 => '0',
		4030 => '0',
		4031 => '0',
		4032 => '0',
		4033 => '0',
		4034 => '0',
		4035 => '0',
		4036 => '0',
		4037 => '0',
		4038 => '0',
		4039 => '0',
		4040 => '0',
		4041 => '0',
		4042 => '0',
		4043 => '0',
		4044 => '0',
		4045 => '0',
		4046 => '0',
		4047 => '0',
		4048 => '0',
		4049 => '0',
		4050 => '1',
		4051 => '0',
		4052 => '0',
		4053 => '1',
		4054 => '1',
		4055 => '0',
		4056 => '1',
		4057 => '1',
		4058 => '1',
		4059 => '1',
		4060 => '1',
		4061 => '1',
		4062 => '1',
		4063 => '1',
		4064 => '1',
		4065 => '0',
		4066 => '0',
		4067 => '0',
		4068 => '0',
		4069 => '0',
		4070 => '0',
		4071 => '0',
		4072 => '0',
		4073 => '0',
		4074 => '0',
		4075 => '0',
		4076 => '0',
		4077 => '0',
		4078 => '0',
		4079 => '0',
		4080 => '0',
		4081 => '0',
		4082 => '0',
		4083 => '0',
		4084 => '0',
		4085 => '0',
		4086 => '0',
		4087 => '0',
		4096 => '0',
		4097 => '0',
		4098 => '0',
		4099 => '0',
		4100 => '0',
		4101 => '0',
		4102 => '0',
		4103 => '0',
		4104 => '0',
		4105 => '0',
		4106 => '0',
		4107 => '0',
		4108 => '0',
		4109 => '0',
		4110 => '0',
		4111 => '0',
		4112 => '0',
		4113 => '0',
		4114 => '0',
		4115 => '0',
		4116 => '0',
		4117 => '0',
		4118 => '0',
		4119 => '1',
		4120 => '1',
		4121 => '1',
		4122 => '1',
		4123 => '1',
		4124 => '1',
		4125 => '1',
		4126 => '1',
		4127 => '0',
		4128 => '0',
		4129 => '0',
		4130 => '1',
		4131 => '1',
		4132 => '1',
		4133 => '0',
		4134 => '0',
		4135 => '0',
		4136 => '0',
		4137 => '1',
		4138 => '1',
		4139 => '1',
		4140 => '0',
		4141 => '0',
		4142 => '0',
		4143 => '0',
		4144 => '0',
		4145 => '0',
		4146 => '0',
		4147 => '0',
		4148 => '0',
		4149 => '0',
		4150 => '0',
		4151 => '0',
		4152 => '0',
		4153 => '0',
		4154 => '0',
		4155 => '0',
		4156 => '0',
		4157 => '0',
		4158 => '0',
		4159 => '0',
		4160 => '0',
		4161 => '0',
		4162 => '0',
		4163 => '0',
		4164 => '0',
		4165 => '0',
		4166 => '0',
		4167 => '0',
		4168 => '0',
		4169 => '0',
		4170 => '0',
		4171 => '0',
		4172 => '0',
		4173 => '0',
		4174 => '0',
		4175 => '0',
		4176 => '0',
		4177 => '0',
		4178 => '0',
		4179 => '0',
		4180 => '1',
		4181 => '0',
		4182 => '0',
		4183 => '1',
		4184 => '0',
		4185 => '1',
		4186 => '1',
		4187 => '1',
		4188 => '1',
		4189 => '1',
		4190 => '1',
		4191 => '1',
		4192 => '1',
		4193 => '1',
		4194 => '0',
		4195 => '0',
		4196 => '0',
		4197 => '0',
		4198 => '0',
		4199 => '0',
		4200 => '0',
		4201 => '0',
		4202 => '0',
		4203 => '0',
		4204 => '0',
		4205 => '0',
		4206 => '0',
		4207 => '0',
		4208 => '0',
		4209 => '0',
		4210 => '0',
		4211 => '0',
		4212 => '0',
		4213 => '0',
		4214 => '0',
		4215 => '0',
		4224 => '0',
		4225 => '0',
		4226 => '0',
		4227 => '0',
		4228 => '0',
		4229 => '0',
		4230 => '0',
		4231 => '0',
		4232 => '0',
		4233 => '0',
		4234 => '0',
		4235 => '0',
		4236 => '0',
		4237 => '0',
		4238 => '0',
		4239 => '0',
		4240 => '0',
		4241 => '0',
		4242 => '0',
		4243 => '0',
		4244 => '0',
		4245 => '0',
		4246 => '1',
		4247 => '1',
		4248 => '1',
		4249 => '1',
		4250 => '1',
		4251 => '1',
		4252 => '1',
		4253 => '1',
		4254 => '0',
		4255 => '0',
		4256 => '0',
		4257 => '1',
		4258 => '1',
		4259 => '1',
		4260 => '0',
		4261 => '0',
		4262 => '0',
		4263 => '0',
		4264 => '1',
		4265 => '1',
		4266 => '0',
		4267 => '0',
		4268 => '0',
		4269 => '0',
		4270 => '0',
		4271 => '0',
		4272 => '0',
		4273 => '0',
		4274 => '0',
		4275 => '0',
		4276 => '0',
		4277 => '0',
		4278 => '0',
		4279 => '0',
		4280 => '0',
		4281 => '0',
		4282 => '0',
		4283 => '0',
		4284 => '0',
		4285 => '0',
		4286 => '0',
		4287 => '0',
		4288 => '0',
		4289 => '0',
		4290 => '0',
		4291 => '0',
		4292 => '0',
		4293 => '0',
		4294 => '0',
		4295 => '0',
		4296 => '0',
		4297 => '0',
		4298 => '0',
		4299 => '0',
		4300 => '0',
		4301 => '0',
		4302 => '0',
		4303 => '0',
		4304 => '0',
		4305 => '0',
		4306 => '0',
		4307 => '0',
		4308 => '0',
		4309 => '0',
		4310 => '0',
		4311 => '0',
		4312 => '1',
		4313 => '0',
		4314 => '1',
		4315 => '1',
		4316 => '1',
		4317 => '1',
		4318 => '1',
		4319 => '1',
		4320 => '1',
		4321 => '1',
		4322 => '0',
		4323 => '0',
		4324 => '0',
		4325 => '0',
		4326 => '0',
		4327 => '0',
		4328 => '0',
		4329 => '0',
		4330 => '0',
		4331 => '0',
		4332 => '0',
		4333 => '0',
		4334 => '0',
		4335 => '0',
		4336 => '0',
		4337 => '0',
		4338 => '0',
		4339 => '0',
		4340 => '0',
		4341 => '0',
		4342 => '0',
		4343 => '0',
		4352 => '0',
		4353 => '0',
		4354 => '0',
		4355 => '0',
		4356 => '0',
		4357 => '0',
		4358 => '0',
		4359 => '0',
		4360 => '0',
		4361 => '0',
		4362 => '0',
		4363 => '0',
		4364 => '0',
		4365 => '0',
		4366 => '0',
		4367 => '0',
		4368 => '0',
		4369 => '0',
		4370 => '0',
		4371 => '0',
		4372 => '0',
		4373 => '1',
		4374 => '1',
		4375 => '1',
		4376 => '1',
		4377 => '1',
		4378 => '1',
		4379 => '1',
		4380 => '1',
		4381 => '0',
		4382 => '0',
		4383 => '0',
		4384 => '1',
		4385 => '1',
		4386 => '1',
		4387 => '0',
		4388 => '0',
		4389 => '0',
		4390 => '1',
		4391 => '1',
		4392 => '1',
		4393 => '0',
		4394 => '0',
		4395 => '0',
		4396 => '0',
		4397 => '0',
		4398 => '0',
		4399 => '0',
		4400 => '0',
		4401 => '0',
		4402 => '0',
		4403 => '0',
		4404 => '0',
		4405 => '0',
		4406 => '0',
		4407 => '0',
		4408 => '0',
		4409 => '0',
		4410 => '0',
		4411 => '0',
		4412 => '0',
		4413 => '0',
		4414 => '0',
		4415 => '0',
		4416 => '0',
		4417 => '0',
		4418 => '0',
		4419 => '0',
		4420 => '0',
		4421 => '0',
		4422 => '0',
		4423 => '0',
		4424 => '0',
		4425 => '0',
		4426 => '0',
		4427 => '0',
		4428 => '0',
		4429 => '0',
		4430 => '0',
		4431 => '0',
		4432 => '0',
		4433 => '0',
		4434 => '0',
		4435 => '0',
		4436 => '0',
		4437 => '0',
		4438 => '0',
		4439 => '1',
		4440 => '0',
		4441 => '1',
		4442 => '0',
		4443 => '1',
		4444 => '1',
		4445 => '1',
		4446 => '1',
		4447 => '1',
		4448 => '1',
		4449 => '1',
		4450 => '1',
		4451 => '0',
		4452 => '0',
		4453 => '0',
		4454 => '0',
		4455 => '0',
		4456 => '0',
		4457 => '0',
		4458 => '0',
		4459 => '0',
		4460 => '0',
		4461 => '0',
		4462 => '0',
		4463 => '0',
		4464 => '0',
		4465 => '0',
		4466 => '0',
		4467 => '0',
		4468 => '0',
		4469 => '0',
		4470 => '0',
		4471 => '0',
		4480 => '0',
		4481 => '0',
		4482 => '0',
		4483 => '0',
		4484 => '0',
		4485 => '0',
		4486 => '0',
		4487 => '0',
		4488 => '0',
		4489 => '0',
		4490 => '0',
		4491 => '0',
		4492 => '0',
		4493 => '0',
		4494 => '0',
		4495 => '0',
		4496 => '0',
		4497 => '0',
		4498 => '0',
		4499 => '0',
		4500 => '0',
		4501 => '1',
		4502 => '1',
		4503 => '1',
		4504 => '1',
		4505 => '1',
		4506 => '1',
		4507 => '1',
		4508 => '0',
		4509 => '0',
		4510 => '0',
		4511 => '1',
		4512 => '1',
		4513 => '1',
		4514 => '0',
		4515 => '0',
		4516 => '0',
		4517 => '1',
		4518 => '1',
		4519 => '0',
		4520 => '0',
		4521 => '0',
		4522 => '0',
		4523 => '0',
		4524 => '0',
		4525 => '0',
		4526 => '0',
		4527 => '0',
		4528 => '0',
		4529 => '0',
		4530 => '0',
		4531 => '0',
		4532 => '0',
		4533 => '0',
		4534 => '0',
		4535 => '0',
		4536 => '0',
		4537 => '0',
		4538 => '0',
		4539 => '0',
		4540 => '0',
		4541 => '0',
		4542 => '0',
		4543 => '0',
		4544 => '0',
		4545 => '0',
		4546 => '0',
		4547 => '0',
		4548 => '0',
		4549 => '0',
		4550 => '0',
		4551 => '0',
		4552 => '0',
		4553 => '0',
		4554 => '0',
		4555 => '0',
		4556 => '0',
		4557 => '0',
		4558 => '0',
		4559 => '0',
		4560 => '0',
		4561 => '0',
		4562 => '0',
		4563 => '0',
		4564 => '0',
		4565 => '0',
		4566 => '0',
		4567 => '0',
		4568 => '0',
		4569 => '0',
		4570 => '1',
		4571 => '0',
		4572 => '1',
		4573 => '1',
		4574 => '1',
		4575 => '1',
		4576 => '1',
		4577 => '1',
		4578 => '1',
		4579 => '1',
		4580 => '0',
		4581 => '0',
		4582 => '0',
		4583 => '0',
		4584 => '0',
		4585 => '0',
		4586 => '0',
		4587 => '0',
		4588 => '0',
		4589 => '0',
		4590 => '0',
		4591 => '0',
		4592 => '0',
		4593 => '0',
		4594 => '0',
		4595 => '0',
		4596 => '0',
		4597 => '0',
		4598 => '0',
		4599 => '0',
		4608 => '0',
		4609 => '0',
		4610 => '0',
		4611 => '0',
		4612 => '0',
		4613 => '0',
		4614 => '0',
		4615 => '0',
		4616 => '0',
		4617 => '0',
		4618 => '0',
		4619 => '0',
		4620 => '0',
		4621 => '0',
		4622 => '0',
		4623 => '0',
		4624 => '0',
		4625 => '0',
		4626 => '0',
		4627 => '0',
		4628 => '1',
		4629 => '1',
		4630 => '1',
		4631 => '1',
		4632 => '1',
		4633 => '1',
		4634 => '1',
		4635 => '1',
		4636 => '0',
		4637 => '0',
		4638 => '1',
		4639 => '1',
		4640 => '1',
		4641 => '0',
		4642 => '0',
		4643 => '0',
		4644 => '1',
		4645 => '1',
		4646 => '0',
		4647 => '0',
		4648 => '0',
		4649 => '0',
		4650 => '0',
		4651 => '0',
		4652 => '0',
		4653 => '0',
		4654 => '0',
		4655 => '0',
		4656 => '0',
		4657 => '0',
		4658 => '0',
		4659 => '0',
		4660 => '0',
		4661 => '0',
		4662 => '0',
		4663 => '0',
		4664 => '0',
		4665 => '0',
		4666 => '0',
		4667 => '0',
		4668 => '0',
		4669 => '0',
		4670 => '0',
		4671 => '0',
		4672 => '0',
		4673 => '0',
		4674 => '0',
		4675 => '0',
		4676 => '0',
		4677 => '0',
		4678 => '0',
		4679 => '0',
		4680 => '0',
		4681 => '0',
		4682 => '0',
		4683 => '0',
		4684 => '0',
		4685 => '0',
		4686 => '0',
		4687 => '0',
		4688 => '0',
		4689 => '0',
		4690 => '0',
		4691 => '0',
		4692 => '0',
		4693 => '0',
		4694 => '0',
		4695 => '0',
		4696 => '0',
		4697 => '0',
		4698 => '0',
		4699 => '1',
		4700 => '1',
		4701 => '1',
		4702 => '1',
		4703 => '1',
		4704 => '1',
		4705 => '1',
		4706 => '1',
		4707 => '1',
		4708 => '0',
		4709 => '0',
		4710 => '0',
		4711 => '0',
		4712 => '0',
		4713 => '0',
		4714 => '0',
		4715 => '0',
		4716 => '0',
		4717 => '0',
		4718 => '0',
		4719 => '0',
		4720 => '0',
		4721 => '0',
		4722 => '0',
		4723 => '0',
		4724 => '0',
		4725 => '0',
		4726 => '0',
		4727 => '0',
		4736 => '0',
		4737 => '0',
		4738 => '0',
		4739 => '0',
		4740 => '0',
		4741 => '0',
		4742 => '0',
		4743 => '0',
		4744 => '0',
		4745 => '0',
		4746 => '0',
		4747 => '0',
		4748 => '0',
		4749 => '0',
		4750 => '0',
		4751 => '0',
		4752 => '0',
		4753 => '0',
		4754 => '0',
		4755 => '0',
		4756 => '1',
		4757 => '1',
		4758 => '1',
		4759 => '1',
		4760 => '1',
		4761 => '1',
		4762 => '1',
		4763 => '0',
		4764 => '0',
		4765 => '1',
		4766 => '1',
		4767 => '1',
		4768 => '0',
		4769 => '0',
		4770 => '0',
		4771 => '1',
		4772 => '1',
		4773 => '0',
		4774 => '0',
		4775 => '0',
		4776 => '0',
		4777 => '0',
		4778 => '0',
		4779 => '0',
		4780 => '0',
		4781 => '0',
		4782 => '0',
		4783 => '0',
		4784 => '0',
		4785 => '0',
		4786 => '0',
		4787 => '0',
		4788 => '0',
		4789 => '0',
		4790 => '0',
		4791 => '0',
		4792 => '0',
		4793 => '0',
		4794 => '0',
		4795 => '0',
		4796 => '0',
		4797 => '0',
		4798 => '0',
		4799 => '0',
		4800 => '0',
		4801 => '0',
		4802 => '0',
		4803 => '0',
		4804 => '0',
		4805 => '0',
		4806 => '0',
		4807 => '0',
		4808 => '0',
		4809 => '0',
		4810 => '0',
		4811 => '0',
		4812 => '0',
		4813 => '0',
		4814 => '0',
		4815 => '0',
		4816 => '0',
		4817 => '0',
		4818 => '0',
		4819 => '0',
		4820 => '0',
		4821 => '0',
		4822 => '0',
		4823 => '0',
		4824 => '0',
		4825 => '0',
		4826 => '0',
		4827 => '0',
		4828 => '0',
		4829 => '1',
		4830 => '1',
		4831 => '1',
		4832 => '1',
		4833 => '1',
		4834 => '1',
		4835 => '1',
		4836 => '1',
		4837 => '0',
		4838 => '0',
		4839 => '0',
		4840 => '0',
		4841 => '0',
		4842 => '0',
		4843 => '0',
		4844 => '0',
		4845 => '0',
		4846 => '0',
		4847 => '0',
		4848 => '0',
		4849 => '0',
		4850 => '0',
		4851 => '0',
		4852 => '0',
		4853 => '0',
		4854 => '0',
		4855 => '0',
		4864 => '0',
		4865 => '0',
		4866 => '0',
		4867 => '0',
		4868 => '0',
		4869 => '0',
		4870 => '0',
		4871 => '0',
		4872 => '0',
		4873 => '0',
		4874 => '0',
		4875 => '0',
		4876 => '0',
		4877 => '0',
		4878 => '0',
		4879 => '0',
		4880 => '0',
		4881 => '0',
		4882 => '0',
		4883 => '1',
		4884 => '1',
		4885 => '1',
		4886 => '1',
		4887 => '1',
		4888 => '1',
		4889 => '1',
		4890 => '0',
		4891 => '0',
		4892 => '0',
		4893 => '1',
		4894 => '1',
		4895 => '0',
		4896 => '0',
		4897 => '0',
		4898 => '1',
		4899 => '1',
		4900 => '0',
		4901 => '0',
		4902 => '0',
		4903 => '0',
		4904 => '0',
		4905 => '0',
		4906 => '0',
		4907 => '0',
		4908 => '0',
		4909 => '0',
		4910 => '0',
		4911 => '0',
		4912 => '0',
		4913 => '0',
		4914 => '0',
		4915 => '0',
		4916 => '0',
		4917 => '0',
		4918 => '0',
		4919 => '0',
		4920 => '0',
		4921 => '0',
		4922 => '0',
		4923 => '0',
		4924 => '0',
		4925 => '0',
		4926 => '0',
		4927 => '0',
		4928 => '0',
		4929 => '0',
		4930 => '0',
		4931 => '0',
		4932 => '0',
		4933 => '0',
		4934 => '0',
		4935 => '0',
		4936 => '0',
		4937 => '0',
		4938 => '0',
		4939 => '0',
		4940 => '0',
		4941 => '0',
		4942 => '0',
		4943 => '0',
		4944 => '0',
		4945 => '0',
		4946 => '0',
		4947 => '0',
		4948 => '0',
		4949 => '0',
		4950 => '0',
		4951 => '0',
		4952 => '0',
		4953 => '0',
		4954 => '0',
		4955 => '0',
		4956 => '1',
		4957 => '0',
		4958 => '1',
		4959 => '1',
		4960 => '1',
		4961 => '1',
		4962 => '1',
		4963 => '1',
		4964 => '1',
		4965 => '0',
		4966 => '0',
		4967 => '0',
		4968 => '0',
		4969 => '0',
		4970 => '0',
		4971 => '0',
		4972 => '0',
		4973 => '0',
		4974 => '0',
		4975 => '0',
		4976 => '0',
		4977 => '0',
		4978 => '0',
		4979 => '0',
		4980 => '0',
		4981 => '0',
		4982 => '0',
		4983 => '0',
		4992 => '0',
		4993 => '0',
		4994 => '0',
		4995 => '0',
		4996 => '0',
		4997 => '0',
		4998 => '0',
		4999 => '0',
		5000 => '0',
		5001 => '0',
		5002 => '0',
		5003 => '0',
		5004 => '0',
		5005 => '0',
		5006 => '0',
		5007 => '0',
		5008 => '0',
		5009 => '0',
		5010 => '0',
		5011 => '1',
		5012 => '1',
		5013 => '1',
		5014 => '1',
		5015 => '1',
		5016 => '1',
		5017 => '1',
		5018 => '0',
		5019 => '0',
		5020 => '1',
		5021 => '1',
		5022 => '0',
		5023 => '0',
		5024 => '0',
		5025 => '1',
		5026 => '1',
		5027 => '0',
		5028 => '0',
		5029 => '0',
		5030 => '0',
		5031 => '0',
		5032 => '0',
		5033 => '0',
		5034 => '0',
		5035 => '0',
		5036 => '0',
		5037 => '0',
		5038 => '0',
		5039 => '0',
		5040 => '0',
		5041 => '0',
		5042 => '0',
		5043 => '0',
		5044 => '0',
		5045 => '0',
		5046 => '0',
		5047 => '0',
		5048 => '0',
		5049 => '0',
		5050 => '0',
		5051 => '0',
		5052 => '0',
		5053 => '0',
		5054 => '0',
		5055 => '0',
		5056 => '0',
		5057 => '0',
		5058 => '0',
		5059 => '0',
		5060 => '0',
		5061 => '0',
		5062 => '0',
		5063 => '0',
		5064 => '0',
		5065 => '0',
		5066 => '0',
		5067 => '0',
		5068 => '0',
		5069 => '0',
		5070 => '0',
		5071 => '0',
		5072 => '0',
		5073 => '0',
		5074 => '0',
		5075 => '0',
		5076 => '0',
		5077 => '0',
		5078 => '0',
		5079 => '0',
		5080 => '0',
		5081 => '0',
		5082 => '0',
		5083 => '0',
		5084 => '0',
		5085 => '1',
		5086 => '1',
		5087 => '1',
		5088 => '1',
		5089 => '1',
		5090 => '1',
		5091 => '1',
		5092 => '1',
		5093 => '1',
		5094 => '0',
		5095 => '0',
		5096 => '0',
		5097 => '0',
		5098 => '0',
		5099 => '0',
		5100 => '0',
		5101 => '0',
		5102 => '0',
		5103 => '0',
		5104 => '0',
		5105 => '0',
		5106 => '0',
		5107 => '0',
		5108 => '0',
		5109 => '0',
		5110 => '0',
		5111 => '0',
		5120 => '0',
		5121 => '0',
		5122 => '0',
		5123 => '0',
		5124 => '0',
		5125 => '0',
		5126 => '0',
		5127 => '0',
		5128 => '0',
		5129 => '0',
		5130 => '0',
		5131 => '0',
		5132 => '0',
		5133 => '0',
		5134 => '0',
		5135 => '0',
		5136 => '0',
		5137 => '0',
		5138 => '1',
		5139 => '1',
		5140 => '1',
		5141 => '1',
		5142 => '1',
		5143 => '1',
		5144 => '1',
		5145 => '0',
		5146 => '0',
		5147 => '1',
		5148 => '1',
		5149 => '1',
		5150 => '0',
		5151 => '0',
		5152 => '1',
		5153 => '1',
		5154 => '0',
		5155 => '0',
		5156 => '0',
		5157 => '0',
		5158 => '0',
		5159 => '0',
		5160 => '0',
		5161 => '0',
		5162 => '0',
		5163 => '0',
		5164 => '0',
		5165 => '0',
		5166 => '0',
		5167 => '0',
		5168 => '0',
		5169 => '0',
		5170 => '0',
		5171 => '0',
		5172 => '0',
		5173 => '0',
		5174 => '0',
		5175 => '0',
		5176 => '0',
		5177 => '0',
		5178 => '0',
		5179 => '0',
		5180 => '0',
		5181 => '0',
		5182 => '0',
		5183 => '0',
		5184 => '0',
		5185 => '0',
		5186 => '0',
		5187 => '0',
		5188 => '0',
		5189 => '0',
		5190 => '0',
		5191 => '0',
		5192 => '0',
		5193 => '0',
		5194 => '0',
		5195 => '0',
		5196 => '0',
		5197 => '0',
		5198 => '0',
		5199 => '0',
		5200 => '0',
		5201 => '0',
		5202 => '0',
		5203 => '0',
		5204 => '0',
		5205 => '0',
		5206 => '0',
		5207 => '0',
		5208 => '0',
		5209 => '0',
		5210 => '0',
		5211 => '0',
		5212 => '0',
		5213 => '0',
		5214 => '0',
		5215 => '1',
		5216 => '1',
		5217 => '1',
		5218 => '1',
		5219 => '1',
		5220 => '1',
		5221 => '1',
		5222 => '0',
		5223 => '0',
		5224 => '0',
		5225 => '0',
		5226 => '0',
		5227 => '0',
		5228 => '0',
		5229 => '0',
		5230 => '0',
		5231 => '0',
		5232 => '0',
		5233 => '0',
		5234 => '0',
		5235 => '0',
		5236 => '0',
		5237 => '0',
		5238 => '0',
		5239 => '0',
		5248 => '0',
		5249 => '0',
		5250 => '0',
		5251 => '0',
		5252 => '0',
		5253 => '0',
		5254 => '0',
		5255 => '0',
		5256 => '0',
		5257 => '0',
		5258 => '0',
		5259 => '0',
		5260 => '0',
		5261 => '0',
		5262 => '0',
		5263 => '0',
		5264 => '0',
		5265 => '0',
		5266 => '1',
		5267 => '1',
		5268 => '1',
		5269 => '1',
		5270 => '1',
		5271 => '1',
		5272 => '1',
		5273 => '0',
		5274 => '0',
		5275 => '1',
		5276 => '1',
		5277 => '0',
		5278 => '0',
		5279 => '1',
		5280 => '1',
		5281 => '0',
		5282 => '0',
		5283 => '0',
		5284 => '0',
		5285 => '0',
		5286 => '0',
		5287 => '0',
		5288 => '0',
		5289 => '0',
		5290 => '0',
		5291 => '0',
		5292 => '0',
		5293 => '0',
		5294 => '0',
		5295 => '0',
		5296 => '0',
		5297 => '0',
		5298 => '0',
		5299 => '0',
		5300 => '0',
		5301 => '0',
		5302 => '0',
		5303 => '0',
		5304 => '0',
		5305 => '0',
		5306 => '0',
		5307 => '0',
		5308 => '0',
		5309 => '0',
		5310 => '0',
		5311 => '0',
		5312 => '0',
		5313 => '0',
		5314 => '0',
		5315 => '0',
		5316 => '0',
		5317 => '0',
		5318 => '0',
		5319 => '0',
		5320 => '0',
		5321 => '0',
		5322 => '0',
		5323 => '0',
		5324 => '0',
		5325 => '0',
		5326 => '0',
		5327 => '0',
		5328 => '0',
		5329 => '0',
		5330 => '0',
		5331 => '0',
		5332 => '0',
		5333 => '0',
		5334 => '0',
		5335 => '0',
		5336 => '0',
		5337 => '0',
		5338 => '0',
		5339 => '0',
		5340 => '0',
		5341 => '0',
		5342 => '1',
		5343 => '1',
		5344 => '1',
		5345 => '1',
		5346 => '1',
		5347 => '1',
		5348 => '1',
		5349 => '1',
		5350 => '1',
		5351 => '0',
		5352 => '0',
		5353 => '0',
		5354 => '0',
		5355 => '0',
		5356 => '0',
		5357 => '0',
		5358 => '0',
		5359 => '0',
		5360 => '0',
		5361 => '0',
		5362 => '0',
		5363 => '0',
		5364 => '0',
		5365 => '0',
		5366 => '0',
		5367 => '0',
		5376 => '0',
		5377 => '0',
		5378 => '0',
		5379 => '0',
		5380 => '0',
		5381 => '0',
		5382 => '0',
		5383 => '0',
		5384 => '0',
		5385 => '0',
		5386 => '0',
		5387 => '0',
		5388 => '0',
		5389 => '0',
		5390 => '0',
		5391 => '0',
		5392 => '0',
		5393 => '1',
		5394 => '1',
		5395 => '1',
		5396 => '1',
		5397 => '1',
		5398 => '1',
		5399 => '1',
		5400 => '0',
		5401 => '0',
		5402 => '1',
		5403 => '1',
		5404 => '0',
		5405 => '0',
		5406 => '0',
		5407 => '1',
		5408 => '0',
		5409 => '0',
		5410 => '0',
		5411 => '0',
		5412 => '0',
		5413 => '0',
		5414 => '0',
		5415 => '0',
		5416 => '0',
		5417 => '0',
		5418 => '0',
		5419 => '0',
		5420 => '0',
		5421 => '0',
		5422 => '0',
		5423 => '0',
		5424 => '0',
		5425 => '0',
		5426 => '0',
		5427 => '0',
		5428 => '0',
		5429 => '0',
		5430 => '0',
		5431 => '0',
		5432 => '0',
		5433 => '0',
		5434 => '0',
		5435 => '0',
		5436 => '0',
		5437 => '0',
		5438 => '0',
		5439 => '0',
		5440 => '0',
		5441 => '0',
		5442 => '0',
		5443 => '0',
		5444 => '0',
		5445 => '0',
		5446 => '0',
		5447 => '0',
		5448 => '0',
		5449 => '0',
		5450 => '0',
		5451 => '0',
		5452 => '0',
		5453 => '0',
		5454 => '0',
		5455 => '0',
		5456 => '0',
		5457 => '0',
		5458 => '0',
		5459 => '0',
		5460 => '0',
		5461 => '0',
		5462 => '0',
		5463 => '0',
		5464 => '0',
		5465 => '0',
		5466 => '0',
		5467 => '0',
		5468 => '0',
		5469 => '0',
		5470 => '0',
		5471 => '0',
		5472 => '1',
		5473 => '1',
		5474 => '1',
		5475 => '1',
		5476 => '1',
		5477 => '1',
		5478 => '1',
		5479 => '0',
		5480 => '0',
		5481 => '0',
		5482 => '0',
		5483 => '0',
		5484 => '0',
		5485 => '0',
		5486 => '0',
		5487 => '0',
		5488 => '0',
		5489 => '0',
		5490 => '0',
		5491 => '0',
		5492 => '0',
		5493 => '0',
		5494 => '0',
		5495 => '0',
		5504 => '0',
		5505 => '0',
		5506 => '0',
		5507 => '0',
		5508 => '0',
		5509 => '0',
		5510 => '0',
		5511 => '0',
		5512 => '0',
		5513 => '0',
		5514 => '0',
		5515 => '0',
		5516 => '0',
		5517 => '0',
		5518 => '0',
		5519 => '0',
		5520 => '0',
		5521 => '1',
		5522 => '1',
		5523 => '1',
		5524 => '1',
		5525 => '1',
		5526 => '1',
		5527 => '1',
		5528 => '0',
		5529 => '0',
		5530 => '1',
		5531 => '1',
		5532 => '0',
		5533 => '0',
		5534 => '1',
		5535 => '1',
		5536 => '0',
		5537 => '0',
		5538 => '0',
		5539 => '0',
		5540 => '0',
		5541 => '0',
		5542 => '0',
		5543 => '0',
		5544 => '0',
		5545 => '0',
		5546 => '0',
		5547 => '0',
		5548 => '0',
		5549 => '0',
		5550 => '0',
		5551 => '0',
		5552 => '0',
		5553 => '0',
		5554 => '0',
		5555 => '0',
		5556 => '0',
		5557 => '0',
		5558 => '0',
		5559 => '0',
		5560 => '0',
		5561 => '0',
		5562 => '0',
		5563 => '0',
		5564 => '0',
		5565 => '0',
		5566 => '0',
		5567 => '0',
		5568 => '0',
		5569 => '0',
		5570 => '0',
		5571 => '0',
		5572 => '0',
		5573 => '0',
		5574 => '0',
		5575 => '0',
		5576 => '0',
		5577 => '0',
		5578 => '0',
		5579 => '0',
		5580 => '0',
		5581 => '0',
		5582 => '0',
		5583 => '0',
		5584 => '0',
		5585 => '0',
		5586 => '0',
		5587 => '0',
		5588 => '0',
		5589 => '0',
		5590 => '0',
		5591 => '0',
		5592 => '0',
		5593 => '0',
		5594 => '0',
		5595 => '0',
		5596 => '0',
		5597 => '0',
		5598 => '0',
		5599 => '1',
		5600 => '1',
		5601 => '1',
		5602 => '1',
		5603 => '1',
		5604 => '1',
		5605 => '1',
		5606 => '1',
		5607 => '1',
		5608 => '0',
		5609 => '0',
		5610 => '0',
		5611 => '0',
		5612 => '0',
		5613 => '0',
		5614 => '0',
		5615 => '0',
		5616 => '0',
		5617 => '0',
		5618 => '0',
		5619 => '0',
		5620 => '0',
		5621 => '0',
		5622 => '0',
		5623 => '0',
		5632 => '0',
		5633 => '0',
		5634 => '0',
		5635 => '0',
		5636 => '0',
		5637 => '0',
		5638 => '0',
		5639 => '0',
		5640 => '0',
		5641 => '0',
		5642 => '0',
		5643 => '0',
		5644 => '0',
		5645 => '0',
		5646 => '0',
		5647 => '0',
		5648 => '1',
		5649 => '1',
		5650 => '1',
		5651 => '1',
		5652 => '1',
		5653 => '1',
		5654 => '1',
		5655 => '0',
		5656 => '0',
		5657 => '1',
		5658 => '1',
		5659 => '0',
		5660 => '0',
		5661 => '1',
		5662 => '1',
		5663 => '0',
		5664 => '0',
		5665 => '0',
		5666 => '0',
		5667 => '0',
		5668 => '0',
		5669 => '0',
		5670 => '0',
		5671 => '0',
		5672 => '0',
		5673 => '0',
		5674 => '0',
		5675 => '0',
		5676 => '0',
		5677 => '0',
		5678 => '0',
		5679 => '0',
		5680 => '0',
		5681 => '0',
		5682 => '0',
		5683 => '0',
		5684 => '0',
		5685 => '0',
		5686 => '0',
		5687 => '0',
		5688 => '0',
		5689 => '0',
		5690 => '0',
		5691 => '0',
		5692 => '0',
		5693 => '0',
		5694 => '0',
		5695 => '0',
		5696 => '0',
		5697 => '0',
		5698 => '0',
		5699 => '0',
		5700 => '0',
		5701 => '0',
		5702 => '0',
		5703 => '0',
		5704 => '0',
		5705 => '0',
		5706 => '0',
		5707 => '0',
		5708 => '0',
		5709 => '0',
		5710 => '0',
		5711 => '0',
		5712 => '0',
		5713 => '0',
		5714 => '0',
		5715 => '0',
		5716 => '0',
		5717 => '0',
		5718 => '0',
		5719 => '0',
		5720 => '0',
		5721 => '0',
		5722 => '0',
		5723 => '0',
		5724 => '0',
		5725 => '0',
		5726 => '0',
		5727 => '0',
		5728 => '0',
		5729 => '1',
		5730 => '1',
		5731 => '1',
		5732 => '1',
		5733 => '1',
		5734 => '1',
		5735 => '1',
		5736 => '0',
		5737 => '0',
		5738 => '0',
		5739 => '0',
		5740 => '0',
		5741 => '0',
		5742 => '0',
		5743 => '0',
		5744 => '0',
		5745 => '0',
		5746 => '0',
		5747 => '0',
		5748 => '0',
		5749 => '0',
		5750 => '0',
		5751 => '0',
		5760 => '0',
		5761 => '0',
		5762 => '0',
		5763 => '0',
		5764 => '0',
		5765 => '0',
		5766 => '0',
		5767 => '0',
		5768 => '0',
		5769 => '0',
		5770 => '0',
		5771 => '0',
		5772 => '0',
		5773 => '0',
		5774 => '0',
		5775 => '0',
		5776 => '1',
		5777 => '1',
		5778 => '1',
		5779 => '1',
		5780 => '1',
		5781 => '1',
		5782 => '1',
		5783 => '0',
		5784 => '0',
		5785 => '1',
		5786 => '1',
		5787 => '0',
		5788 => '0',
		5789 => '1',
		5790 => '0',
		5791 => '0',
		5792 => '0',
		5793 => '0',
		5794 => '0',
		5795 => '0',
		5796 => '0',
		5797 => '0',
		5798 => '0',
		5799 => '0',
		5800 => '0',
		5801 => '0',
		5802 => '0',
		5803 => '0',
		5804 => '0',
		5805 => '0',
		5806 => '0',
		5807 => '0',
		5808 => '0',
		5809 => '0',
		5810 => '0',
		5811 => '0',
		5812 => '0',
		5813 => '0',
		5814 => '0',
		5815 => '0',
		5816 => '0',
		5817 => '0',
		5818 => '0',
		5819 => '0',
		5820 => '0',
		5821 => '0',
		5822 => '0',
		5823 => '0',
		5824 => '0',
		5825 => '0',
		5826 => '0',
		5827 => '0',
		5828 => '0',
		5829 => '0',
		5830 => '0',
		5831 => '0',
		5832 => '0',
		5833 => '0',
		5834 => '0',
		5835 => '0',
		5836 => '0',
		5837 => '0',
		5838 => '0',
		5839 => '0',
		5840 => '0',
		5841 => '0',
		5842 => '0',
		5843 => '0',
		5844 => '0',
		5845 => '0',
		5846 => '0',
		5847 => '0',
		5848 => '0',
		5849 => '0',
		5850 => '0',
		5851 => '0',
		5852 => '0',
		5853 => '0',
		5854 => '0',
		5855 => '0',
		5856 => '1',
		5857 => '1',
		5858 => '1',
		5859 => '1',
		5860 => '1',
		5861 => '1',
		5862 => '1',
		5863 => '1',
		5864 => '1',
		5865 => '0',
		5866 => '0',
		5867 => '0',
		5868 => '0',
		5869 => '0',
		5870 => '0',
		5871 => '0',
		5872 => '0',
		5873 => '0',
		5874 => '0',
		5875 => '0',
		5876 => '0',
		5877 => '0',
		5878 => '0',
		5879 => '0',
		5888 => '0',
		5889 => '0',
		5890 => '0',
		5891 => '0',
		5892 => '0',
		5893 => '0',
		5894 => '0',
		5895 => '0',
		5896 => '0',
		5897 => '0',
		5898 => '0',
		5899 => '0',
		5900 => '0',
		5901 => '0',
		5902 => '0',
		5903 => '0',
		5904 => '1',
		5905 => '1',
		5906 => '1',
		5907 => '1',
		5908 => '1',
		5909 => '1',
		5910 => '0',
		5911 => '0',
		5912 => '1',
		5913 => '1',
		5914 => '0',
		5915 => '0',
		5916 => '1',
		5917 => '1',
		5918 => '0',
		5919 => '0',
		5920 => '0',
		5921 => '0',
		5922 => '0',
		5923 => '0',
		5924 => '0',
		5925 => '0',
		5926 => '0',
		5927 => '0',
		5928 => '0',
		5929 => '0',
		5930 => '0',
		5931 => '0',
		5932 => '0',
		5933 => '0',
		5934 => '0',
		5935 => '0',
		5936 => '0',
		5937 => '0',
		5938 => '0',
		5939 => '0',
		5940 => '0',
		5941 => '0',
		5942 => '0',
		5943 => '0',
		5944 => '0',
		5945 => '0',
		5946 => '0',
		5947 => '0',
		5948 => '0',
		5949 => '0',
		5950 => '0',
		5951 => '0',
		5952 => '0',
		5953 => '0',
		5954 => '0',
		5955 => '0',
		5956 => '0',
		5957 => '0',
		5958 => '0',
		5959 => '0',
		5960 => '0',
		5961 => '0',
		5962 => '0',
		5963 => '0',
		5964 => '0',
		5965 => '0',
		5966 => '0',
		5967 => '0',
		5968 => '0',
		5969 => '0',
		5970 => '0',
		5971 => '0',
		5972 => '0',
		5973 => '0',
		5974 => '0',
		5975 => '0',
		5976 => '0',
		5977 => '0',
		5978 => '0',
		5979 => '0',
		5980 => '0',
		5981 => '0',
		5982 => '0',
		5983 => '0',
		5984 => '0',
		5985 => '0',
		5986 => '1',
		5987 => '1',
		5988 => '1',
		5989 => '1',
		5990 => '1',
		5991 => '1',
		5992 => '0',
		5993 => '0',
		5994 => '0',
		5995 => '0',
		5996 => '0',
		5997 => '0',
		5998 => '0',
		5999 => '0',
		6000 => '0',
		6001 => '0',
		6002 => '0',
		6003 => '0',
		6004 => '0',
		6005 => '0',
		6006 => '0',
		6007 => '0',
		6016 => '0',
		6017 => '0',
		6018 => '0',
		6019 => '0',
		6020 => '0',
		6021 => '0',
		6022 => '0',
		6023 => '0',
		6024 => '0',
		6025 => '0',
		6026 => '0',
		6027 => '0',
		6028 => '0',
		6029 => '0',
		6030 => '0',
		6031 => '1',
		6032 => '1',
		6033 => '1',
		6034 => '1',
		6035 => '1',
		6036 => '1',
		6037 => '1',
		6038 => '0',
		6039 => '0',
		6040 => '1',
		6041 => '1',
		6042 => '0',
		6043 => '0',
		6044 => '1',
		6045 => '0',
		6046 => '0',
		6047 => '0',
		6048 => '0',
		6049 => '0',
		6050 => '0',
		6051 => '0',
		6052 => '0',
		6053 => '0',
		6054 => '0',
		6055 => '0',
		6056 => '0',
		6057 => '0',
		6058 => '0',
		6059 => '0',
		6060 => '0',
		6061 => '0',
		6062 => '0',
		6063 => '0',
		6064 => '0',
		6065 => '0',
		6066 => '0',
		6067 => '0',
		6068 => '0',
		6069 => '0',
		6070 => '0',
		6071 => '0',
		6072 => '0',
		6073 => '0',
		6074 => '0',
		6075 => '0',
		6076 => '0',
		6077 => '0',
		6078 => '0',
		6079 => '0',
		6080 => '0',
		6081 => '0',
		6082 => '0',
		6083 => '0',
		6084 => '0',
		6085 => '0',
		6086 => '0',
		6087 => '0',
		6088 => '0',
		6089 => '0',
		6090 => '0',
		6091 => '0',
		6092 => '0',
		6093 => '0',
		6094 => '0',
		6095 => '0',
		6096 => '0',
		6097 => '0',
		6098 => '0',
		6099 => '0',
		6100 => '0',
		6101 => '0',
		6102 => '0',
		6103 => '0',
		6104 => '0',
		6105 => '0',
		6106 => '0',
		6107 => '0',
		6108 => '0',
		6109 => '0',
		6110 => '0',
		6111 => '0',
		6112 => '0',
		6113 => '1',
		6114 => '1',
		6115 => '1',
		6116 => '1',
		6117 => '1',
		6118 => '1',
		6119 => '1',
		6120 => '1',
		6121 => '1',
		6122 => '0',
		6123 => '0',
		6124 => '0',
		6125 => '0',
		6126 => '0',
		6127 => '0',
		6128 => '0',
		6129 => '0',
		6130 => '0',
		6131 => '0',
		6132 => '0',
		6133 => '0',
		6134 => '0',
		6135 => '0',
		6144 => '0',
		6145 => '0',
		6146 => '0',
		6147 => '0',
		6148 => '0',
		6149 => '0',
		6150 => '0',
		6151 => '0',
		6152 => '0',
		6153 => '0',
		6154 => '0',
		6155 => '0',
		6156 => '0',
		6157 => '0',
		6158 => '0',
		6159 => '1',
		6160 => '1',
		6161 => '1',
		6162 => '1',
		6163 => '1',
		6164 => '1',
		6165 => '1',
		6166 => '0',
		6167 => '1',
		6168 => '1',
		6169 => '0',
		6170 => '0',
		6171 => '1',
		6172 => '1',
		6173 => '0',
		6174 => '0',
		6175 => '0',
		6176 => '0',
		6177 => '0',
		6178 => '0',
		6179 => '0',
		6180 => '0',
		6181 => '0',
		6182 => '0',
		6183 => '0',
		6184 => '0',
		6185 => '0',
		6186 => '0',
		6187 => '0',
		6188 => '0',
		6189 => '0',
		6190 => '0',
		6191 => '0',
		6192 => '0',
		6193 => '0',
		6194 => '0',
		6195 => '0',
		6196 => '0',
		6197 => '0',
		6198 => '0',
		6199 => '0',
		6200 => '0',
		6201 => '0',
		6202 => '0',
		6203 => '0',
		6204 => '0',
		6205 => '0',
		6206 => '0',
		6207 => '0',
		6208 => '0',
		6209 => '0',
		6210 => '0',
		6211 => '0',
		6212 => '0',
		6213 => '0',
		6214 => '0',
		6215 => '0',
		6216 => '0',
		6217 => '0',
		6218 => '0',
		6219 => '0',
		6220 => '0',
		6221 => '0',
		6222 => '0',
		6223 => '0',
		6224 => '0',
		6225 => '0',
		6226 => '0',
		6227 => '0',
		6228 => '0',
		6229 => '0',
		6230 => '0',
		6231 => '0',
		6232 => '0',
		6233 => '0',
		6234 => '0',
		6235 => '0',
		6236 => '0',
		6237 => '0',
		6238 => '0',
		6239 => '0',
		6240 => '0',
		6241 => '0',
		6242 => '1',
		6243 => '1',
		6244 => '1',
		6245 => '1',
		6246 => '1',
		6247 => '1',
		6248 => '1',
		6249 => '1',
		6250 => '0',
		6251 => '0',
		6252 => '0',
		6253 => '0',
		6254 => '0',
		6255 => '0',
		6256 => '0',
		6257 => '0',
		6258 => '0',
		6259 => '0',
		6260 => '0',
		6261 => '0',
		6262 => '0',
		6263 => '0',
		6272 => '0',
		6273 => '0',
		6274 => '0',
		6275 => '0',
		6276 => '0',
		6277 => '0',
		6278 => '0',
		6279 => '0',
		6280 => '0',
		6281 => '0',
		6282 => '0',
		6283 => '0',
		6284 => '0',
		6285 => '0',
		6286 => '0',
		6287 => '1',
		6288 => '1',
		6289 => '1',
		6290 => '1',
		6291 => '1',
		6292 => '1',
		6293 => '0',
		6294 => '0',
		6295 => '1',
		6296 => '1',
		6297 => '0',
		6298 => '0',
		6299 => '1',
		6300 => '0',
		6301 => '0',
		6302 => '0',
		6303 => '0',
		6304 => '0',
		6305 => '0',
		6306 => '0',
		6307 => '0',
		6308 => '0',
		6309 => '0',
		6310 => '0',
		6311 => '0',
		6312 => '0',
		6313 => '0',
		6314 => '0',
		6315 => '0',
		6316 => '0',
		6317 => '0',
		6318 => '0',
		6319 => '0',
		6320 => '0',
		6321 => '0',
		6322 => '0',
		6323 => '0',
		6324 => '0',
		6325 => '0',
		6326 => '0',
		6327 => '0',
		6328 => '0',
		6329 => '0',
		6330 => '0',
		6331 => '0',
		6332 => '0',
		6333 => '0',
		6334 => '0',
		6335 => '0',
		6336 => '0',
		6337 => '0',
		6338 => '0',
		6339 => '0',
		6340 => '0',
		6341 => '0',
		6342 => '0',
		6343 => '0',
		6344 => '0',
		6345 => '0',
		6346 => '0',
		6347 => '0',
		6348 => '0',
		6349 => '0',
		6350 => '0',
		6351 => '0',
		6352 => '0',
		6353 => '0',
		6354 => '0',
		6355 => '0',
		6356 => '0',
		6357 => '0',
		6358 => '0',
		6359 => '0',
		6360 => '0',
		6361 => '0',
		6362 => '0',
		6363 => '0',
		6364 => '0',
		6365 => '0',
		6366 => '0',
		6367 => '0',
		6368 => '0',
		6369 => '0',
		6370 => '0',
		6371 => '1',
		6372 => '1',
		6373 => '1',
		6374 => '1',
		6375 => '1',
		6376 => '1',
		6377 => '0',
		6378 => '1',
		6379 => '0',
		6380 => '0',
		6381 => '0',
		6382 => '0',
		6383 => '0',
		6384 => '0',
		6385 => '0',
		6386 => '0',
		6387 => '0',
		6388 => '0',
		6389 => '0',
		6390 => '0',
		6391 => '0',
		6400 => '0',
		6401 => '0',
		6402 => '0',
		6403 => '0',
		6404 => '0',
		6405 => '0',
		6406 => '0',
		6407 => '0',
		6408 => '0',
		6409 => '0',
		6410 => '0',
		6411 => '0',
		6412 => '0',
		6413 => '0',
		6414 => '0',
		6415 => '1',
		6416 => '1',
		6417 => '1',
		6418 => '1',
		6419 => '1',
		6420 => '1',
		6421 => '0',
		6422 => '0',
		6423 => '1',
		6424 => '0',
		6425 => '0',
		6426 => '1',
		6427 => '1',
		6428 => '0',
		6429 => '0',
		6430 => '0',
		6431 => '0',
		6432 => '0',
		6433 => '0',
		6434 => '0',
		6435 => '0',
		6436 => '0',
		6437 => '0',
		6438 => '0',
		6439 => '0',
		6440 => '0',
		6441 => '0',
		6442 => '0',
		6443 => '0',
		6444 => '0',
		6445 => '0',
		6446 => '0',
		6447 => '0',
		6448 => '0',
		6449 => '0',
		6450 => '0',
		6451 => '0',
		6452 => '0',
		6453 => '0',
		6454 => '0',
		6455 => '0',
		6456 => '0',
		6457 => '0',
		6458 => '0',
		6459 => '0',
		6460 => '0',
		6461 => '0',
		6462 => '0',
		6463 => '0',
		6464 => '0',
		6465 => '0',
		6466 => '0',
		6467 => '0',
		6468 => '0',
		6469 => '0',
		6470 => '0',
		6471 => '0',
		6472 => '0',
		6473 => '0',
		6474 => '0',
		6475 => '0',
		6476 => '0',
		6477 => '0',
		6478 => '0',
		6479 => '0',
		6480 => '0',
		6481 => '0',
		6482 => '0',
		6483 => '0',
		6484 => '0',
		6485 => '0',
		6486 => '0',
		6487 => '0',
		6488 => '0',
		6489 => '0',
		6490 => '0',
		6491 => '0',
		6492 => '0',
		6493 => '0',
		6494 => '0',
		6495 => '0',
		6496 => '0',
		6497 => '0',
		6498 => '1',
		6499 => '1',
		6500 => '1',
		6501 => '1',
		6502 => '1',
		6503 => '1',
		6504 => '1',
		6505 => '0',
		6506 => '0',
		6507 => '0',
		6508 => '0',
		6509 => '0',
		6510 => '0',
		6511 => '0',
		6512 => '0',
		6513 => '0',
		6514 => '0',
		6515 => '0',
		6516 => '0',
		6517 => '0',
		6518 => '0',
		6519 => '0',
		6528 => '0',
		6529 => '0',
		6530 => '0',
		6531 => '0',
		6532 => '0',
		6533 => '0',
		6534 => '0',
		6535 => '0',
		6536 => '0',
		6537 => '0',
		6538 => '0',
		6539 => '0',
		6540 => '0',
		6541 => '0',
		6542 => '0',
		6543 => '1',
		6544 => '1',
		6545 => '1',
		6546 => '1',
		6547 => '1',
		6548 => '1',
		6549 => '0',
		6550 => '1',
		6551 => '1',
		6552 => '0',
		6553 => '0',
		6554 => '1',
		6555 => '0',
		6556 => '0',
		6557 => '0',
		6558 => '0',
		6559 => '0',
		6560 => '0',
		6561 => '0',
		6562 => '0',
		6563 => '0',
		6564 => '0',
		6565 => '0',
		6566 => '0',
		6567 => '0',
		6568 => '0',
		6569 => '0',
		6570 => '0',
		6571 => '0',
		6572 => '0',
		6573 => '0',
		6574 => '0',
		6575 => '0',
		6576 => '0',
		6577 => '0',
		6578 => '0',
		6579 => '0',
		6580 => '0',
		6581 => '0',
		6582 => '0',
		6583 => '0',
		6584 => '0',
		6585 => '0',
		6586 => '0',
		6587 => '0',
		6588 => '0',
		6589 => '0',
		6590 => '0',
		6591 => '0',
		6592 => '0',
		6593 => '0',
		6594 => '0',
		6595 => '0',
		6596 => '0',
		6597 => '0',
		6598 => '0',
		6599 => '0',
		6600 => '0',
		6601 => '0',
		6602 => '0',
		6603 => '0',
		6604 => '0',
		6605 => '0',
		6606 => '0',
		6607 => '0',
		6608 => '0',
		6609 => '0',
		6610 => '0',
		6611 => '0',
		6612 => '0',
		6613 => '0',
		6614 => '0',
		6615 => '0',
		6616 => '0',
		6617 => '0',
		6618 => '0',
		6619 => '0',
		6620 => '0',
		6621 => '0',
		6622 => '0',
		6623 => '0',
		6624 => '0',
		6625 => '0',
		6626 => '0',
		6627 => '1',
		6628 => '1',
		6629 => '1',
		6630 => '1',
		6631 => '1',
		6632 => '1',
		6633 => '0',
		6634 => '1',
		6635 => '1',
		6636 => '0',
		6637 => '0',
		6638 => '0',
		6639 => '0',
		6640 => '0',
		6641 => '0',
		6642 => '0',
		6643 => '0',
		6644 => '0',
		6645 => '0',
		6646 => '0',
		6647 => '0',
		6656 => '0',
		6657 => '0',
		6658 => '0',
		6659 => '0',
		6660 => '0',
		6661 => '0',
		6662 => '0',
		6663 => '0',
		6664 => '0',
		6665 => '0',
		6666 => '0',
		6667 => '0',
		6668 => '0',
		6669 => '0',
		6670 => '1',
		6671 => '1',
		6672 => '1',
		6673 => '1',
		6674 => '1',
		6675 => '1',
		6676 => '1',
		6677 => '0',
		6678 => '1',
		6679 => '1',
		6680 => '0',
		6681 => '1',
		6682 => '1',
		6683 => '0',
		6684 => '0',
		6685 => '0',
		6686 => '0',
		6687 => '0',
		6688 => '0',
		6689 => '0',
		6690 => '0',
		6691 => '0',
		6692 => '0',
		6693 => '0',
		6694 => '0',
		6695 => '0',
		6696 => '0',
		6697 => '0',
		6698 => '0',
		6699 => '0',
		6700 => '0',
		6701 => '0',
		6702 => '0',
		6703 => '0',
		6704 => '0',
		6705 => '0',
		6706 => '0',
		6707 => '0',
		6708 => '0',
		6709 => '0',
		6710 => '0',
		6711 => '0',
		6712 => '0',
		6713 => '0',
		6714 => '0',
		6715 => '0',
		6716 => '0',
		6717 => '0',
		6718 => '0',
		6719 => '0',
		6720 => '0',
		6721 => '0',
		6722 => '0',
		6723 => '0',
		6724 => '0',
		6725 => '0',
		6726 => '0',
		6727 => '0',
		6728 => '0',
		6729 => '0',
		6730 => '0',
		6731 => '0',
		6732 => '0',
		6733 => '0',
		6734 => '0',
		6735 => '0',
		6736 => '0',
		6737 => '0',
		6738 => '0',
		6739 => '0',
		6740 => '0',
		6741 => '0',
		6742 => '0',
		6743 => '0',
		6744 => '0',
		6745 => '0',
		6746 => '0',
		6747 => '0',
		6748 => '0',
		6749 => '0',
		6750 => '0',
		6751 => '0',
		6752 => '0',
		6753 => '0',
		6754 => '0',
		6755 => '1',
		6756 => '1',
		6757 => '1',
		6758 => '1',
		6759 => '1',
		6760 => '1',
		6761 => '1',
		6762 => '1',
		6763 => '1',
		6764 => '0',
		6765 => '0',
		6766 => '0',
		6767 => '0',
		6768 => '0',
		6769 => '0',
		6770 => '0',
		6771 => '0',
		6772 => '0',
		6773 => '0',
		6774 => '0',
		6775 => '0',
		6784 => '0',
		6785 => '0',
		6786 => '0',
		6787 => '0',
		6788 => '0',
		6789 => '0',
		6790 => '0',
		6791 => '0',
		6792 => '0',
		6793 => '0',
		6794 => '0',
		6795 => '0',
		6796 => '0',
		6797 => '0',
		6798 => '1',
		6799 => '1',
		6800 => '1',
		6801 => '1',
		6802 => '1',
		6803 => '1',
		6804 => '1',
		6805 => '0',
		6806 => '1',
		6807 => '0',
		6808 => '0',
		6809 => '1',
		6810 => '0',
		6811 => '0',
		6812 => '0',
		6813 => '0',
		6814 => '0',
		6815 => '0',
		6816 => '0',
		6817 => '0',
		6818 => '0',
		6819 => '0',
		6820 => '0',
		6821 => '0',
		6822 => '0',
		6823 => '0',
		6824 => '0',
		6825 => '0',
		6826 => '0',
		6827 => '0',
		6828 => '0',
		6829 => '0',
		6830 => '0',
		6831 => '0',
		6832 => '0',
		6833 => '0',
		6834 => '0',
		6835 => '0',
		6836 => '0',
		6837 => '0',
		6838 => '0',
		6839 => '0',
		6840 => '0',
		6841 => '0',
		6842 => '0',
		6843 => '0',
		6844 => '0',
		6845 => '0',
		6846 => '0',
		6847 => '0',
		6848 => '0',
		6849 => '0',
		6850 => '0',
		6851 => '0',
		6852 => '0',
		6853 => '0',
		6854 => '0',
		6855 => '0',
		6856 => '0',
		6857 => '0',
		6858 => '0',
		6859 => '0',
		6860 => '0',
		6861 => '0',
		6862 => '0',
		6863 => '0',
		6864 => '0',
		6865 => '0',
		6866 => '0',
		6867 => '0',
		6868 => '0',
		6869 => '0',
		6870 => '0',
		6871 => '0',
		6872 => '0',
		6873 => '0',
		6874 => '0',
		6875 => '0',
		6876 => '0',
		6877 => '0',
		6878 => '0',
		6879 => '0',
		6880 => '0',
		6881 => '0',
		6882 => '0',
		6883 => '1',
		6884 => '1',
		6885 => '1',
		6886 => '1',
		6887 => '1',
		6888 => '1',
		6889 => '1',
		6890 => '1',
		6891 => '0',
		6892 => '0',
		6893 => '0',
		6894 => '0',
		6895 => '0',
		6896 => '0',
		6897 => '0',
		6898 => '0',
		6899 => '0',
		6900 => '0',
		6901 => '0',
		6902 => '0',
		6903 => '0',
		6912 => '0',
		6913 => '0',
		6914 => '0',
		6915 => '0',
		6916 => '0',
		6917 => '0',
		6918 => '0',
		6919 => '0',
		6920 => '0',
		6921 => '0',
		6922 => '0',
		6923 => '0',
		6924 => '0',
		6925 => '0',
		6926 => '1',
		6927 => '1',
		6928 => '1',
		6929 => '1',
		6930 => '1',
		6931 => '1',
		6932 => '0',
		6933 => '0',
		6934 => '1',
		6935 => '0',
		6936 => '0',
		6937 => '1',
		6938 => '0',
		6939 => '0',
		6940 => '0',
		6941 => '0',
		6942 => '0',
		6943 => '0',
		6944 => '0',
		6945 => '0',
		6946 => '0',
		6947 => '0',
		6948 => '0',
		6949 => '0',
		6950 => '0',
		6951 => '0',
		6952 => '0',
		6953 => '0',
		6954 => '0',
		6955 => '0',
		6956 => '0',
		6957 => '0',
		6958 => '0',
		6959 => '0',
		6960 => '0',
		6961 => '0',
		6962 => '0',
		6963 => '0',
		6964 => '0',
		6965 => '0',
		6966 => '0',
		6967 => '0',
		6968 => '0',
		6969 => '0',
		6970 => '0',
		6971 => '0',
		6972 => '0',
		6973 => '0',
		6974 => '0',
		6975 => '0',
		6976 => '0',
		6977 => '0',
		6978 => '0',
		6979 => '0',
		6980 => '0',
		6981 => '0',
		6982 => '0',
		6983 => '0',
		6984 => '0',
		6985 => '0',
		6986 => '0',
		6987 => '0',
		6988 => '0',
		6989 => '0',
		6990 => '0',
		6991 => '0',
		6992 => '0',
		6993 => '0',
		6994 => '0',
		6995 => '0',
		6996 => '0',
		6997 => '0',
		6998 => '0',
		6999 => '0',
		7000 => '0',
		7001 => '0',
		7002 => '0',
		7003 => '0',
		7004 => '0',
		7005 => '0',
		7006 => '0',
		7007 => '0',
		7008 => '0',
		7009 => '0',
		7010 => '0',
		7011 => '0',
		7012 => '1',
		7013 => '1',
		7014 => '1',
		7015 => '1',
		7016 => '1',
		7017 => '1',
		7018 => '0',
		7019 => '0',
		7020 => '1',
		7021 => '0',
		7022 => '0',
		7023 => '0',
		7024 => '0',
		7025 => '0',
		7026 => '0',
		7027 => '0',
		7028 => '0',
		7029 => '0',
		7030 => '0',
		7031 => '0',
		7040 => '0',
		7041 => '0',
		7042 => '0',
		7043 => '0',
		7044 => '0',
		7045 => '0',
		7046 => '0',
		7047 => '0',
		7048 => '0',
		7049 => '0',
		7050 => '0',
		7051 => '0',
		7052 => '0',
		7053 => '0',
		7054 => '1',
		7055 => '1',
		7056 => '1',
		7057 => '1',
		7058 => '1',
		7059 => '1',
		7060 => '0',
		7061 => '0',
		7062 => '1',
		7063 => '0',
		7064 => '1',
		7065 => '1',
		7066 => '0',
		7067 => '0',
		7068 => '0',
		7069 => '0',
		7070 => '0',
		7071 => '0',
		7072 => '0',
		7073 => '0',
		7074 => '0',
		7075 => '0',
		7076 => '0',
		7077 => '0',
		7078 => '0',
		7079 => '0',
		7080 => '0',
		7081 => '0',
		7082 => '0',
		7083 => '0',
		7084 => '0',
		7085 => '0',
		7086 => '0',
		7087 => '0',
		7088 => '0',
		7089 => '0',
		7090 => '0',
		7091 => '0',
		7092 => '0',
		7093 => '0',
		7094 => '0',
		7095 => '0',
		7096 => '0',
		7097 => '0',
		7098 => '0',
		7099 => '0',
		7100 => '0',
		7101 => '0',
		7102 => '0',
		7103 => '0',
		7104 => '0',
		7105 => '0',
		7106 => '0',
		7107 => '0',
		7108 => '0',
		7109 => '0',
		7110 => '0',
		7111 => '0',
		7112 => '0',
		7113 => '0',
		7114 => '0',
		7115 => '0',
		7116 => '0',
		7117 => '0',
		7118 => '0',
		7119 => '0',
		7120 => '0',
		7121 => '0',
		7122 => '0',
		7123 => '0',
		7124 => '0',
		7125 => '0',
		7126 => '0',
		7127 => '0',
		7128 => '0',
		7129 => '0',
		7130 => '0',
		7131 => '0',
		7132 => '0',
		7133 => '0',
		7134 => '0',
		7135 => '0',
		7136 => '0',
		7137 => '0',
		7138 => '0',
		7139 => '1',
		7140 => '1',
		7141 => '1',
		7142 => '1',
		7143 => '1',
		7144 => '1',
		7145 => '1',
		7146 => '0',
		7147 => '0',
		7148 => '1',
		7149 => '0',
		7150 => '0',
		7151 => '0',
		7152 => '0',
		7153 => '0',
		7154 => '0',
		7155 => '0',
		7156 => '0',
		7157 => '0',
		7158 => '0',
		7159 => '0',
		7168 => '0',
		7169 => '0',
		7170 => '0',
		7171 => '0',
		7172 => '0',
		7173 => '0',
		7174 => '0',
		7175 => '0',
		7176 => '0',
		7177 => '0',
		7178 => '0',
		7179 => '0',
		7180 => '0',
		7181 => '0',
		7182 => '1',
		7183 => '1',
		7184 => '1',
		7185 => '1',
		7186 => '1',
		7187 => '1',
		7188 => '0',
		7189 => '1',
		7190 => '1',
		7191 => '0',
		7192 => '1',
		7193 => '0',
		7194 => '0',
		7195 => '0',
		7196 => '0',
		7197 => '0',
		7198 => '0',
		7199 => '0',
		7200 => '0',
		7201 => '0',
		7202 => '0',
		7203 => '0',
		7204 => '0',
		7205 => '0',
		7206 => '0',
		7207 => '0',
		7208 => '0',
		7209 => '0',
		7210 => '0',
		7211 => '0',
		7212 => '0',
		7213 => '0',
		7214 => '0',
		7215 => '0',
		7216 => '0',
		7217 => '0',
		7218 => '0',
		7219 => '0',
		7220 => '0',
		7221 => '0',
		7222 => '0',
		7223 => '0',
		7224 => '0',
		7225 => '0',
		7226 => '0',
		7227 => '0',
		7228 => '0',
		7229 => '0',
		7230 => '0',
		7231 => '0',
		7232 => '0',
		7233 => '0',
		7234 => '0',
		7235 => '0',
		7236 => '0',
		7237 => '0',
		7238 => '0',
		7239 => '0',
		7240 => '0',
		7241 => '0',
		7242 => '0',
		7243 => '0',
		7244 => '0',
		7245 => '0',
		7246 => '0',
		7247 => '0',
		7248 => '0',
		7249 => '0',
		7250 => '0',
		7251 => '0',
		7252 => '0',
		7253 => '0',
		7254 => '0',
		7255 => '0',
		7256 => '0',
		7257 => '0',
		7258 => '0',
		7259 => '0',
		7260 => '0',
		7261 => '0',
		7262 => '0',
		7263 => '0',
		7264 => '0',
		7265 => '0',
		7266 => '0',
		7267 => '0',
		7268 => '1',
		7269 => '1',
		7270 => '1',
		7271 => '1',
		7272 => '1',
		7273 => '1',
		7274 => '0',
		7275 => '1',
		7276 => '1',
		7277 => '0',
		7278 => '0',
		7279 => '0',
		7280 => '0',
		7281 => '0',
		7282 => '0',
		7283 => '0',
		7284 => '0',
		7285 => '0',
		7286 => '0',
		7287 => '0',
		7296 => '0',
		7297 => '0',
		7298 => '0',
		7299 => '0',
		7300 => '0',
		7301 => '0',
		7302 => '0',
		7303 => '0',
		7304 => '0',
		7305 => '0',
		7306 => '0',
		7307 => '0',
		7308 => '0',
		7309 => '0',
		7310 => '1',
		7311 => '1',
		7312 => '1',
		7313 => '1',
		7314 => '1',
		7315 => '1',
		7316 => '0',
		7317 => '1',
		7318 => '1',
		7319 => '0',
		7320 => '1',
		7321 => '0',
		7322 => '0',
		7323 => '0',
		7324 => '0',
		7325 => '0',
		7326 => '0',
		7327 => '0',
		7328 => '0',
		7329 => '0',
		7330 => '0',
		7331 => '0',
		7332 => '0',
		7333 => '0',
		7334 => '0',
		7335 => '0',
		7336 => '0',
		7337 => '0',
		7338 => '0',
		7339 => '0',
		7340 => '0',
		7341 => '0',
		7342 => '0',
		7343 => '0',
		7344 => '0',
		7345 => '0',
		7346 => '0',
		7347 => '0',
		7348 => '0',
		7349 => '0',
		7350 => '0',
		7351 => '0',
		7352 => '0',
		7353 => '0',
		7354 => '0',
		7355 => '0',
		7356 => '0',
		7357 => '0',
		7358 => '0',
		7359 => '0',
		7360 => '0',
		7361 => '0',
		7362 => '0',
		7363 => '0',
		7364 => '0',
		7365 => '0',
		7366 => '0',
		7367 => '0',
		7368 => '0',
		7369 => '0',
		7370 => '0',
		7371 => '0',
		7372 => '0',
		7373 => '0',
		7374 => '0',
		7375 => '0',
		7376 => '0',
		7377 => '0',
		7378 => '0',
		7379 => '0',
		7380 => '0',
		7381 => '0',
		7382 => '0',
		7383 => '0',
		7384 => '0',
		7385 => '0',
		7386 => '0',
		7387 => '0',
		7388 => '0',
		7389 => '0',
		7390 => '0',
		7391 => '0',
		7392 => '0',
		7393 => '0',
		7394 => '0',
		7395 => '0',
		7396 => '1',
		7397 => '1',
		7398 => '1',
		7399 => '1',
		7400 => '1',
		7401 => '1',
		7402 => '0',
		7403 => '1',
		7404 => '1',
		7405 => '0',
		7406 => '0',
		7407 => '0',
		7408 => '0',
		7409 => '0',
		7410 => '0',
		7411 => '0',
		7412 => '0',
		7413 => '0',
		7414 => '0',
		7415 => '0',
		7424 => '0',
		7425 => '0',
		7426 => '0',
		7427 => '0',
		7428 => '0',
		7429 => '0',
		7430 => '0',
		7431 => '0',
		7432 => '0',
		7433 => '0',
		7434 => '0',
		7435 => '0',
		7436 => '0',
		7437 => '0',
		7438 => '1',
		7439 => '1',
		7440 => '1',
		7441 => '1',
		7442 => '1',
		7443 => '1',
		7444 => '0',
		7445 => '1',
		7446 => '0',
		7447 => '0',
		7448 => '1',
		7449 => '0',
		7450 => '0',
		7451 => '0',
		7452 => '0',
		7453 => '0',
		7454 => '0',
		7455 => '0',
		7456 => '0',
		7457 => '0',
		7458 => '0',
		7459 => '0',
		7460 => '0',
		7461 => '0',
		7462 => '0',
		7463 => '0',
		7464 => '0',
		7465 => '0',
		7466 => '0',
		7467 => '0',
		7468 => '0',
		7469 => '0',
		7470 => '0',
		7471 => '0',
		7472 => '0',
		7473 => '0',
		7474 => '0',
		7475 => '0',
		7476 => '0',
		7477 => '0',
		7478 => '0',
		7479 => '0',
		7480 => '0',
		7481 => '0',
		7482 => '0',
		7483 => '0',
		7484 => '0',
		7485 => '0',
		7486 => '0',
		7487 => '0',
		7488 => '0',
		7489 => '0',
		7490 => '0',
		7491 => '0',
		7492 => '0',
		7493 => '0',
		7494 => '0',
		7495 => '0',
		7496 => '0',
		7497 => '0',
		7498 => '0',
		7499 => '0',
		7500 => '0',
		7501 => '0',
		7502 => '0',
		7503 => '0',
		7504 => '0',
		7505 => '0',
		7506 => '0',
		7507 => '0',
		7508 => '0',
		7509 => '0',
		7510 => '0',
		7511 => '0',
		7512 => '0',
		7513 => '0',
		7514 => '0',
		7515 => '0',
		7516 => '0',
		7517 => '0',
		7518 => '0',
		7519 => '0',
		7520 => '0',
		7521 => '0',
		7522 => '0',
		7523 => '0',
		7524 => '1',
		7525 => '1',
		7526 => '1',
		7527 => '1',
		7528 => '1',
		7529 => '1',
		7530 => '0',
		7531 => '1',
		7532 => '0',
		7533 => '0',
		7534 => '0',
		7535 => '0',
		7536 => '0',
		7537 => '0',
		7538 => '0',
		7539 => '0',
		7540 => '0',
		7541 => '0',
		7542 => '0',
		7543 => '0',
		7552 => '0',
		7553 => '0',
		7554 => '0',
		7555 => '0',
		7556 => '0',
		7557 => '0',
		7558 => '0',
		7559 => '0',
		7560 => '0',
		7561 => '0',
		7562 => '0',
		7563 => '0',
		7564 => '0',
		7565 => '0',
		7566 => '1',
		7567 => '1',
		7568 => '1',
		7569 => '1',
		7570 => '1',
		7571 => '1',
		7572 => '0',
		7573 => '1',
		7574 => '0',
		7575 => '0',
		7576 => '1',
		7577 => '0',
		7578 => '0',
		7579 => '0',
		7580 => '0',
		7581 => '0',
		7582 => '0',
		7583 => '0',
		7584 => '0',
		7585 => '0',
		7586 => '0',
		7587 => '0',
		7588 => '0',
		7589 => '0',
		7590 => '0',
		7591 => '0',
		7592 => '0',
		7593 => '0',
		7594 => '0',
		7595 => '0',
		7596 => '0',
		7597 => '0',
		7598 => '0',
		7599 => '0',
		7600 => '0',
		7601 => '0',
		7602 => '0',
		7603 => '0',
		7604 => '0',
		7605 => '0',
		7606 => '0',
		7607 => '0',
		7608 => '0',
		7609 => '0',
		7610 => '0',
		7611 => '0',
		7612 => '0',
		7613 => '0',
		7614 => '0',
		7615 => '0',
		7616 => '0',
		7617 => '0',
		7618 => '0',
		7619 => '0',
		7620 => '0',
		7621 => '0',
		7622 => '0',
		7623 => '0',
		7624 => '0',
		7625 => '0',
		7626 => '0',
		7627 => '0',
		7628 => '0',
		7629 => '0',
		7630 => '0',
		7631 => '0',
		7632 => '0',
		7633 => '0',
		7634 => '0',
		7635 => '0',
		7636 => '0',
		7637 => '0',
		7638 => '0',
		7639 => '0',
		7640 => '0',
		7641 => '0',
		7642 => '0',
		7643 => '0',
		7644 => '0',
		7645 => '0',
		7646 => '0',
		7647 => '0',
		7648 => '0',
		7649 => '0',
		7650 => '0',
		7651 => '0',
		7652 => '1',
		7653 => '1',
		7654 => '1',
		7655 => '1',
		7656 => '1',
		7657 => '1',
		7658 => '0',
		7659 => '1',
		7660 => '0',
		7661 => '1',
		7662 => '0',
		7663 => '0',
		7664 => '0',
		7665 => '0',
		7666 => '0',
		7667 => '0',
		7668 => '0',
		7669 => '0',
		7670 => '0',
		7671 => '0',
		7680 => '0',
		7681 => '0',
		7682 => '0',
		7683 => '0',
		7684 => '0',
		7685 => '0',
		7686 => '0',
		7687 => '0',
		7688 => '0',
		7689 => '0',
		7690 => '0',
		7691 => '0',
		7692 => '0',
		7693 => '0',
		7694 => '1',
		7695 => '1',
		7696 => '1',
		7697 => '1',
		7698 => '1',
		7699 => '1',
		7700 => '0',
		7701 => '1',
		7702 => '0',
		7703 => '1',
		7704 => '1',
		7705 => '0',
		7706 => '0',
		7707 => '0',
		7708 => '0',
		7709 => '0',
		7710 => '0',
		7711 => '0',
		7712 => '0',
		7713 => '0',
		7714 => '0',
		7715 => '0',
		7716 => '0',
		7717 => '0',
		7718 => '0',
		7719 => '0',
		7720 => '0',
		7721 => '0',
		7722 => '0',
		7723 => '0',
		7724 => '0',
		7725 => '0',
		7726 => '0',
		7727 => '0',
		7728 => '0',
		7729 => '0',
		7730 => '0',
		7731 => '0',
		7732 => '0',
		7733 => '0',
		7734 => '0',
		7735 => '0',
		7736 => '0',
		7737 => '0',
		7738 => '0',
		7739 => '0',
		7740 => '0',
		7741 => '0',
		7742 => '0',
		7743 => '0',
		7744 => '0',
		7745 => '0',
		7746 => '0',
		7747 => '0',
		7748 => '0',
		7749 => '0',
		7750 => '0',
		7751 => '0',
		7752 => '0',
		7753 => '0',
		7754 => '0',
		7755 => '0',
		7756 => '0',
		7757 => '0',
		7758 => '0',
		7759 => '0',
		7760 => '0',
		7761 => '0',
		7762 => '0',
		7763 => '0',
		7764 => '0',
		7765 => '0',
		7766 => '0',
		7767 => '0',
		7768 => '0',
		7769 => '0',
		7770 => '0',
		7771 => '0',
		7772 => '0',
		7773 => '0',
		7774 => '0',
		7775 => '0',
		7776 => '0',
		7777 => '0',
		7778 => '0',
		7779 => '0',
		7780 => '1',
		7781 => '1',
		7782 => '1',
		7783 => '1',
		7784 => '1',
		7785 => '1',
		7786 => '0',
		7787 => '1',
		7788 => '0',
		7789 => '1',
		7790 => '0',
		7791 => '0',
		7792 => '0',
		7793 => '0',
		7794 => '0',
		7795 => '0',
		7796 => '0',
		7797 => '0',
		7798 => '0',
		7799 => '0',
		7808 => '0',
		7809 => '0',
		7810 => '0',
		7811 => '0',
		7812 => '0',
		7813 => '0',
		7814 => '0',
		7815 => '0',
		7816 => '0',
		7817 => '0',
		7818 => '0',
		7819 => '0',
		7820 => '0',
		7821 => '0',
		7822 => '1',
		7823 => '1',
		7824 => '1',
		7825 => '1',
		7826 => '1',
		7827 => '1',
		7828 => '0',
		7829 => '1',
		7830 => '0',
		7831 => '1',
		7832 => '0',
		7833 => '0',
		7834 => '0',
		7835 => '0',
		7836 => '0',
		7837 => '0',
		7838 => '0',
		7839 => '0',
		7840 => '0',
		7841 => '0',
		7842 => '0',
		7843 => '0',
		7844 => '0',
		7845 => '0',
		7846 => '0',
		7847 => '0',
		7848 => '0',
		7849 => '0',
		7850 => '0',
		7851 => '0',
		7852 => '0',
		7853 => '0',
		7854 => '0',
		7855 => '0',
		7856 => '0',
		7857 => '0',
		7858 => '0',
		7859 => '0',
		7860 => '0',
		7861 => '0',
		7862 => '0',
		7863 => '0',
		7864 => '0',
		7865 => '0',
		7866 => '0',
		7867 => '0',
		7868 => '0',
		7869 => '0',
		7870 => '0',
		7871 => '0',
		7872 => '0',
		7873 => '0',
		7874 => '0',
		7875 => '0',
		7876 => '0',
		7877 => '0',
		7878 => '0',
		7879 => '0',
		7880 => '0',
		7881 => '0',
		7882 => '0',
		7883 => '0',
		7884 => '0',
		7885 => '0',
		7886 => '0',
		7887 => '0',
		7888 => '0',
		7889 => '0',
		7890 => '0',
		7891 => '0',
		7892 => '0',
		7893 => '0',
		7894 => '0',
		7895 => '0',
		7896 => '0',
		7897 => '0',
		7898 => '0',
		7899 => '0',
		7900 => '0',
		7901 => '0',
		7902 => '0',
		7903 => '0',
		7904 => '0',
		7905 => '0',
		7906 => '0',
		7907 => '0',
		7908 => '1',
		7909 => '1',
		7910 => '1',
		7911 => '1',
		7912 => '1',
		7913 => '1',
		7914 => '0',
		7915 => '1',
		7916 => '0',
		7917 => '1',
		7918 => '0',
		7919 => '0',
		7920 => '0',
		7921 => '0',
		7922 => '0',
		7923 => '0',
		7924 => '0',
		7925 => '0',
		7926 => '0',
		7927 => '0',
		7936 => '0',
		7937 => '0',
		7938 => '0',
		7939 => '0',
		7940 => '0',
		7941 => '0',
		7942 => '0',
		7943 => '0',
		7944 => '0',
		7945 => '0',
		7946 => '0',
		7947 => '0',
		7948 => '0',
		7949 => '0',
		7950 => '1',
		7951 => '1',
		7952 => '1',
		7953 => '1',
		7954 => '1',
		7955 => '1',
		7956 => '0',
		7957 => '1',
		7958 => '0',
		7959 => '1',
		7960 => '0',
		7961 => '0',
		7962 => '0',
		7963 => '0',
		7964 => '0',
		7965 => '0',
		7966 => '0',
		7967 => '0',
		7968 => '0',
		7969 => '0',
		7970 => '0',
		7971 => '0',
		7972 => '0',
		7973 => '0',
		7974 => '0',
		7975 => '0',
		7976 => '0',
		7977 => '0',
		7978 => '0',
		7979 => '0',
		7980 => '0',
		7981 => '0',
		7982 => '0',
		7983 => '0',
		7984 => '0',
		7985 => '0',
		7986 => '0',
		7987 => '0',
		7988 => '0',
		7989 => '0',
		7990 => '0',
		7991 => '0',
		7992 => '0',
		7993 => '0',
		7994 => '0',
		7995 => '0',
		7996 => '0',
		7997 => '0',
		7998 => '0',
		7999 => '0',
		8000 => '0',
		8001 => '0',
		8002 => '0',
		8003 => '0',
		8004 => '0',
		8005 => '0',
		8006 => '0',
		8007 => '0',
		8008 => '0',
		8009 => '0',
		8010 => '0',
		8011 => '0',
		8012 => '0',
		8013 => '0',
		8014 => '0',
		8015 => '0',
		8016 => '0',
		8017 => '0',
		8018 => '0',
		8019 => '0',
		8020 => '0',
		8021 => '0',
		8022 => '0',
		8023 => '0',
		8024 => '0',
		8025 => '0',
		8026 => '0',
		8027 => '0',
		8028 => '0',
		8029 => '0',
		8030 => '0',
		8031 => '0',
		8032 => '0',
		8033 => '0',
		8034 => '0',
		8035 => '0',
		8036 => '1',
		8037 => '1',
		8038 => '1',
		8039 => '1',
		8040 => '1',
		8041 => '1',
		8042 => '0',
		8043 => '1',
		8044 => '0',
		8045 => '1',
		8046 => '0',
		8047 => '0',
		8048 => '0',
		8049 => '0',
		8050 => '0',
		8051 => '0',
		8052 => '0',
		8053 => '0',
		8054 => '0',
		8055 => '0',
		8064 => '0',
		8065 => '0',
		8066 => '0',
		8067 => '0',
		8068 => '0',
		8069 => '0',
		8070 => '0',
		8071 => '0',
		8072 => '0',
		8073 => '0',
		8074 => '0',
		8075 => '0',
		8076 => '0',
		8077 => '0',
		8078 => '1',
		8079 => '1',
		8080 => '1',
		8081 => '1',
		8082 => '1',
		8083 => '1',
		8084 => '0',
		8085 => '1',
		8086 => '0',
		8087 => '1',
		8088 => '0',
		8089 => '0',
		8090 => '0',
		8091 => '0',
		8092 => '0',
		8093 => '0',
		8094 => '0',
		8095 => '0',
		8096 => '0',
		8097 => '0',
		8098 => '0',
		8099 => '0',
		8100 => '0',
		8101 => '0',
		8102 => '0',
		8103 => '0',
		8104 => '0',
		8105 => '0',
		8106 => '0',
		8107 => '0',
		8108 => '0',
		8109 => '0',
		8110 => '0',
		8111 => '0',
		8112 => '0',
		8113 => '0',
		8114 => '0',
		8115 => '0',
		8116 => '0',
		8117 => '0',
		8118 => '0',
		8119 => '0',
		8120 => '0',
		8121 => '0',
		8122 => '0',
		8123 => '0',
		8124 => '0',
		8125 => '0',
		8126 => '0',
		8127 => '0',
		8128 => '0',
		8129 => '0',
		8130 => '0',
		8131 => '0',
		8132 => '0',
		8133 => '0',
		8134 => '0',
		8135 => '0',
		8136 => '0',
		8137 => '0',
		8138 => '0',
		8139 => '0',
		8140 => '0',
		8141 => '0',
		8142 => '0',
		8143 => '0',
		8144 => '0',
		8145 => '0',
		8146 => '0',
		8147 => '0',
		8148 => '0',
		8149 => '0',
		8150 => '0',
		8151 => '0',
		8152 => '0',
		8153 => '0',
		8154 => '0',
		8155 => '0',
		8156 => '0',
		8157 => '0',
		8158 => '0',
		8159 => '0',
		8160 => '0',
		8161 => '0',
		8162 => '0',
		8163 => '0',
		8164 => '1',
		8165 => '1',
		8166 => '1',
		8167 => '1',
		8168 => '1',
		8169 => '1',
		8170 => '0',
		8171 => '1',
		8172 => '0',
		8173 => '1',
		8174 => '0',
		8175 => '0',
		8176 => '0',
		8177 => '0',
		8178 => '0',
		8179 => '0',
		8180 => '0',
		8181 => '0',
		8182 => '0',
		8183 => '0',
		8192 => '0',
		8193 => '0',
		8194 => '0',
		8195 => '0',
		8196 => '0',
		8197 => '0',
		8198 => '0',
		8199 => '0',
		8200 => '0',
		8201 => '0',
		8202 => '0',
		8203 => '0',
		8204 => '0',
		8205 => '0',
		8206 => '1',
		8207 => '1',
		8208 => '1',
		8209 => '1',
		8210 => '1',
		8211 => '1',
		8212 => '0',
		8213 => '1',
		8214 => '0',
		8215 => '1',
		8216 => '0',
		8217 => '0',
		8218 => '0',
		8219 => '0',
		8220 => '0',
		8221 => '0',
		8222 => '0',
		8223 => '0',
		8224 => '0',
		8225 => '0',
		8226 => '0',
		8227 => '0',
		8228 => '0',
		8229 => '0',
		8230 => '0',
		8231 => '0',
		8232 => '0',
		8233 => '0',
		8234 => '0',
		8235 => '0',
		8236 => '0',
		8237 => '0',
		8238 => '0',
		8239 => '0',
		8240 => '0',
		8241 => '0',
		8242 => '0',
		8243 => '0',
		8244 => '0',
		8245 => '0',
		8246 => '0',
		8247 => '0',
		8248 => '0',
		8249 => '0',
		8250 => '0',
		8251 => '0',
		8252 => '0',
		8253 => '0',
		8254 => '0',
		8255 => '0',
		8256 => '0',
		8257 => '0',
		8258 => '0',
		8259 => '0',
		8260 => '0',
		8261 => '0',
		8262 => '0',
		8263 => '0',
		8264 => '0',
		8265 => '0',
		8266 => '0',
		8267 => '0',
		8268 => '0',
		8269 => '0',
		8270 => '0',
		8271 => '0',
		8272 => '0',
		8273 => '0',
		8274 => '0',
		8275 => '0',
		8276 => '0',
		8277 => '0',
		8278 => '0',
		8279 => '0',
		8280 => '0',
		8281 => '0',
		8282 => '0',
		8283 => '0',
		8284 => '0',
		8285 => '0',
		8286 => '0',
		8287 => '0',
		8288 => '0',
		8289 => '0',
		8290 => '0',
		8291 => '0',
		8292 => '1',
		8293 => '1',
		8294 => '1',
		8295 => '1',
		8296 => '1',
		8297 => '1',
		8298 => '0',
		8299 => '1',
		8300 => '0',
		8301 => '1',
		8302 => '0',
		8303 => '0',
		8304 => '0',
		8305 => '0',
		8306 => '0',
		8307 => '0',
		8308 => '0',
		8309 => '0',
		8310 => '0',
		8311 => '0',
		8320 => '0',
		8321 => '0',
		8322 => '0',
		8323 => '0',
		8324 => '0',
		8325 => '0',
		8326 => '0',
		8327 => '0',
		8328 => '0',
		8329 => '0',
		8330 => '0',
		8331 => '0',
		8332 => '0',
		8333 => '0',
		8334 => '1',
		8335 => '1',
		8336 => '1',
		8337 => '1',
		8338 => '1',
		8339 => '1',
		8340 => '0',
		8341 => '1',
		8342 => '0',
		8343 => '1',
		8344 => '0',
		8345 => '0',
		8346 => '0',
		8347 => '0',
		8348 => '0',
		8349 => '0',
		8350 => '0',
		8351 => '0',
		8352 => '0',
		8353 => '0',
		8354 => '0',
		8355 => '0',
		8356 => '0',
		8357 => '0',
		8358 => '0',
		8359 => '0',
		8360 => '0',
		8361 => '0',
		8362 => '0',
		8363 => '0',
		8364 => '0',
		8365 => '0',
		8366 => '0',
		8367 => '0',
		8368 => '0',
		8369 => '0',
		8370 => '0',
		8371 => '0',
		8372 => '0',
		8373 => '0',
		8374 => '0',
		8375 => '0',
		8376 => '0',
		8377 => '0',
		8378 => '0',
		8379 => '0',
		8380 => '0',
		8381 => '0',
		8382 => '0',
		8383 => '0',
		8384 => '0',
		8385 => '0',
		8386 => '0',
		8387 => '0',
		8388 => '0',
		8389 => '0',
		8390 => '0',
		8391 => '0',
		8392 => '0',
		8393 => '0',
		8394 => '0',
		8395 => '0',
		8396 => '0',
		8397 => '0',
		8398 => '0',
		8399 => '0',
		8400 => '0',
		8401 => '0',
		8402 => '0',
		8403 => '0',
		8404 => '0',
		8405 => '0',
		8406 => '0',
		8407 => '0',
		8408 => '0',
		8409 => '0',
		8410 => '0',
		8411 => '0',
		8412 => '0',
		8413 => '0',
		8414 => '0',
		8415 => '0',
		8416 => '0',
		8417 => '0',
		8418 => '0',
		8419 => '0',
		8420 => '1',
		8421 => '1',
		8422 => '1',
		8423 => '1',
		8424 => '1',
		8425 => '1',
		8426 => '0',
		8427 => '1',
		8428 => '0',
		8429 => '1',
		8430 => '0',
		8431 => '0',
		8432 => '0',
		8433 => '0',
		8434 => '0',
		8435 => '0',
		8436 => '0',
		8437 => '0',
		8438 => '0',
		8439 => '0',
		8448 => '0',
		8449 => '0',
		8450 => '0',
		8451 => '0',
		8452 => '0',
		8453 => '0',
		8454 => '0',
		8455 => '0',
		8456 => '0',
		8457 => '0',
		8458 => '0',
		8459 => '0',
		8460 => '0',
		8461 => '0',
		8462 => '1',
		8463 => '1',
		8464 => '1',
		8465 => '1',
		8466 => '1',
		8467 => '1',
		8468 => '1',
		8469 => '1',
		8470 => '0',
		8471 => '1',
		8472 => '0',
		8473 => '0',
		8474 => '0',
		8475 => '0',
		8476 => '0',
		8477 => '0',
		8478 => '0',
		8479 => '0',
		8480 => '0',
		8481 => '0',
		8482 => '0',
		8483 => '0',
		8484 => '0',
		8485 => '0',
		8486 => '0',
		8487 => '0',
		8488 => '0',
		8489 => '0',
		8490 => '0',
		8491 => '0',
		8492 => '0',
		8493 => '0',
		8494 => '0',
		8495 => '0',
		8496 => '0',
		8497 => '0',
		8498 => '0',
		8499 => '0',
		8500 => '0',
		8501 => '0',
		8502 => '0',
		8503 => '0',
		8504 => '0',
		8505 => '0',
		8506 => '0',
		8507 => '0',
		8508 => '0',
		8509 => '0',
		8510 => '0',
		8511 => '0',
		8512 => '0',
		8513 => '0',
		8514 => '0',
		8515 => '0',
		8516 => '0',
		8517 => '0',
		8518 => '0',
		8519 => '0',
		8520 => '0',
		8521 => '0',
		8522 => '0',
		8523 => '0',
		8524 => '0',
		8525 => '0',
		8526 => '0',
		8527 => '0',
		8528 => '0',
		8529 => '0',
		8530 => '0',
		8531 => '0',
		8532 => '0',
		8533 => '0',
		8534 => '0',
		8535 => '0',
		8536 => '0',
		8537 => '0',
		8538 => '0',
		8539 => '0',
		8540 => '0',
		8541 => '0',
		8542 => '0',
		8543 => '0',
		8544 => '0',
		8545 => '0',
		8546 => '0',
		8547 => '1',
		8548 => '1',
		8549 => '1',
		8550 => '1',
		8551 => '1',
		8552 => '1',
		8553 => '1',
		8554 => '0',
		8555 => '1',
		8556 => '0',
		8557 => '1',
		8558 => '0',
		8559 => '0',
		8560 => '0',
		8561 => '0',
		8562 => '0',
		8563 => '0',
		8564 => '0',
		8565 => '0',
		8566 => '0',
		8567 => '0',
		8576 => '0',
		8577 => '0',
		8578 => '0',
		8579 => '0',
		8580 => '0',
		8581 => '0',
		8582 => '0',
		8583 => '0',
		8584 => '0',
		8585 => '0',
		8586 => '0',
		8587 => '0',
		8588 => '0',
		8589 => '0',
		8590 => '1',
		8591 => '1',
		8592 => '1',
		8593 => '1',
		8594 => '1',
		8595 => '1',
		8596 => '1',
		8597 => '1',
		8598 => '0',
		8599 => '1',
		8600 => '0',
		8601 => '0',
		8602 => '0',
		8603 => '0',
		8604 => '0',
		8605 => '0',
		8606 => '0',
		8607 => '0',
		8608 => '0',
		8609 => '0',
		8610 => '0',
		8611 => '0',
		8612 => '0',
		8613 => '0',
		8614 => '0',
		8615 => '0',
		8616 => '0',
		8617 => '0',
		8618 => '0',
		8619 => '0',
		8620 => '0',
		8621 => '0',
		8622 => '0',
		8623 => '0',
		8624 => '0',
		8625 => '0',
		8626 => '0',
		8627 => '0',
		8628 => '0',
		8629 => '0',
		8630 => '0',
		8631 => '0',
		8632 => '0',
		8633 => '0',
		8634 => '0',
		8635 => '0',
		8636 => '0',
		8637 => '0',
		8638 => '0',
		8639 => '0',
		8640 => '0',
		8641 => '0',
		8642 => '0',
		8643 => '0',
		8644 => '0',
		8645 => '0',
		8646 => '0',
		8647 => '0',
		8648 => '0',
		8649 => '0',
		8650 => '0',
		8651 => '0',
		8652 => '0',
		8653 => '0',
		8654 => '0',
		8655 => '0',
		8656 => '0',
		8657 => '0',
		8658 => '0',
		8659 => '0',
		8660 => '0',
		8661 => '0',
		8662 => '0',
		8663 => '0',
		8664 => '0',
		8665 => '0',
		8666 => '0',
		8667 => '0',
		8668 => '0',
		8669 => '0',
		8670 => '0',
		8671 => '0',
		8672 => '0',
		8673 => '0',
		8674 => '0',
		8675 => '1',
		8676 => '1',
		8677 => '1',
		8678 => '1',
		8679 => '1',
		8680 => '1',
		8681 => '1',
		8682 => '0',
		8683 => '1',
		8684 => '0',
		8685 => '1',
		8686 => '0',
		8687 => '0',
		8688 => '0',
		8689 => '0',
		8690 => '0',
		8691 => '0',
		8692 => '0',
		8693 => '0',
		8694 => '0',
		8695 => '0',
		8704 => '0',
		8705 => '0',
		8706 => '0',
		8707 => '0',
		8708 => '0',
		8709 => '0',
		8710 => '0',
		8711 => '0',
		8712 => '0',
		8713 => '0',
		8714 => '0',
		8715 => '0',
		8716 => '0',
		8717 => '0',
		8718 => '0',
		8719 => '1',
		8720 => '1',
		8721 => '1',
		8722 => '1',
		8723 => '1',
		8724 => '1',
		8725 => '0',
		8726 => '0',
		8727 => '1',
		8728 => '0',
		8729 => '0',
		8730 => '0',
		8731 => '0',
		8732 => '0',
		8733 => '0',
		8734 => '0',
		8735 => '0',
		8736 => '0',
		8737 => '0',
		8738 => '0',
		8739 => '0',
		8740 => '0',
		8741 => '0',
		8742 => '0',
		8743 => '0',
		8744 => '0',
		8745 => '0',
		8746 => '0',
		8747 => '0',
		8748 => '0',
		8749 => '0',
		8750 => '0',
		8751 => '0',
		8752 => '0',
		8753 => '0',
		8754 => '0',
		8755 => '0',
		8756 => '0',
		8757 => '0',
		8758 => '0',
		8759 => '0',
		8760 => '0',
		8761 => '0',
		8762 => '0',
		8763 => '0',
		8764 => '0',
		8765 => '0',
		8766 => '0',
		8767 => '0',
		8768 => '0',
		8769 => '0',
		8770 => '0',
		8771 => '0',
		8772 => '0',
		8773 => '0',
		8774 => '0',
		8775 => '0',
		8776 => '0',
		8777 => '0',
		8778 => '0',
		8779 => '0',
		8780 => '0',
		8781 => '0',
		8782 => '0',
		8783 => '0',
		8784 => '0',
		8785 => '0',
		8786 => '0',
		8787 => '0',
		8788 => '0',
		8789 => '0',
		8790 => '0',
		8791 => '0',
		8792 => '0',
		8793 => '0',
		8794 => '0',
		8795 => '0',
		8796 => '0',
		8797 => '0',
		8798 => '0',
		8799 => '0',
		8800 => '0',
		8801 => '0',
		8802 => '0',
		8803 => '1',
		8804 => '1',
		8805 => '1',
		8806 => '1',
		8807 => '1',
		8808 => '1',
		8809 => '0',
		8810 => '0',
		8811 => '1',
		8812 => '0',
		8813 => '1',
		8814 => '0',
		8815 => '0',
		8816 => '0',
		8817 => '0',
		8818 => '0',
		8819 => '0',
		8820 => '0',
		8821 => '0',
		8822 => '0',
		8823 => '0',
		8832 => '0',
		8833 => '0',
		8834 => '0',
		8835 => '0',
		8836 => '0',
		8837 => '0',
		8838 => '0',
		8839 => '0',
		8840 => '0',
		8841 => '0',
		8842 => '0',
		8843 => '0',
		8844 => '0',
		8845 => '0',
		8846 => '1',
		8847 => '1',
		8848 => '1',
		8849 => '1',
		8850 => '1',
		8851 => '1',
		8852 => '1',
		8853 => '0',
		8854 => '0',
		8855 => '1',
		8856 => '0',
		8857 => '0',
		8858 => '0',
		8859 => '0',
		8860 => '0',
		8861 => '0',
		8862 => '0',
		8863 => '0',
		8864 => '0',
		8865 => '0',
		8866 => '0',
		8867 => '0',
		8868 => '0',
		8869 => '0',
		8870 => '0',
		8871 => '0',
		8872 => '0',
		8873 => '0',
		8874 => '0',
		8875 => '0',
		8876 => '0',
		8877 => '0',
		8878 => '0',
		8879 => '0',
		8880 => '0',
		8881 => '0',
		8882 => '0',
		8883 => '0',
		8884 => '0',
		8885 => '0',
		8886 => '0',
		8887 => '0',
		8888 => '0',
		8889 => '0',
		8890 => '0',
		8891 => '0',
		8892 => '0',
		8893 => '0',
		8894 => '0',
		8895 => '0',
		8896 => '0',
		8897 => '0',
		8898 => '0',
		8899 => '0',
		8900 => '0',
		8901 => '0',
		8902 => '0',
		8903 => '0',
		8904 => '0',
		8905 => '0',
		8906 => '0',
		8907 => '0',
		8908 => '0',
		8909 => '0',
		8910 => '0',
		8911 => '0',
		8912 => '0',
		8913 => '0',
		8914 => '0',
		8915 => '0',
		8916 => '0',
		8917 => '0',
		8918 => '0',
		8919 => '0',
		8920 => '0',
		8921 => '0',
		8922 => '0',
		8923 => '0',
		8924 => '0',
		8925 => '0',
		8926 => '0',
		8927 => '0',
		8928 => '0',
		8929 => '0',
		8930 => '0',
		8931 => '1',
		8932 => '1',
		8933 => '1',
		8934 => '1',
		8935 => '1',
		8936 => '1',
		8937 => '0',
		8938 => '0',
		8939 => '1',
		8940 => '0',
		8941 => '1',
		8942 => '0',
		8943 => '0',
		8944 => '0',
		8945 => '0',
		8946 => '0',
		8947 => '0',
		8948 => '0',
		8949 => '0',
		8950 => '0',
		8951 => '0',
		8960 => '0',
		8961 => '0',
		8962 => '0',
		8963 => '0',
		8964 => '0',
		8965 => '0',
		8966 => '0',
		8967 => '0',
		8968 => '0',
		8969 => '0',
		8970 => '0',
		8971 => '0',
		8972 => '0',
		8973 => '0',
		8974 => '0',
		8975 => '1',
		8976 => '1',
		8977 => '1',
		8978 => '1',
		8979 => '1',
		8980 => '1',
		8981 => '0',
		8982 => '1',
		8983 => '1',
		8984 => '0',
		8985 => '0',
		8986 => '0',
		8987 => '0',
		8988 => '0',
		8989 => '0',
		8990 => '0',
		8991 => '0',
		8992 => '0',
		8993 => '0',
		8994 => '0',
		8995 => '0',
		8996 => '0',
		8997 => '0',
		8998 => '0',
		8999 => '0',
		9000 => '0',
		9001 => '0',
		9002 => '0',
		9003 => '0',
		9004 => '0',
		9005 => '0',
		9006 => '0',
		9007 => '0',
		9008 => '0',
		9009 => '0',
		9010 => '0',
		9011 => '0',
		9012 => '0',
		9013 => '0',
		9014 => '0',
		9015 => '0',
		9016 => '0',
		9017 => '0',
		9018 => '0',
		9019 => '0',
		9020 => '0',
		9021 => '0',
		9022 => '0',
		9023 => '0',
		9024 => '0',
		9025 => '0',
		9026 => '0',
		9027 => '0',
		9028 => '0',
		9029 => '0',
		9030 => '0',
		9031 => '0',
		9032 => '0',
		9033 => '0',
		9034 => '0',
		9035 => '0',
		9036 => '0',
		9037 => '0',
		9038 => '0',
		9039 => '0',
		9040 => '0',
		9041 => '0',
		9042 => '0',
		9043 => '0',
		9044 => '0',
		9045 => '0',
		9046 => '0',
		9047 => '0',
		9048 => '0',
		9049 => '0',
		9050 => '0',
		9051 => '0',
		9052 => '0',
		9053 => '0',
		9054 => '0',
		9055 => '0',
		9056 => '0',
		9057 => '0',
		9058 => '0',
		9059 => '1',
		9060 => '1',
		9061 => '1',
		9062 => '1',
		9063 => '1',
		9064 => '1',
		9065 => '0',
		9066 => '1',
		9067 => '1',
		9068 => '0',
		9069 => '1',
		9070 => '0',
		9071 => '0',
		9072 => '0',
		9073 => '0',
		9074 => '0',
		9075 => '0',
		9076 => '0',
		9077 => '0',
		9078 => '0',
		9079 => '0',
		9088 => '0',
		9089 => '0',
		9090 => '0',
		9091 => '0',
		9092 => '0',
		9093 => '0',
		9094 => '0',
		9095 => '0',
		9096 => '0',
		9097 => '0',
		9098 => '0',
		9099 => '0',
		9100 => '0',
		9101 => '0',
		9102 => '0',
		9103 => '1',
		9104 => '1',
		9105 => '1',
		9106 => '1',
		9107 => '1',
		9108 => '1',
		9109 => '1',
		9110 => '1',
		9111 => '1',
		9112 => '0',
		9113 => '0',
		9114 => '0',
		9115 => '0',
		9116 => '0',
		9117 => '0',
		9118 => '0',
		9119 => '0',
		9120 => '0',
		9121 => '0',
		9122 => '0',
		9123 => '0',
		9124 => '0',
		9125 => '0',
		9126 => '0',
		9127 => '0',
		9128 => '0',
		9129 => '0',
		9130 => '0',
		9131 => '0',
		9132 => '0',
		9133 => '0',
		9134 => '0',
		9135 => '0',
		9136 => '0',
		9137 => '0',
		9138 => '0',
		9139 => '0',
		9140 => '0',
		9141 => '0',
		9142 => '0',
		9143 => '0',
		9144 => '0',
		9145 => '0',
		9146 => '0',
		9147 => '0',
		9148 => '0',
		9149 => '0',
		9150 => '0',
		9151 => '0',
		9152 => '0',
		9153 => '0',
		9154 => '0',
		9155 => '0',
		9156 => '0',
		9157 => '0',
		9158 => '0',
		9159 => '0',
		9160 => '0',
		9161 => '0',
		9162 => '0',
		9163 => '0',
		9164 => '0',
		9165 => '0',
		9166 => '0',
		9167 => '0',
		9168 => '0',
		9169 => '0',
		9170 => '0',
		9171 => '0',
		9172 => '0',
		9173 => '0',
		9174 => '0',
		9175 => '0',
		9176 => '0',
		9177 => '0',
		9178 => '0',
		9179 => '0',
		9180 => '0',
		9181 => '0',
		9182 => '0',
		9183 => '0',
		9184 => '0',
		9185 => '0',
		9186 => '1',
		9187 => '1',
		9188 => '1',
		9189 => '1',
		9190 => '1',
		9191 => '1',
		9192 => '1',
		9193 => '0',
		9194 => '1',
		9195 => '1',
		9196 => '0',
		9197 => '1',
		9198 => '0',
		9199 => '0',
		9200 => '0',
		9201 => '0',
		9202 => '0',
		9203 => '0',
		9204 => '0',
		9205 => '0',
		9206 => '0',
		9207 => '0',
		9216 => '0',
		9217 => '0',
		9218 => '0',
		9219 => '0',
		9220 => '0',
		9221 => '0',
		9222 => '0',
		9223 => '0',
		9224 => '0',
		9225 => '0',
		9226 => '0',
		9227 => '0',
		9228 => '0',
		9229 => '0',
		9230 => '0',
		9231 => '1',
		9232 => '1',
		9233 => '1',
		9234 => '1',
		9235 => '1',
		9236 => '1',
		9237 => '1',
		9238 => '1',
		9239 => '0',
		9240 => '0',
		9241 => '0',
		9242 => '0',
		9243 => '0',
		9244 => '0',
		9245 => '0',
		9246 => '0',
		9247 => '0',
		9248 => '0',
		9249 => '0',
		9250 => '0',
		9251 => '0',
		9252 => '0',
		9253 => '0',
		9254 => '0',
		9255 => '0',
		9256 => '0',
		9257 => '0',
		9258 => '0',
		9259 => '0',
		9260 => '0',
		9261 => '0',
		9262 => '0',
		9263 => '0',
		9264 => '0',
		9265 => '0',
		9266 => '0',
		9267 => '0',
		9268 => '0',
		9269 => '0',
		9270 => '0',
		9271 => '0',
		9272 => '0',
		9273 => '0',
		9274 => '0',
		9275 => '0',
		9276 => '0',
		9277 => '0',
		9278 => '0',
		9279 => '0',
		9280 => '0',
		9281 => '0',
		9282 => '0',
		9283 => '0',
		9284 => '0',
		9285 => '0',
		9286 => '0',
		9287 => '0',
		9288 => '0',
		9289 => '0',
		9290 => '0',
		9291 => '0',
		9292 => '0',
		9293 => '0',
		9294 => '0',
		9295 => '0',
		9296 => '0',
		9297 => '0',
		9298 => '0',
		9299 => '0',
		9300 => '0',
		9301 => '0',
		9302 => '0',
		9303 => '0',
		9304 => '0',
		9305 => '0',
		9306 => '0',
		9307 => '0',
		9308 => '0',
		9309 => '0',
		9310 => '0',
		9311 => '0',
		9312 => '0',
		9313 => '0',
		9314 => '1',
		9315 => '1',
		9316 => '1',
		9317 => '1',
		9318 => '1',
		9319 => '1',
		9320 => '1',
		9321 => '0',
		9322 => '1',
		9323 => '0',
		9324 => '0',
		9325 => '1',
		9326 => '0',
		9327 => '0',
		9328 => '0',
		9329 => '0',
		9330 => '0',
		9331 => '0',
		9332 => '0',
		9333 => '0',
		9334 => '0',
		9335 => '0',
		9344 => '0',
		9345 => '0',
		9346 => '0',
		9347 => '0',
		9348 => '0',
		9349 => '0',
		9350 => '0',
		9351 => '0',
		9352 => '0',
		9353 => '0',
		9354 => '0',
		9355 => '0',
		9356 => '0',
		9357 => '0',
		9358 => '0',
		9359 => '0',
		9360 => '1',
		9361 => '1',
		9362 => '1',
		9363 => '1',
		9364 => '1',
		9365 => '1',
		9366 => '0',
		9367 => '0',
		9368 => '1',
		9369 => '0',
		9370 => '0',
		9371 => '0',
		9372 => '0',
		9373 => '0',
		9374 => '0',
		9375 => '0',
		9376 => '0',
		9377 => '0',
		9378 => '0',
		9379 => '0',
		9380 => '0',
		9381 => '0',
		9382 => '0',
		9383 => '0',
		9384 => '0',
		9385 => '0',
		9386 => '0',
		9387 => '0',
		9388 => '0',
		9389 => '0',
		9390 => '0',
		9391 => '0',
		9392 => '0',
		9393 => '0',
		9394 => '0',
		9395 => '0',
		9396 => '0',
		9397 => '0',
		9398 => '0',
		9399 => '0',
		9400 => '0',
		9401 => '0',
		9402 => '0',
		9403 => '0',
		9404 => '0',
		9405 => '0',
		9406 => '0',
		9407 => '0',
		9408 => '0',
		9409 => '0',
		9410 => '0',
		9411 => '0',
		9412 => '0',
		9413 => '0',
		9414 => '0',
		9415 => '0',
		9416 => '0',
		9417 => '0',
		9418 => '0',
		9419 => '0',
		9420 => '0',
		9421 => '0',
		9422 => '0',
		9423 => '0',
		9424 => '0',
		9425 => '0',
		9426 => '0',
		9427 => '0',
		9428 => '0',
		9429 => '0',
		9430 => '0',
		9431 => '0',
		9432 => '0',
		9433 => '0',
		9434 => '0',
		9435 => '0',
		9436 => '0',
		9437 => '0',
		9438 => '0',
		9439 => '0',
		9440 => '0',
		9441 => '0',
		9442 => '1',
		9443 => '1',
		9444 => '1',
		9445 => '1',
		9446 => '1',
		9447 => '1',
		9448 => '0',
		9449 => '0',
		9450 => '1',
		9451 => '0',
		9452 => '0',
		9453 => '1',
		9454 => '0',
		9455 => '0',
		9456 => '0',
		9457 => '0',
		9458 => '0',
		9459 => '0',
		9460 => '0',
		9461 => '0',
		9462 => '0',
		9463 => '0',
		9472 => '0',
		9473 => '0',
		9474 => '0',
		9475 => '0',
		9476 => '0',
		9477 => '0',
		9478 => '0',
		9479 => '0',
		9480 => '0',
		9481 => '0',
		9482 => '0',
		9483 => '0',
		9484 => '0',
		9485 => '0',
		9486 => '0',
		9487 => '1',
		9488 => '1',
		9489 => '1',
		9490 => '1',
		9491 => '1',
		9492 => '1',
		9493 => '1',
		9494 => '1',
		9495 => '0',
		9496 => '1',
		9497 => '0',
		9498 => '0',
		9499 => '0',
		9500 => '0',
		9501 => '0',
		9502 => '0',
		9503 => '0',
		9504 => '0',
		9505 => '0',
		9506 => '0',
		9507 => '0',
		9508 => '0',
		9509 => '0',
		9510 => '0',
		9511 => '0',
		9512 => '0',
		9513 => '0',
		9514 => '0',
		9515 => '0',
		9516 => '0',
		9517 => '0',
		9518 => '0',
		9519 => '0',
		9520 => '0',
		9521 => '0',
		9522 => '0',
		9523 => '0',
		9524 => '0',
		9525 => '0',
		9526 => '0',
		9527 => '0',
		9528 => '0',
		9529 => '0',
		9530 => '0',
		9531 => '0',
		9532 => '0',
		9533 => '0',
		9534 => '0',
		9535 => '0',
		9536 => '0',
		9537 => '0',
		9538 => '0',
		9539 => '0',
		9540 => '0',
		9541 => '0',
		9542 => '0',
		9543 => '0',
		9544 => '0',
		9545 => '0',
		9546 => '0',
		9547 => '0',
		9548 => '0',
		9549 => '0',
		9550 => '0',
		9551 => '0',
		9552 => '0',
		9553 => '0',
		9554 => '0',
		9555 => '0',
		9556 => '0',
		9557 => '0',
		9558 => '0',
		9559 => '0',
		9560 => '0',
		9561 => '0',
		9562 => '0',
		9563 => '0',
		9564 => '0',
		9565 => '0',
		9566 => '0',
		9567 => '0',
		9568 => '0',
		9569 => '1',
		9570 => '1',
		9571 => '1',
		9572 => '1',
		9573 => '1',
		9574 => '1',
		9575 => '1',
		9576 => '0',
		9577 => '0',
		9578 => '1',
		9579 => '0',
		9580 => '1',
		9581 => '1',
		9582 => '0',
		9583 => '0',
		9584 => '0',
		9585 => '0',
		9586 => '0',
		9587 => '0',
		9588 => '0',
		9589 => '0',
		9590 => '0',
		9591 => '0',
		9600 => '0',
		9601 => '0',
		9602 => '0',
		9603 => '0',
		9604 => '0',
		9605 => '0',
		9606 => '0',
		9607 => '0',
		9608 => '0',
		9609 => '0',
		9610 => '0',
		9611 => '0',
		9612 => '0',
		9613 => '0',
		9614 => '0',
		9615 => '0',
		9616 => '1',
		9617 => '1',
		9618 => '1',
		9619 => '1',
		9620 => '1',
		9621 => '1',
		9622 => '1',
		9623 => '1',
		9624 => '1',
		9625 => '0',
		9626 => '0',
		9627 => '0',
		9628 => '0',
		9629 => '0',
		9630 => '0',
		9631 => '0',
		9632 => '0',
		9633 => '0',
		9634 => '0',
		9635 => '0',
		9636 => '0',
		9637 => '0',
		9638 => '0',
		9639 => '0',
		9640 => '0',
		9641 => '0',
		9642 => '0',
		9643 => '0',
		9644 => '0',
		9645 => '0',
		9646 => '0',
		9647 => '0',
		9648 => '0',
		9649 => '0',
		9650 => '0',
		9651 => '0',
		9652 => '0',
		9653 => '0',
		9654 => '0',
		9655 => '0',
		9656 => '0',
		9657 => '0',
		9658 => '0',
		9659 => '0',
		9660 => '0',
		9661 => '0',
		9662 => '0',
		9663 => '0',
		9664 => '0',
		9665 => '0',
		9666 => '0',
		9667 => '0',
		9668 => '0',
		9669 => '0',
		9670 => '0',
		9671 => '0',
		9672 => '0',
		9673 => '0',
		9674 => '0',
		9675 => '0',
		9676 => '0',
		9677 => '0',
		9678 => '0',
		9679 => '0',
		9680 => '0',
		9681 => '0',
		9682 => '0',
		9683 => '0',
		9684 => '0',
		9685 => '0',
		9686 => '0',
		9687 => '0',
		9688 => '0',
		9689 => '0',
		9690 => '0',
		9691 => '0',
		9692 => '0',
		9693 => '0',
		9694 => '0',
		9695 => '0',
		9696 => '0',
		9697 => '1',
		9698 => '1',
		9699 => '1',
		9700 => '1',
		9701 => '1',
		9702 => '1',
		9703 => '1',
		9704 => '0',
		9705 => '1',
		9706 => '1',
		9707 => '0',
		9708 => '1',
		9709 => '0',
		9710 => '0',
		9711 => '0',
		9712 => '0',
		9713 => '0',
		9714 => '0',
		9715 => '0',
		9716 => '0',
		9717 => '0',
		9718 => '0',
		9719 => '0',
		9728 => '0',
		9729 => '0',
		9730 => '0',
		9731 => '0',
		9732 => '0',
		9733 => '0',
		9734 => '0',
		9735 => '0',
		9736 => '0',
		9737 => '0',
		9738 => '0',
		9739 => '0',
		9740 => '0',
		9741 => '0',
		9742 => '0',
		9743 => '0',
		9744 => '0',
		9745 => '1',
		9746 => '1',
		9747 => '1',
		9748 => '1',
		9749 => '1',
		9750 => '1',
		9751 => '1',
		9752 => '1',
		9753 => '0',
		9754 => '0',
		9755 => '0',
		9756 => '0',
		9757 => '0',
		9758 => '0',
		9759 => '0',
		9760 => '0',
		9761 => '0',
		9762 => '0',
		9763 => '0',
		9764 => '0',
		9765 => '0',
		9766 => '0',
		9767 => '0',
		9768 => '0',
		9769 => '0',
		9770 => '0',
		9771 => '0',
		9772 => '0',
		9773 => '0',
		9774 => '0',
		9775 => '0',
		9776 => '0',
		9777 => '0',
		9778 => '0',
		9779 => '0',
		9780 => '0',
		9781 => '0',
		9782 => '0',
		9783 => '0',
		9784 => '0',
		9785 => '0',
		9786 => '0',
		9787 => '0',
		9788 => '0',
		9789 => '0',
		9790 => '0',
		9791 => '0',
		9792 => '0',
		9793 => '0',
		9794 => '0',
		9795 => '0',
		9796 => '0',
		9797 => '0',
		9798 => '0',
		9799 => '0',
		9800 => '0',
		9801 => '0',
		9802 => '0',
		9803 => '0',
		9804 => '0',
		9805 => '0',
		9806 => '0',
		9807 => '0',
		9808 => '0',
		9809 => '0',
		9810 => '0',
		9811 => '0',
		9812 => '0',
		9813 => '0',
		9814 => '0',
		9815 => '0',
		9816 => '0',
		9817 => '0',
		9818 => '0',
		9819 => '0',
		9820 => '0',
		9821 => '0',
		9822 => '0',
		9823 => '0',
		9824 => '1',
		9825 => '1',
		9826 => '1',
		9827 => '1',
		9828 => '1',
		9829 => '1',
		9830 => '1',
		9831 => '0',
		9832 => '0',
		9833 => '1',
		9834 => '1',
		9835 => '0',
		9836 => '1',
		9837 => '0',
		9838 => '0',
		9839 => '0',
		9840 => '0',
		9841 => '0',
		9842 => '0',
		9843 => '0',
		9844 => '0',
		9845 => '0',
		9846 => '0',
		9847 => '0',
		9856 => '0',
		9857 => '0',
		9858 => '0',
		9859 => '0',
		9860 => '0',
		9861 => '0',
		9862 => '0',
		9863 => '0',
		9864 => '0',
		9865 => '0',
		9866 => '0',
		9867 => '0',
		9868 => '0',
		9869 => '0',
		9870 => '0',
		9871 => '0',
		9872 => '1',
		9873 => '1',
		9874 => '1',
		9875 => '1',
		9876 => '1',
		9877 => '1',
		9878 => '1',
		9879 => '1',
		9880 => '0',
		9881 => '0',
		9882 => '0',
		9883 => '0',
		9884 => '0',
		9885 => '0',
		9886 => '0',
		9887 => '0',
		9888 => '0',
		9889 => '0',
		9890 => '0',
		9891 => '0',
		9892 => '0',
		9893 => '0',
		9894 => '0',
		9895 => '0',
		9896 => '0',
		9897 => '0',
		9898 => '0',
		9899 => '0',
		9900 => '0',
		9901 => '0',
		9902 => '0',
		9903 => '0',
		9904 => '0',
		9905 => '0',
		9906 => '0',
		9907 => '0',
		9908 => '0',
		9909 => '0',
		9910 => '0',
		9911 => '0',
		9912 => '0',
		9913 => '0',
		9914 => '0',
		9915 => '0',
		9916 => '0',
		9917 => '0',
		9918 => '0',
		9919 => '0',
		9920 => '0',
		9921 => '0',
		9922 => '0',
		9923 => '0',
		9924 => '0',
		9925 => '0',
		9926 => '0',
		9927 => '0',
		9928 => '0',
		9929 => '0',
		9930 => '0',
		9931 => '0',
		9932 => '0',
		9933 => '0',
		9934 => '0',
		9935 => '0',
		9936 => '0',
		9937 => '0',
		9938 => '0',
		9939 => '0',
		9940 => '0',
		9941 => '0',
		9942 => '0',
		9943 => '0',
		9944 => '0',
		9945 => '0',
		9946 => '0',
		9947 => '0',
		9948 => '0',
		9949 => '0',
		9950 => '0',
		9951 => '0',
		9952 => '1',
		9953 => '1',
		9954 => '1',
		9955 => '1',
		9956 => '1',
		9957 => '1',
		9958 => '1',
		9959 => '0',
		9960 => '0',
		9961 => '1',
		9962 => '0',
		9963 => '0',
		9964 => '1',
		9965 => '0',
		9966 => '0',
		9967 => '0',
		9968 => '0',
		9969 => '0',
		9970 => '0',
		9971 => '0',
		9972 => '0',
		9973 => '0',
		9974 => '0',
		9975 => '0',
		9984 => '0',
		9985 => '0',
		9986 => '0',
		9987 => '0',
		9988 => '0',
		9989 => '0',
		9990 => '0',
		9991 => '0',
		9992 => '0',
		9993 => '0',
		9994 => '0',
		9995 => '0',
		9996 => '0',
		9997 => '0',
		9998 => '0',
		9999 => '0',
		10000 => '0',
		10001 => '0',
		10002 => '1',
		10003 => '1',
		10004 => '1',
		10005 => '1',
		10006 => '1',
		10007 => '1',
		10008 => '1',
		10009 => '1',
		10010 => '0',
		10011 => '0',
		10012 => '0',
		10013 => '0',
		10014 => '0',
		10015 => '0',
		10016 => '0',
		10017 => '0',
		10018 => '0',
		10019 => '0',
		10020 => '0',
		10021 => '0',
		10022 => '0',
		10023 => '0',
		10024 => '0',
		10025 => '0',
		10026 => '0',
		10027 => '0',
		10028 => '0',
		10029 => '0',
		10030 => '0',
		10031 => '0',
		10032 => '0',
		10033 => '0',
		10034 => '0',
		10035 => '0',
		10036 => '0',
		10037 => '0',
		10038 => '0',
		10039 => '0',
		10040 => '0',
		10041 => '0',
		10042 => '0',
		10043 => '0',
		10044 => '0',
		10045 => '0',
		10046 => '0',
		10047 => '0',
		10048 => '0',
		10049 => '0',
		10050 => '0',
		10051 => '0',
		10052 => '0',
		10053 => '0',
		10054 => '0',
		10055 => '0',
		10056 => '0',
		10057 => '0',
		10058 => '0',
		10059 => '0',
		10060 => '0',
		10061 => '0',
		10062 => '0',
		10063 => '0',
		10064 => '0',
		10065 => '0',
		10066 => '0',
		10067 => '0',
		10068 => '0',
		10069 => '0',
		10070 => '0',
		10071 => '0',
		10072 => '0',
		10073 => '0',
		10074 => '0',
		10075 => '0',
		10076 => '0',
		10077 => '0',
		10078 => '0',
		10079 => '1',
		10080 => '1',
		10081 => '1',
		10082 => '1',
		10083 => '1',
		10084 => '1',
		10085 => '1',
		10086 => '0',
		10087 => '0',
		10088 => '1',
		10089 => '1',
		10090 => '0',
		10091 => '0',
		10092 => '1',
		10093 => '0',
		10094 => '0',
		10095 => '0',
		10096 => '0',
		10097 => '0',
		10098 => '0',
		10099 => '0',
		10100 => '0',
		10101 => '0',
		10102 => '0',
		10103 => '0',
		10112 => '0',
		10113 => '0',
		10114 => '0',
		10115 => '0',
		10116 => '0',
		10117 => '0',
		10118 => '0',
		10119 => '0',
		10120 => '0',
		10121 => '0',
		10122 => '0',
		10123 => '0',
		10124 => '0',
		10125 => '0',
		10126 => '0',
		10127 => '0',
		10128 => '0',
		10129 => '1',
		10130 => '1',
		10131 => '1',
		10132 => '1',
		10133 => '1',
		10134 => '1',
		10135 => '1',
		10136 => '1',
		10137 => '1',
		10138 => '0',
		10139 => '0',
		10140 => '0',
		10141 => '0',
		10142 => '0',
		10143 => '0',
		10144 => '0',
		10145 => '0',
		10146 => '0',
		10147 => '0',
		10148 => '0',
		10149 => '0',
		10150 => '0',
		10151 => '0',
		10152 => '0',
		10153 => '0',
		10154 => '0',
		10155 => '0',
		10156 => '0',
		10157 => '0',
		10158 => '0',
		10159 => '0',
		10160 => '0',
		10161 => '0',
		10162 => '0',
		10163 => '0',
		10164 => '0',
		10165 => '0',
		10166 => '0',
		10167 => '0',
		10168 => '0',
		10169 => '0',
		10170 => '0',
		10171 => '0',
		10172 => '0',
		10173 => '0',
		10174 => '0',
		10175 => '0',
		10176 => '0',
		10177 => '0',
		10178 => '0',
		10179 => '0',
		10180 => '0',
		10181 => '0',
		10182 => '0',
		10183 => '0',
		10184 => '0',
		10185 => '0',
		10186 => '0',
		10187 => '0',
		10188 => '0',
		10189 => '0',
		10190 => '0',
		10191 => '0',
		10192 => '0',
		10193 => '0',
		10194 => '0',
		10195 => '0',
		10196 => '0',
		10197 => '0',
		10198 => '0',
		10199 => '0',
		10200 => '0',
		10201 => '0',
		10202 => '0',
		10203 => '0',
		10204 => '0',
		10205 => '0',
		10206 => '0',
		10207 => '1',
		10208 => '1',
		10209 => '1',
		10210 => '1',
		10211 => '1',
		10212 => '1',
		10213 => '1',
		10214 => '0',
		10215 => '0',
		10216 => '1',
		10217 => '1',
		10218 => '0',
		10219 => '1',
		10220 => '1',
		10221 => '0',
		10222 => '0',
		10223 => '0',
		10224 => '0',
		10225 => '0',
		10226 => '0',
		10227 => '0',
		10228 => '0',
		10229 => '0',
		10230 => '0',
		10231 => '0',
		10240 => '0',
		10241 => '0',
		10242 => '0',
		10243 => '0',
		10244 => '0',
		10245 => '0',
		10246 => '0',
		10247 => '0',
		10248 => '0',
		10249 => '0',
		10250 => '0',
		10251 => '0',
		10252 => '0',
		10253 => '0',
		10254 => '0',
		10255 => '0',
		10256 => '0',
		10257 => '0',
		10258 => '0',
		10259 => '1',
		10260 => '1',
		10261 => '1',
		10262 => '1',
		10263 => '1',
		10264 => '1',
		10265 => '1',
		10266 => '0',
		10267 => '0',
		10268 => '0',
		10269 => '0',
		10270 => '0',
		10271 => '0',
		10272 => '0',
		10273 => '0',
		10274 => '0',
		10275 => '0',
		10276 => '0',
		10277 => '0',
		10278 => '0',
		10279 => '0',
		10280 => '0',
		10281 => '0',
		10282 => '0',
		10283 => '0',
		10284 => '0',
		10285 => '0',
		10286 => '0',
		10287 => '0',
		10288 => '0',
		10289 => '0',
		10290 => '0',
		10291 => '0',
		10292 => '0',
		10293 => '0',
		10294 => '0',
		10295 => '0',
		10296 => '0',
		10297 => '0',
		10298 => '0',
		10299 => '0',
		10300 => '0',
		10301 => '0',
		10302 => '0',
		10303 => '0',
		10304 => '0',
		10305 => '0',
		10306 => '0',
		10307 => '0',
		10308 => '0',
		10309 => '0',
		10310 => '0',
		10311 => '0',
		10312 => '0',
		10313 => '0',
		10314 => '0',
		10315 => '0',
		10316 => '0',
		10317 => '0',
		10318 => '0',
		10319 => '0',
		10320 => '0',
		10321 => '0',
		10322 => '0',
		10323 => '0',
		10324 => '0',
		10325 => '0',
		10326 => '0',
		10327 => '0',
		10328 => '0',
		10329 => '0',
		10330 => '0',
		10331 => '0',
		10332 => '0',
		10333 => '0',
		10334 => '1',
		10335 => '1',
		10336 => '1',
		10337 => '1',
		10338 => '1',
		10339 => '1',
		10340 => '1',
		10341 => '0',
		10342 => '0',
		10343 => '1',
		10344 => '1',
		10345 => '0',
		10346 => '0',
		10347 => '1',
		10348 => '0',
		10349 => '0',
		10350 => '0',
		10351 => '0',
		10352 => '0',
		10353 => '0',
		10354 => '0',
		10355 => '0',
		10356 => '0',
		10357 => '0',
		10358 => '0',
		10359 => '0',
		10368 => '0',
		10369 => '0',
		10370 => '0',
		10371 => '0',
		10372 => '0',
		10373 => '0',
		10374 => '0',
		10375 => '0',
		10376 => '0',
		10377 => '0',
		10378 => '0',
		10379 => '0',
		10380 => '0',
		10381 => '0',
		10382 => '0',
		10383 => '0',
		10384 => '0',
		10385 => '0',
		10386 => '1',
		10387 => '1',
		10388 => '1',
		10389 => '1',
		10390 => '1',
		10391 => '1',
		10392 => '1',
		10393 => '1',
		10394 => '1',
		10395 => '0',
		10396 => '0',
		10397 => '0',
		10398 => '0',
		10399 => '0',
		10400 => '0',
		10401 => '0',
		10402 => '0',
		10403 => '0',
		10404 => '0',
		10405 => '0',
		10406 => '0',
		10407 => '0',
		10408 => '0',
		10409 => '0',
		10410 => '0',
		10411 => '0',
		10412 => '0',
		10413 => '0',
		10414 => '0',
		10415 => '0',
		10416 => '0',
		10417 => '0',
		10418 => '0',
		10419 => '0',
		10420 => '0',
		10421 => '0',
		10422 => '0',
		10423 => '0',
		10424 => '0',
		10425 => '0',
		10426 => '0',
		10427 => '0',
		10428 => '0',
		10429 => '0',
		10430 => '0',
		10431 => '0',
		10432 => '0',
		10433 => '0',
		10434 => '0',
		10435 => '0',
		10436 => '0',
		10437 => '0',
		10438 => '0',
		10439 => '0',
		10440 => '0',
		10441 => '0',
		10442 => '0',
		10443 => '0',
		10444 => '0',
		10445 => '0',
		10446 => '0',
		10447 => '0',
		10448 => '0',
		10449 => '0',
		10450 => '0',
		10451 => '0',
		10452 => '0',
		10453 => '0',
		10454 => '0',
		10455 => '0',
		10456 => '0',
		10457 => '0',
		10458 => '0',
		10459 => '0',
		10460 => '0',
		10461 => '0',
		10462 => '1',
		10463 => '1',
		10464 => '1',
		10465 => '1',
		10466 => '1',
		10467 => '1',
		10468 => '1',
		10469 => '0',
		10470 => '0',
		10471 => '1',
		10472 => '1',
		10473 => '0',
		10474 => '0',
		10475 => '1',
		10476 => '0',
		10477 => '0',
		10478 => '0',
		10479 => '0',
		10480 => '0',
		10481 => '0',
		10482 => '0',
		10483 => '0',
		10484 => '0',
		10485 => '0',
		10486 => '0',
		10487 => '0',
		10496 => '0',
		10497 => '0',
		10498 => '0',
		10499 => '0',
		10500 => '0',
		10501 => '0',
		10502 => '0',
		10503 => '0',
		10504 => '0',
		10505 => '0',
		10506 => '0',
		10507 => '0',
		10508 => '0',
		10509 => '0',
		10510 => '0',
		10511 => '0',
		10512 => '0',
		10513 => '0',
		10514 => '0',
		10515 => '0',
		10516 => '1',
		10517 => '1',
		10518 => '1',
		10519 => '1',
		10520 => '1',
		10521 => '1',
		10522 => '1',
		10523 => '0',
		10524 => '0',
		10525 => '0',
		10526 => '0',
		10527 => '0',
		10528 => '0',
		10529 => '0',
		10530 => '0',
		10531 => '0',
		10532 => '0',
		10533 => '0',
		10534 => '0',
		10535 => '0',
		10536 => '0',
		10537 => '0',
		10538 => '0',
		10539 => '0',
		10540 => '0',
		10541 => '0',
		10542 => '0',
		10543 => '0',
		10544 => '0',
		10545 => '0',
		10546 => '0',
		10547 => '0',
		10548 => '0',
		10549 => '0',
		10550 => '0',
		10551 => '0',
		10552 => '0',
		10553 => '0',
		10554 => '0',
		10555 => '0',
		10556 => '0',
		10557 => '0',
		10558 => '0',
		10559 => '0',
		10560 => '0',
		10561 => '0',
		10562 => '0',
		10563 => '0',
		10564 => '0',
		10565 => '0',
		10566 => '0',
		10567 => '0',
		10568 => '0',
		10569 => '0',
		10570 => '0',
		10571 => '0',
		10572 => '0',
		10573 => '0',
		10574 => '0',
		10575 => '0',
		10576 => '0',
		10577 => '0',
		10578 => '0',
		10579 => '0',
		10580 => '0',
		10581 => '0',
		10582 => '0',
		10583 => '0',
		10584 => '0',
		10585 => '0',
		10586 => '0',
		10587 => '0',
		10588 => '0',
		10589 => '1',
		10590 => '1',
		10591 => '1',
		10592 => '1',
		10593 => '1',
		10594 => '1',
		10595 => '1',
		10596 => '0',
		10597 => '0',
		10598 => '1',
		10599 => '1',
		10600 => '0',
		10601 => '0',
		10602 => '1',
		10603 => '1',
		10604 => '0',
		10605 => '0',
		10606 => '0',
		10607 => '0',
		10608 => '0',
		10609 => '0',
		10610 => '0',
		10611 => '0',
		10612 => '0',
		10613 => '0',
		10614 => '0',
		10615 => '0',
		10624 => '0',
		10625 => '0',
		10626 => '0',
		10627 => '0',
		10628 => '0',
		10629 => '0',
		10630 => '0',
		10631 => '0',
		10632 => '0',
		10633 => '0',
		10634 => '0',
		10635 => '0',
		10636 => '0',
		10637 => '0',
		10638 => '0',
		10639 => '0',
		10640 => '0',
		10641 => '0',
		10642 => '0',
		10643 => '1',
		10644 => '1',
		10645 => '1',
		10646 => '1',
		10647 => '1',
		10648 => '1',
		10649 => '1',
		10650 => '1',
		10651 => '1',
		10652 => '0',
		10653 => '0',
		10654 => '0',
		10655 => '0',
		10656 => '0',
		10657 => '0',
		10658 => '0',
		10659 => '0',
		10660 => '0',
		10661 => '0',
		10662 => '0',
		10663 => '0',
		10664 => '0',
		10665 => '0',
		10666 => '0',
		10667 => '0',
		10668 => '0',
		10669 => '0',
		10670 => '0',
		10671 => '0',
		10672 => '0',
		10673 => '0',
		10674 => '0',
		10675 => '0',
		10676 => '0',
		10677 => '0',
		10678 => '0',
		10679 => '0',
		10680 => '0',
		10681 => '0',
		10682 => '0',
		10683 => '0',
		10684 => '0',
		10685 => '0',
		10686 => '0',
		10687 => '0',
		10688 => '0',
		10689 => '0',
		10690 => '0',
		10691 => '0',
		10692 => '0',
		10693 => '0',
		10694 => '0',
		10695 => '0',
		10696 => '0',
		10697 => '0',
		10698 => '0',
		10699 => '0',
		10700 => '0',
		10701 => '0',
		10702 => '0',
		10703 => '0',
		10704 => '0',
		10705 => '0',
		10706 => '0',
		10707 => '0',
		10708 => '0',
		10709 => '0',
		10710 => '0',
		10711 => '0',
		10712 => '0',
		10713 => '0',
		10714 => '0',
		10715 => '0',
		10716 => '1',
		10717 => '1',
		10718 => '1',
		10719 => '1',
		10720 => '1',
		10721 => '1',
		10722 => '1',
		10723 => '1',
		10724 => '0',
		10725 => '0',
		10726 => '1',
		10727 => '1',
		10728 => '0',
		10729 => '0',
		10730 => '1',
		10731 => '0',
		10732 => '0',
		10733 => '0',
		10734 => '0',
		10735 => '0',
		10736 => '0',
		10737 => '0',
		10738 => '0',
		10739 => '0',
		10740 => '0',
		10741 => '0',
		10742 => '0',
		10743 => '0',
		10752 => '0',
		10753 => '0',
		10754 => '0',
		10755 => '0',
		10756 => '0',
		10757 => '0',
		10758 => '0',
		10759 => '0',
		10760 => '0',
		10761 => '0',
		10762 => '0',
		10763 => '0',
		10764 => '0',
		10765 => '0',
		10766 => '0',
		10767 => '0',
		10768 => '0',
		10769 => '0',
		10770 => '0',
		10771 => '0',
		10772 => '0',
		10773 => '1',
		10774 => '1',
		10775 => '1',
		10776 => '1',
		10777 => '1',
		10778 => '1',
		10779 => '1',
		10780 => '1',
		10781 => '0',
		10782 => '0',
		10783 => '0',
		10784 => '0',
		10785 => '0',
		10786 => '0',
		10787 => '0',
		10788 => '0',
		10789 => '0',
		10790 => '0',
		10791 => '0',
		10792 => '0',
		10793 => '0',
		10794 => '0',
		10795 => '0',
		10796 => '0',
		10797 => '0',
		10798 => '0',
		10799 => '0',
		10800 => '0',
		10801 => '0',
		10802 => '0',
		10803 => '0',
		10804 => '0',
		10805 => '0',
		10806 => '0',
		10807 => '0',
		10808 => '0',
		10809 => '0',
		10810 => '0',
		10811 => '0',
		10812 => '0',
		10813 => '0',
		10814 => '0',
		10815 => '0',
		10816 => '0',
		10817 => '0',
		10818 => '0',
		10819 => '0',
		10820 => '0',
		10821 => '0',
		10822 => '0',
		10823 => '0',
		10824 => '0',
		10825 => '0',
		10826 => '0',
		10827 => '0',
		10828 => '0',
		10829 => '0',
		10830 => '0',
		10831 => '0',
		10832 => '0',
		10833 => '0',
		10834 => '0',
		10835 => '0',
		10836 => '0',
		10837 => '0',
		10838 => '0',
		10839 => '0',
		10840 => '0',
		10841 => '0',
		10842 => '0',
		10843 => '0',
		10844 => '1',
		10845 => '1',
		10846 => '1',
		10847 => '1',
		10848 => '1',
		10849 => '1',
		10850 => '1',
		10851 => '0',
		10852 => '0',
		10853 => '1',
		10854 => '1',
		10855 => '0',
		10856 => '0',
		10857 => '1',
		10858 => '1',
		10859 => '0',
		10860 => '0',
		10861 => '0',
		10862 => '0',
		10863 => '0',
		10864 => '0',
		10865 => '0',
		10866 => '0',
		10867 => '0',
		10868 => '0',
		10869 => '0',
		10870 => '0',
		10871 => '0',
		10880 => '0',
		10881 => '0',
		10882 => '0',
		10883 => '0',
		10884 => '0',
		10885 => '0',
		10886 => '0',
		10887 => '0',
		10888 => '0',
		10889 => '0',
		10890 => '0',
		10891 => '0',
		10892 => '0',
		10893 => '0',
		10894 => '0',
		10895 => '0',
		10896 => '0',
		10897 => '0',
		10898 => '0',
		10899 => '0',
		10900 => '1',
		10901 => '1',
		10902 => '1',
		10903 => '1',
		10904 => '1',
		10905 => '1',
		10906 => '1',
		10907 => '1',
		10908 => '1',
		10909 => '0',
		10910 => '0',
		10911 => '0',
		10912 => '0',
		10913 => '0',
		10914 => '0',
		10915 => '0',
		10916 => '0',
		10917 => '0',
		10918 => '0',
		10919 => '0',
		10920 => '0',
		10921 => '0',
		10922 => '0',
		10923 => '0',
		10924 => '0',
		10925 => '0',
		10926 => '0',
		10927 => '0',
		10928 => '0',
		10929 => '0',
		10930 => '0',
		10931 => '0',
		10932 => '0',
		10933 => '0',
		10934 => '0',
		10935 => '0',
		10936 => '0',
		10937 => '0',
		10938 => '0',
		10939 => '0',
		10940 => '0',
		10941 => '0',
		10942 => '0',
		10943 => '0',
		10944 => '0',
		10945 => '0',
		10946 => '0',
		10947 => '0',
		10948 => '0',
		10949 => '0',
		10950 => '0',
		10951 => '0',
		10952 => '0',
		10953 => '0',
		10954 => '0',
		10955 => '0',
		10956 => '0',
		10957 => '0',
		10958 => '0',
		10959 => '0',
		10960 => '0',
		10961 => '0',
		10962 => '0',
		10963 => '0',
		10964 => '0',
		10965 => '0',
		10966 => '0',
		10967 => '0',
		10968 => '0',
		10969 => '0',
		10970 => '0',
		10971 => '1',
		10972 => '1',
		10973 => '1',
		10974 => '1',
		10975 => '1',
		10976 => '1',
		10977 => '1',
		10978 => '1',
		10979 => '0',
		10980 => '0',
		10981 => '1',
		10982 => '1',
		10983 => '0',
		10984 => '0',
		10985 => '1',
		10986 => '0',
		10987 => '0',
		10988 => '0',
		10989 => '0',
		10990 => '0',
		10991 => '0',
		10992 => '0',
		10993 => '0',
		10994 => '0',
		10995 => '0',
		10996 => '0',
		10997 => '0',
		10998 => '0',
		10999 => '0',
		11008 => '0',
		11009 => '0',
		11010 => '0',
		11011 => '0',
		11012 => '0',
		11013 => '0',
		11014 => '0',
		11015 => '0',
		11016 => '0',
		11017 => '0',
		11018 => '0',
		11019 => '0',
		11020 => '0',
		11021 => '0',
		11022 => '0',
		11023 => '0',
		11024 => '0',
		11025 => '0',
		11026 => '0',
		11027 => '0',
		11028 => '0',
		11029 => '0',
		11030 => '1',
		11031 => '1',
		11032 => '1',
		11033 => '1',
		11034 => '1',
		11035 => '1',
		11036 => '1',
		11037 => '1',
		11038 => '0',
		11039 => '0',
		11040 => '0',
		11041 => '0',
		11042 => '0',
		11043 => '0',
		11044 => '0',
		11045 => '0',
		11046 => '0',
		11047 => '0',
		11048 => '0',
		11049 => '0',
		11050 => '0',
		11051 => '0',
		11052 => '0',
		11053 => '0',
		11054 => '0',
		11055 => '0',
		11056 => '0',
		11057 => '0',
		11058 => '0',
		11059 => '0',
		11060 => '0',
		11061 => '0',
		11062 => '0',
		11063 => '0',
		11064 => '0',
		11065 => '0',
		11066 => '0',
		11067 => '0',
		11068 => '0',
		11069 => '0',
		11070 => '0',
		11071 => '0',
		11072 => '0',
		11073 => '0',
		11074 => '0',
		11075 => '0',
		11076 => '0',
		11077 => '0',
		11078 => '0',
		11079 => '0',
		11080 => '0',
		11081 => '0',
		11082 => '0',
		11083 => '0',
		11084 => '0',
		11085 => '0',
		11086 => '0',
		11087 => '0',
		11088 => '0',
		11089 => '0',
		11090 => '0',
		11091 => '0',
		11092 => '0',
		11093 => '0',
		11094 => '0',
		11095 => '0',
		11096 => '0',
		11097 => '0',
		11098 => '1',
		11099 => '1',
		11100 => '1',
		11101 => '1',
		11102 => '1',
		11103 => '1',
		11104 => '1',
		11105 => '1',
		11106 => '0',
		11107 => '0',
		11108 => '1',
		11109 => '1',
		11110 => '0',
		11111 => '0',
		11112 => '1',
		11113 => '1',
		11114 => '0',
		11115 => '0',
		11116 => '0',
		11117 => '0',
		11118 => '0',
		11119 => '0',
		11120 => '0',
		11121 => '0',
		11122 => '0',
		11123 => '0',
		11124 => '0',
		11125 => '0',
		11126 => '0',
		11127 => '0',
		11136 => '0',
		11137 => '0',
		11138 => '0',
		11139 => '0',
		11140 => '0',
		11141 => '0',
		11142 => '0',
		11143 => '0',
		11144 => '0',
		11145 => '0',
		11146 => '0',
		11147 => '0',
		11148 => '0',
		11149 => '0',
		11150 => '0',
		11151 => '0',
		11152 => '0',
		11153 => '0',
		11154 => '0',
		11155 => '0',
		11156 => '0',
		11157 => '1',
		11158 => '0',
		11159 => '1',
		11160 => '1',
		11161 => '1',
		11162 => '1',
		11163 => '1',
		11164 => '1',
		11165 => '1',
		11166 => '1',
		11167 => '0',
		11168 => '0',
		11169 => '0',
		11170 => '0',
		11171 => '0',
		11172 => '0',
		11173 => '0',
		11174 => '0',
		11175 => '0',
		11176 => '0',
		11177 => '0',
		11178 => '0',
		11179 => '0',
		11180 => '0',
		11181 => '0',
		11182 => '0',
		11183 => '0',
		11184 => '0',
		11185 => '0',
		11186 => '0',
		11187 => '0',
		11188 => '0',
		11189 => '0',
		11190 => '0',
		11191 => '0',
		11192 => '0',
		11193 => '0',
		11194 => '0',
		11195 => '0',
		11196 => '0',
		11197 => '0',
		11198 => '0',
		11199 => '0',
		11200 => '0',
		11201 => '0',
		11202 => '0',
		11203 => '0',
		11204 => '0',
		11205 => '0',
		11206 => '0',
		11207 => '0',
		11208 => '0',
		11209 => '0',
		11210 => '0',
		11211 => '0',
		11212 => '0',
		11213 => '0',
		11214 => '0',
		11215 => '0',
		11216 => '0',
		11217 => '0',
		11218 => '0',
		11219 => '0',
		11220 => '0',
		11221 => '0',
		11222 => '0',
		11223 => '0',
		11224 => '0',
		11225 => '1',
		11226 => '1',
		11227 => '1',
		11228 => '1',
		11229 => '1',
		11230 => '1',
		11231 => '1',
		11232 => '1',
		11233 => '0',
		11234 => '0',
		11235 => '0',
		11236 => '1',
		11237 => '1',
		11238 => '0',
		11239 => '0',
		11240 => '1',
		11241 => '0',
		11242 => '0',
		11243 => '0',
		11244 => '0',
		11245 => '0',
		11246 => '0',
		11247 => '0',
		11248 => '0',
		11249 => '0',
		11250 => '0',
		11251 => '0',
		11252 => '0',
		11253 => '0',
		11254 => '0',
		11255 => '0',
		11264 => '0',
		11265 => '0',
		11266 => '0',
		11267 => '0',
		11268 => '0',
		11269 => '0',
		11270 => '0',
		11271 => '0',
		11272 => '0',
		11273 => '0',
		11274 => '0',
		11275 => '0',
		11276 => '0',
		11277 => '0',
		11278 => '0',
		11279 => '0',
		11280 => '0',
		11281 => '0',
		11282 => '0',
		11283 => '0',
		11284 => '0',
		11285 => '0',
		11286 => '1',
		11287 => '1',
		11288 => '1',
		11289 => '1',
		11290 => '1',
		11291 => '1',
		11292 => '1',
		11293 => '1',
		11294 => '1',
		11295 => '1',
		11296 => '0',
		11297 => '0',
		11298 => '0',
		11299 => '0',
		11300 => '0',
		11301 => '0',
		11302 => '0',
		11303 => '0',
		11304 => '0',
		11305 => '0',
		11306 => '0',
		11307 => '0',
		11308 => '0',
		11309 => '0',
		11310 => '0',
		11311 => '0',
		11312 => '0',
		11313 => '0',
		11314 => '0',
		11315 => '0',
		11316 => '0',
		11317 => '0',
		11318 => '0',
		11319 => '0',
		11320 => '0',
		11321 => '0',
		11322 => '0',
		11323 => '0',
		11324 => '0',
		11325 => '0',
		11326 => '0',
		11327 => '0',
		11328 => '0',
		11329 => '0',
		11330 => '0',
		11331 => '0',
		11332 => '0',
		11333 => '0',
		11334 => '0',
		11335 => '0',
		11336 => '0',
		11337 => '0',
		11338 => '0',
		11339 => '0',
		11340 => '0',
		11341 => '0',
		11342 => '0',
		11343 => '0',
		11344 => '0',
		11345 => '0',
		11346 => '0',
		11347 => '0',
		11348 => '0',
		11349 => '0',
		11350 => '0',
		11351 => '0',
		11352 => '1',
		11353 => '1',
		11354 => '1',
		11355 => '1',
		11356 => '1',
		11357 => '1',
		11358 => '1',
		11359 => '1',
		11360 => '1',
		11361 => '0',
		11362 => '0',
		11363 => '1',
		11364 => '1',
		11365 => '0',
		11366 => '0',
		11367 => '1',
		11368 => '1',
		11369 => '0',
		11370 => '0',
		11371 => '0',
		11372 => '0',
		11373 => '0',
		11374 => '0',
		11375 => '0',
		11376 => '0',
		11377 => '0',
		11378 => '0',
		11379 => '0',
		11380 => '0',
		11381 => '0',
		11382 => '0',
		11383 => '0',
		11392 => '0',
		11393 => '0',
		11394 => '0',
		11395 => '0',
		11396 => '0',
		11397 => '0',
		11398 => '0',
		11399 => '0',
		11400 => '0',
		11401 => '0',
		11402 => '0',
		11403 => '0',
		11404 => '0',
		11405 => '0',
		11406 => '0',
		11407 => '0',
		11408 => '0',
		11409 => '0',
		11410 => '0',
		11411 => '0',
		11412 => '0',
		11413 => '0',
		11414 => '0',
		11415 => '0',
		11416 => '1',
		11417 => '1',
		11418 => '1',
		11419 => '1',
		11420 => '1',
		11421 => '1',
		11422 => '1',
		11423 => '1',
		11424 => '1',
		11425 => '0',
		11426 => '0',
		11427 => '0',
		11428 => '0',
		11429 => '0',
		11430 => '0',
		11431 => '0',
		11432 => '0',
		11433 => '0',
		11434 => '0',
		11435 => '0',
		11436 => '0',
		11437 => '0',
		11438 => '0',
		11439 => '0',
		11440 => '0',
		11441 => '0',
		11442 => '0',
		11443 => '0',
		11444 => '0',
		11445 => '0',
		11446 => '0',
		11447 => '0',
		11448 => '0',
		11449 => '0',
		11450 => '0',
		11451 => '0',
		11452 => '0',
		11453 => '0',
		11454 => '0',
		11455 => '0',
		11456 => '0',
		11457 => '0',
		11458 => '0',
		11459 => '0',
		11460 => '0',
		11461 => '0',
		11462 => '0',
		11463 => '0',
		11464 => '0',
		11465 => '0',
		11466 => '0',
		11467 => '0',
		11468 => '0',
		11469 => '0',
		11470 => '0',
		11471 => '0',
		11472 => '0',
		11473 => '0',
		11474 => '0',
		11475 => '0',
		11476 => '0',
		11477 => '0',
		11478 => '0',
		11479 => '1',
		11480 => '1',
		11481 => '1',
		11482 => '1',
		11483 => '1',
		11484 => '1',
		11485 => '1',
		11486 => '1',
		11487 => '1',
		11488 => '0',
		11489 => '0',
		11490 => '1',
		11491 => '1',
		11492 => '1',
		11493 => '0',
		11494 => '0',
		11495 => '1',
		11496 => '0',
		11497 => '0',
		11498 => '0',
		11499 => '0',
		11500 => '0',
		11501 => '0',
		11502 => '0',
		11503 => '0',
		11504 => '0',
		11505 => '0',
		11506 => '0',
		11507 => '0',
		11508 => '0',
		11509 => '0',
		11510 => '0',
		11511 => '0',
		11520 => '0',
		11521 => '0',
		11522 => '0',
		11523 => '0',
		11524 => '0',
		11525 => '0',
		11526 => '0',
		11527 => '0',
		11528 => '0',
		11529 => '0',
		11530 => '0',
		11531 => '0',
		11532 => '0',
		11533 => '0',
		11534 => '0',
		11535 => '0',
		11536 => '0',
		11537 => '0',
		11538 => '0',
		11539 => '0',
		11540 => '0',
		11541 => '0',
		11542 => '0',
		11543 => '1',
		11544 => '0',
		11545 => '1',
		11546 => '1',
		11547 => '1',
		11548 => '1',
		11549 => '1',
		11550 => '1',
		11551 => '1',
		11552 => '1',
		11553 => '1',
		11554 => '0',
		11555 => '0',
		11556 => '0',
		11557 => '0',
		11558 => '0',
		11559 => '0',
		11560 => '0',
		11561 => '0',
		11562 => '0',
		11563 => '0',
		11564 => '0',
		11565 => '0',
		11566 => '0',
		11567 => '0',
		11568 => '0',
		11569 => '0',
		11570 => '0',
		11571 => '0',
		11572 => '0',
		11573 => '0',
		11574 => '0',
		11575 => '0',
		11576 => '0',
		11577 => '0',
		11578 => '0',
		11579 => '0',
		11580 => '0',
		11581 => '0',
		11582 => '0',
		11583 => '0',
		11584 => '0',
		11585 => '0',
		11586 => '0',
		11587 => '0',
		11588 => '0',
		11589 => '0',
		11590 => '0',
		11591 => '0',
		11592 => '0',
		11593 => '0',
		11594 => '0',
		11595 => '0',
		11596 => '0',
		11597 => '0',
		11598 => '0',
		11599 => '0',
		11600 => '0',
		11601 => '0',
		11602 => '0',
		11603 => '0',
		11604 => '0',
		11605 => '0',
		11606 => '1',
		11607 => '1',
		11608 => '1',
		11609 => '1',
		11610 => '1',
		11611 => '1',
		11612 => '1',
		11613 => '1',
		11614 => '1',
		11615 => '0',
		11616 => '0',
		11617 => '0',
		11618 => '1',
		11619 => '1',
		11620 => '0',
		11621 => '0',
		11622 => '1',
		11623 => '1',
		11624 => '0',
		11625 => '0',
		11626 => '0',
		11627 => '0',
		11628 => '0',
		11629 => '0',
		11630 => '0',
		11631 => '0',
		11632 => '0',
		11633 => '0',
		11634 => '0',
		11635 => '0',
		11636 => '0',
		11637 => '0',
		11638 => '0',
		11639 => '0',
		11648 => '0',
		11649 => '0',
		11650 => '0',
		11651 => '0',
		11652 => '0',
		11653 => '0',
		11654 => '0',
		11655 => '0',
		11656 => '0',
		11657 => '0',
		11658 => '0',
		11659 => '0',
		11660 => '0',
		11661 => '0',
		11662 => '0',
		11663 => '0',
		11664 => '0',
		11665 => '0',
		11666 => '0',
		11667 => '0',
		11668 => '0',
		11669 => '0',
		11670 => '0',
		11671 => '0',
		11672 => '1',
		11673 => '0',
		11674 => '1',
		11675 => '1',
		11676 => '1',
		11677 => '1',
		11678 => '1',
		11679 => '1',
		11680 => '1',
		11681 => '1',
		11682 => '1',
		11683 => '0',
		11684 => '0',
		11685 => '0',
		11686 => '0',
		11687 => '0',
		11688 => '0',
		11689 => '0',
		11690 => '0',
		11691 => '0',
		11692 => '0',
		11693 => '0',
		11694 => '0',
		11695 => '0',
		11696 => '0',
		11697 => '0',
		11698 => '0',
		11699 => '0',
		11700 => '0',
		11701 => '0',
		11702 => '0',
		11703 => '0',
		11704 => '0',
		11705 => '0',
		11706 => '0',
		11707 => '0',
		11708 => '0',
		11709 => '0',
		11710 => '0',
		11711 => '0',
		11712 => '0',
		11713 => '0',
		11714 => '0',
		11715 => '0',
		11716 => '0',
		11717 => '0',
		11718 => '0',
		11719 => '0',
		11720 => '0',
		11721 => '0',
		11722 => '0',
		11723 => '0',
		11724 => '0',
		11725 => '0',
		11726 => '0',
		11727 => '0',
		11728 => '0',
		11729 => '0',
		11730 => '0',
		11731 => '0',
		11732 => '0',
		11733 => '1',
		11734 => '1',
		11735 => '1',
		11736 => '1',
		11737 => '1',
		11738 => '1',
		11739 => '1',
		11740 => '1',
		11741 => '1',
		11742 => '0',
		11743 => '0',
		11744 => '0',
		11745 => '1',
		11746 => '1',
		11747 => '0',
		11748 => '0',
		11749 => '0',
		11750 => '1',
		11751 => '0',
		11752 => '0',
		11753 => '0',
		11754 => '0',
		11755 => '0',
		11756 => '0',
		11757 => '0',
		11758 => '0',
		11759 => '0',
		11760 => '0',
		11761 => '0',
		11762 => '0',
		11763 => '0',
		11764 => '0',
		11765 => '0',
		11766 => '0',
		11767 => '0',
		11776 => '0',
		11777 => '0',
		11778 => '0',
		11779 => '0',
		11780 => '0',
		11781 => '0',
		11782 => '0',
		11783 => '0',
		11784 => '0',
		11785 => '0',
		11786 => '0',
		11787 => '0',
		11788 => '0',
		11789 => '0',
		11790 => '0',
		11791 => '0',
		11792 => '0',
		11793 => '0',
		11794 => '0',
		11795 => '0',
		11796 => '0',
		11797 => '0',
		11798 => '0',
		11799 => '0',
		11800 => '0',
		11801 => '1',
		11802 => '0',
		11803 => '1',
		11804 => '1',
		11805 => '1',
		11806 => '1',
		11807 => '1',
		11808 => '1',
		11809 => '1',
		11810 => '1',
		11811 => '1',
		11812 => '1',
		11813 => '0',
		11814 => '0',
		11815 => '0',
		11816 => '0',
		11817 => '0',
		11818 => '0',
		11819 => '0',
		11820 => '0',
		11821 => '0',
		11822 => '0',
		11823 => '0',
		11824 => '0',
		11825 => '0',
		11826 => '0',
		11827 => '0',
		11828 => '0',
		11829 => '0',
		11830 => '0',
		11831 => '0',
		11832 => '0',
		11833 => '0',
		11834 => '0',
		11835 => '0',
		11836 => '0',
		11837 => '0',
		11838 => '0',
		11839 => '0',
		11840 => '0',
		11841 => '0',
		11842 => '0',
		11843 => '0',
		11844 => '0',
		11845 => '0',
		11846 => '0',
		11847 => '0',
		11848 => '0',
		11849 => '0',
		11850 => '0',
		11851 => '0',
		11852 => '0',
		11853 => '0',
		11854 => '0',
		11855 => '0',
		11856 => '0',
		11857 => '0',
		11858 => '0',
		11859 => '1',
		11860 => '1',
		11861 => '1',
		11862 => '1',
		11863 => '1',
		11864 => '1',
		11865 => '1',
		11866 => '1',
		11867 => '1',
		11868 => '1',
		11869 => '0',
		11870 => '0',
		11871 => '0',
		11872 => '1',
		11873 => '1',
		11874 => '1',
		11875 => '0',
		11876 => '0',
		11877 => '1',
		11878 => '1',
		11879 => '0',
		11880 => '0',
		11881 => '0',
		11882 => '0',
		11883 => '0',
		11884 => '0',
		11885 => '0',
		11886 => '0',
		11887 => '0',
		11888 => '0',
		11889 => '0',
		11890 => '0',
		11891 => '0',
		11892 => '0',
		11893 => '0',
		11894 => '0',
		11895 => '0',
		11904 => '0',
		11905 => '0',
		11906 => '0',
		11907 => '0',
		11908 => '0',
		11909 => '0',
		11910 => '0',
		11911 => '0',
		11912 => '0',
		11913 => '0',
		11914 => '0',
		11915 => '0',
		11916 => '0',
		11917 => '0',
		11918 => '0',
		11919 => '0',
		11920 => '0',
		11921 => '0',
		11922 => '0',
		11923 => '0',
		11924 => '0',
		11925 => '0',
		11926 => '0',
		11927 => '0',
		11928 => '0',
		11929 => '0',
		11930 => '1',
		11931 => '0',
		11932 => '1',
		11933 => '1',
		11934 => '1',
		11935 => '1',
		11936 => '1',
		11937 => '1',
		11938 => '1',
		11939 => '1',
		11940 => '1',
		11941 => '1',
		11942 => '0',
		11943 => '0',
		11944 => '0',
		11945 => '0',
		11946 => '0',
		11947 => '0',
		11948 => '0',
		11949 => '0',
		11950 => '0',
		11951 => '0',
		11952 => '0',
		11953 => '0',
		11954 => '0',
		11955 => '0',
		11956 => '0',
		11957 => '0',
		11958 => '0',
		11959 => '0',
		11960 => '0',
		11961 => '0',
		11962 => '0',
		11963 => '0',
		11964 => '0',
		11965 => '0',
		11966 => '0',
		11967 => '0',
		11968 => '0',
		11969 => '0',
		11970 => '0',
		11971 => '0',
		11972 => '0',
		11973 => '0',
		11974 => '0',
		11975 => '0',
		11976 => '0',
		11977 => '0',
		11978 => '0',
		11979 => '0',
		11980 => '0',
		11981 => '0',
		11982 => '0',
		11983 => '0',
		11984 => '0',
		11985 => '0',
		11986 => '1',
		11987 => '1',
		11988 => '1',
		11989 => '1',
		11990 => '1',
		11991 => '1',
		11992 => '1',
		11993 => '1',
		11994 => '1',
		11995 => '1',
		11996 => '0',
		11997 => '0',
		11998 => '0',
		11999 => '1',
		12000 => '1',
		12001 => '1',
		12002 => '0',
		12003 => '0',
		12004 => '1',
		12005 => '1',
		12006 => '0',
		12007 => '0',
		12008 => '0',
		12009 => '0',
		12010 => '0',
		12011 => '0',
		12012 => '0',
		12013 => '0',
		12014 => '0',
		12015 => '0',
		12016 => '0',
		12017 => '0',
		12018 => '0',
		12019 => '0',
		12020 => '0',
		12021 => '0',
		12022 => '0',
		12023 => '0',
		12032 => '0',
		12033 => '0',
		12034 => '0',
		12035 => '0',
		12036 => '0',
		12037 => '0',
		12038 => '0',
		12039 => '0',
		12040 => '0',
		12041 => '0',
		12042 => '0',
		12043 => '0',
		12044 => '0',
		12045 => '0',
		12046 => '0',
		12047 => '0',
		12048 => '0',
		12049 => '0',
		12050 => '0',
		12051 => '0',
		12052 => '0',
		12053 => '0',
		12054 => '0',
		12055 => '0',
		12056 => '0',
		12057 => '0',
		12058 => '0',
		12059 => '1',
		12060 => '0',
		12061 => '1',
		12062 => '1',
		12063 => '1',
		12064 => '1',
		12065 => '1',
		12066 => '1',
		12067 => '1',
		12068 => '1',
		12069 => '1',
		12070 => '1',
		12071 => '1',
		12072 => '0',
		12073 => '0',
		12074 => '0',
		12075 => '0',
		12076 => '0',
		12077 => '0',
		12078 => '0',
		12079 => '0',
		12080 => '0',
		12081 => '0',
		12082 => '0',
		12083 => '0',
		12084 => '0',
		12085 => '0',
		12086 => '0',
		12087 => '0',
		12088 => '0',
		12089 => '0',
		12090 => '0',
		12091 => '0',
		12092 => '0',
		12093 => '0',
		12094 => '0',
		12095 => '0',
		12096 => '0',
		12097 => '0',
		12098 => '0',
		12099 => '0',
		12100 => '0',
		12101 => '0',
		12102 => '0',
		12103 => '0',
		12104 => '0',
		12105 => '0',
		12106 => '0',
		12107 => '0',
		12108 => '0',
		12109 => '0',
		12110 => '0',
		12111 => '0',
		12112 => '1',
		12113 => '1',
		12114 => '1',
		12115 => '1',
		12116 => '1',
		12117 => '1',
		12118 => '1',
		12119 => '1',
		12120 => '1',
		12121 => '1',
		12122 => '1',
		12123 => '0',
		12124 => '0',
		12125 => '0',
		12126 => '1',
		12127 => '1',
		12128 => '1',
		12129 => '0',
		12130 => '0',
		12131 => '0',
		12132 => '1',
		12133 => '0',
		12134 => '0',
		12135 => '0',
		12136 => '0',
		12137 => '0',
		12138 => '0',
		12139 => '0',
		12140 => '0',
		12141 => '0',
		12142 => '0',
		12143 => '0',
		12144 => '0',
		12145 => '0',
		12146 => '0',
		12147 => '0',
		12148 => '0',
		12149 => '0',
		12150 => '0',
		12151 => '0',
		12160 => '0',
		12161 => '0',
		12162 => '0',
		12163 => '0',
		12164 => '0',
		12165 => '0',
		12166 => '0',
		12167 => '0',
		12168 => '0',
		12169 => '0',
		12170 => '0',
		12171 => '0',
		12172 => '0',
		12173 => '0',
		12174 => '0',
		12175 => '0',
		12176 => '0',
		12177 => '0',
		12178 => '0',
		12179 => '0',
		12180 => '0',
		12181 => '0',
		12182 => '0',
		12183 => '0',
		12184 => '0',
		12185 => '0',
		12186 => '0',
		12187 => '0',
		12188 => '1',
		12189 => '0',
		12190 => '1',
		12191 => '1',
		12192 => '1',
		12193 => '1',
		12194 => '1',
		12195 => '1',
		12196 => '1',
		12197 => '1',
		12198 => '1',
		12199 => '1',
		12200 => '1',
		12201 => '1',
		12202 => '0',
		12203 => '0',
		12204 => '0',
		12205 => '0',
		12206 => '0',
		12207 => '0',
		12208 => '0',
		12209 => '0',
		12210 => '0',
		12211 => '0',
		12212 => '0',
		12213 => '0',
		12214 => '0',
		12215 => '0',
		12216 => '0',
		12217 => '0',
		12218 => '0',
		12219 => '0',
		12220 => '0',
		12221 => '0',
		12222 => '0',
		12223 => '0',
		12224 => '0',
		12225 => '0',
		12226 => '0',
		12227 => '0',
		12228 => '0',
		12229 => '0',
		12230 => '0',
		12231 => '0',
		12232 => '0',
		12233 => '0',
		12234 => '0',
		12235 => '0',
		12236 => '0',
		12237 => '0',
		12238 => '1',
		12239 => '1',
		12240 => '1',
		12241 => '1',
		12242 => '1',
		12243 => '1',
		12244 => '1',
		12245 => '1',
		12246 => '1',
		12247 => '1',
		12248 => '1',
		12249 => '1',
		12250 => '0',
		12251 => '0',
		12252 => '0',
		12253 => '1',
		12254 => '1',
		12255 => '1',
		12256 => '0',
		12257 => '0',
		12258 => '0',
		12259 => '1',
		12260 => '1',
		12261 => '0',
		12262 => '0',
		12263 => '0',
		12264 => '0',
		12265 => '0',
		12266 => '0',
		12267 => '0',
		12268 => '0',
		12269 => '0',
		12270 => '0',
		12271 => '0',
		12272 => '0',
		12273 => '0',
		12274 => '0',
		12275 => '0',
		12276 => '0',
		12277 => '0',
		12278 => '0',
		12279 => '0',
		12288 => '0',
		12289 => '0',
		12290 => '0',
		12291 => '0',
		12292 => '0',
		12293 => '0',
		12294 => '0',
		12295 => '0',
		12296 => '0',
		12297 => '0',
		12298 => '0',
		12299 => '0',
		12300 => '0',
		12301 => '0',
		12302 => '0',
		12303 => '0',
		12304 => '0',
		12305 => '0',
		12306 => '0',
		12307 => '0',
		12308 => '0',
		12309 => '0',
		12310 => '0',
		12311 => '0',
		12312 => '0',
		12313 => '0',
		12314 => '0',
		12315 => '0',
		12316 => '0',
		12317 => '1',
		12318 => '0',
		12319 => '1',
		12320 => '1',
		12321 => '1',
		12322 => '1',
		12323 => '1',
		12324 => '1',
		12325 => '1',
		12326 => '1',
		12327 => '1',
		12328 => '1',
		12329 => '1',
		12330 => '1',
		12331 => '1',
		12332 => '0',
		12333 => '0',
		12334 => '0',
		12335 => '0',
		12336 => '0',
		12337 => '0',
		12338 => '0',
		12339 => '0',
		12340 => '0',
		12341 => '0',
		12342 => '0',
		12343 => '0',
		12344 => '0',
		12345 => '0',
		12346 => '0',
		12347 => '0',
		12348 => '0',
		12349 => '0',
		12350 => '0',
		12351 => '0',
		12352 => '0',
		12353 => '0',
		12354 => '0',
		12355 => '0',
		12356 => '0',
		12357 => '0',
		12358 => '0',
		12359 => '0',
		12360 => '0',
		12361 => '0',
		12362 => '0',
		12363 => '0',
		12364 => '1',
		12365 => '1',
		12366 => '1',
		12367 => '1',
		12368 => '1',
		12369 => '1',
		12370 => '1',
		12371 => '1',
		12372 => '1',
		12373 => '1',
		12374 => '1',
		12375 => '1',
		12376 => '1',
		12377 => '0',
		12378 => '0',
		12379 => '0',
		12380 => '1',
		12381 => '1',
		12382 => '1',
		12383 => '0',
		12384 => '0',
		12385 => '0',
		12386 => '1',
		12387 => '1',
		12388 => '0',
		12389 => '0',
		12390 => '0',
		12391 => '0',
		12392 => '0',
		12393 => '0',
		12394 => '0',
		12395 => '0',
		12396 => '0',
		12397 => '0',
		12398 => '0',
		12399 => '0',
		12400 => '0',
		12401 => '0',
		12402 => '0',
		12403 => '0',
		12404 => '0',
		12405 => '0',
		12406 => '0',
		12407 => '0',
		12416 => '0',
		12417 => '0',
		12418 => '0',
		12419 => '0',
		12420 => '0',
		12421 => '0',
		12422 => '0',
		12423 => '0',
		12424 => '0',
		12425 => '0',
		12426 => '0',
		12427 => '0',
		12428 => '0',
		12429 => '0',
		12430 => '0',
		12431 => '0',
		12432 => '0',
		12433 => '0',
		12434 => '0',
		12435 => '0',
		12436 => '0',
		12437 => '0',
		12438 => '0',
		12439 => '0',
		12440 => '0',
		12441 => '0',
		12442 => '0',
		12443 => '0',
		12444 => '0',
		12445 => '0',
		12446 => '1',
		12447 => '0',
		12448 => '0',
		12449 => '1',
		12450 => '1',
		12451 => '1',
		12452 => '1',
		12453 => '1',
		12454 => '1',
		12455 => '1',
		12456 => '1',
		12457 => '1',
		12458 => '1',
		12459 => '1',
		12460 => '1',
		12461 => '1',
		12462 => '0',
		12463 => '0',
		12464 => '0',
		12465 => '0',
		12466 => '0',
		12467 => '0',
		12468 => '0',
		12469 => '0',
		12470 => '0',
		12471 => '0',
		12472 => '0',
		12473 => '0',
		12474 => '0',
		12475 => '0',
		12476 => '0',
		12477 => '0',
		12478 => '0',
		12479 => '0',
		12480 => '0',
		12481 => '0',
		12482 => '0',
		12483 => '0',
		12484 => '0',
		12485 => '0',
		12486 => '0',
		12487 => '0',
		12488 => '0',
		12489 => '0',
		12490 => '1',
		12491 => '1',
		12492 => '1',
		12493 => '1',
		12494 => '1',
		12495 => '1',
		12496 => '1',
		12497 => '1',
		12498 => '1',
		12499 => '1',
		12500 => '1',
		12501 => '1',
		12502 => '1',
		12503 => '0',
		12504 => '0',
		12505 => '0',
		12506 => '0',
		12507 => '1',
		12508 => '1',
		12509 => '1',
		12510 => '0',
		12511 => '0',
		12512 => '0',
		12513 => '1',
		12514 => '1',
		12515 => '0',
		12516 => '0',
		12517 => '0',
		12518 => '0',
		12519 => '0',
		12520 => '0',
		12521 => '0',
		12522 => '0',
		12523 => '0',
		12524 => '0',
		12525 => '0',
		12526 => '0',
		12527 => '0',
		12528 => '0',
		12529 => '0',
		12530 => '0',
		12531 => '0',
		12532 => '0',
		12533 => '0',
		12534 => '0',
		12535 => '0',
		12544 => '0',
		12545 => '0',
		12546 => '0',
		12547 => '0',
		12548 => '0',
		12549 => '0',
		12550 => '0',
		12551 => '0',
		12552 => '0',
		12553 => '0',
		12554 => '0',
		12555 => '0',
		12556 => '0',
		12557 => '0',
		12558 => '0',
		12559 => '0',
		12560 => '0',
		12561 => '0',
		12562 => '0',
		12563 => '0',
		12564 => '0',
		12565 => '0',
		12566 => '0',
		12567 => '0',
		12568 => '0',
		12569 => '0',
		12570 => '0',
		12571 => '0',
		12572 => '0',
		12573 => '0',
		12574 => '0',
		12575 => '1',
		12576 => '0',
		12577 => '0',
		12578 => '1',
		12579 => '1',
		12580 => '1',
		12581 => '1',
		12582 => '1',
		12583 => '1',
		12584 => '1',
		12585 => '1',
		12586 => '1',
		12587 => '1',
		12588 => '1',
		12589 => '1',
		12590 => '1',
		12591 => '1',
		12592 => '1',
		12593 => '0',
		12594 => '0',
		12595 => '0',
		12596 => '0',
		12597 => '0',
		12598 => '0',
		12599 => '0',
		12600 => '0',
		12601 => '0',
		12602 => '0',
		12603 => '0',
		12604 => '0',
		12605 => '0',
		12606 => '0',
		12607 => '0',
		12608 => '0',
		12609 => '0',
		12610 => '0',
		12611 => '0',
		12612 => '0',
		12613 => '0',
		12614 => '0',
		12615 => '1',
		12616 => '1',
		12617 => '1',
		12618 => '1',
		12619 => '1',
		12620 => '1',
		12621 => '1',
		12622 => '1',
		12623 => '1',
		12624 => '1',
		12625 => '1',
		12626 => '1',
		12627 => '1',
		12628 => '1',
		12629 => '1',
		12630 => '0',
		12631 => '0',
		12632 => '0',
		12633 => '0',
		12634 => '1',
		12635 => '1',
		12636 => '1',
		12637 => '0',
		12638 => '0',
		12639 => '0',
		12640 => '1',
		12641 => '1',
		12642 => '0',
		12643 => '0',
		12644 => '0',
		12645 => '0',
		12646 => '0',
		12647 => '0',
		12648 => '0',
		12649 => '0',
		12650 => '0',
		12651 => '0',
		12652 => '0',
		12653 => '0',
		12654 => '0',
		12655 => '0',
		12656 => '0',
		12657 => '0',
		12658 => '0',
		12659 => '0',
		12660 => '0',
		12661 => '0',
		12662 => '0',
		12663 => '0',
		12672 => '0',
		12673 => '0',
		12674 => '0',
		12675 => '0',
		12676 => '0',
		12677 => '0',
		12678 => '0',
		12679 => '0',
		12680 => '0',
		12681 => '0',
		12682 => '0',
		12683 => '0',
		12684 => '0',
		12685 => '0',
		12686 => '0',
		12687 => '0',
		12688 => '0',
		12689 => '0',
		12690 => '0',
		12691 => '0',
		12692 => '0',
		12693 => '0',
		12694 => '0',
		12695 => '0',
		12696 => '0',
		12697 => '0',
		12698 => '0',
		12699 => '0',
		12700 => '0',
		12701 => '0',
		12702 => '0',
		12703 => '0',
		12704 => '1',
		12705 => '1',
		12706 => '0',
		12707 => '0',
		12708 => '1',
		12709 => '1',
		12710 => '1',
		12711 => '1',
		12712 => '1',
		12713 => '1',
		12714 => '1',
		12715 => '1',
		12716 => '1',
		12717 => '1',
		12718 => '1',
		12719 => '1',
		12720 => '1',
		12721 => '1',
		12722 => '1',
		12723 => '1',
		12724 => '1',
		12725 => '1',
		12726 => '0',
		12727 => '0',
		12728 => '0',
		12729 => '0',
		12730 => '0',
		12731 => '0',
		12732 => '0',
		12733 => '0',
		12734 => '0',
		12735 => '0',
		12736 => '0',
		12737 => '0',
		12738 => '1',
		12739 => '1',
		12740 => '1',
		12741 => '1',
		12742 => '1',
		12743 => '1',
		12744 => '1',
		12745 => '1',
		12746 => '1',
		12747 => '1',
		12748 => '1',
		12749 => '1',
		12750 => '1',
		12751 => '1',
		12752 => '1',
		12753 => '1',
		12754 => '1',
		12755 => '1',
		12756 => '0',
		12757 => '0',
		12758 => '0',
		12759 => '0',
		12760 => '1',
		12761 => '1',
		12762 => '1',
		12763 => '1',
		12764 => '0',
		12765 => '0',
		12766 => '0',
		12767 => '1',
		12768 => '1',
		12769 => '0',
		12770 => '0',
		12771 => '0',
		12772 => '0',
		12773 => '0',
		12774 => '0',
		12775 => '0',
		12776 => '0',
		12777 => '0',
		12778 => '0',
		12779 => '0',
		12780 => '0',
		12781 => '0',
		12782 => '0',
		12783 => '0',
		12784 => '0',
		12785 => '0',
		12786 => '0',
		12787 => '0',
		12788 => '0',
		12789 => '0',
		12790 => '0',
		12791 => '0',
		12800 => '0',
		12801 => '0',
		12802 => '0',
		12803 => '0',
		12804 => '0',
		12805 => '0',
		12806 => '0',
		12807 => '0',
		12808 => '0',
		12809 => '0',
		12810 => '0',
		12811 => '0',
		12812 => '0',
		12813 => '0',
		12814 => '0',
		12815 => '0',
		12816 => '0',
		12817 => '0',
		12818 => '0',
		12819 => '0',
		12820 => '0',
		12821 => '0',
		12822 => '0',
		12823 => '0',
		12824 => '0',
		12825 => '0',
		12826 => '0',
		12827 => '0',
		12828 => '0',
		12829 => '0',
		12830 => '0',
		12831 => '0',
		12832 => '0',
		12833 => '1',
		12834 => '1',
		12835 => '0',
		12836 => '0',
		12837 => '0',
		12838 => '1',
		12839 => '1',
		12840 => '1',
		12841 => '1',
		12842 => '1',
		12843 => '1',
		12844 => '1',
		12845 => '1',
		12846 => '1',
		12847 => '1',
		12848 => '1',
		12849 => '1',
		12850 => '1',
		12851 => '1',
		12852 => '1',
		12853 => '1',
		12854 => '1',
		12855 => '1',
		12856 => '1',
		12857 => '1',
		12858 => '1',
		12859 => '1',
		12860 => '1',
		12861 => '1',
		12862 => '1',
		12863 => '1',
		12864 => '1',
		12865 => '1',
		12866 => '1',
		12867 => '1',
		12868 => '1',
		12869 => '1',
		12870 => '1',
		12871 => '1',
		12872 => '1',
		12873 => '1',
		12874 => '1',
		12875 => '1',
		12876 => '1',
		12877 => '1',
		12878 => '1',
		12879 => '1',
		12880 => '1',
		12881 => '1',
		12882 => '0',
		12883 => '0',
		12884 => '0',
		12885 => '0',
		12886 => '0',
		12887 => '1',
		12888 => '1',
		12889 => '1',
		12890 => '1',
		12891 => '0',
		12892 => '0',
		12893 => '0',
		12894 => '1',
		12895 => '1',
		12896 => '0',
		12897 => '0',
		12898 => '0',
		12899 => '0',
		12900 => '0',
		12901 => '0',
		12902 => '0',
		12903 => '0',
		12904 => '0',
		12905 => '0',
		12906 => '0',
		12907 => '0',
		12908 => '0',
		12909 => '0',
		12910 => '0',
		12911 => '0',
		12912 => '0',
		12913 => '0',
		12914 => '0',
		12915 => '0',
		12916 => '0',
		12917 => '0',
		12918 => '0',
		12919 => '0',
		12928 => '0',
		12929 => '0',
		12930 => '0',
		12931 => '0',
		12932 => '0',
		12933 => '0',
		12934 => '0',
		12935 => '0',
		12936 => '0',
		12937 => '0',
		12938 => '0',
		12939 => '0',
		12940 => '0',
		12941 => '0',
		12942 => '0',
		12943 => '0',
		12944 => '0',
		12945 => '0',
		12946 => '0',
		12947 => '0',
		12948 => '0',
		12949 => '0',
		12950 => '0',
		12951 => '0',
		12952 => '0',
		12953 => '0',
		12954 => '0',
		12955 => '0',
		12956 => '0',
		12957 => '0',
		12958 => '0',
		12959 => '0',
		12960 => '0',
		12961 => '0',
		12962 => '0',
		12963 => '1',
		12964 => '1',
		12965 => '0',
		12966 => '0',
		12967 => '0',
		12968 => '1',
		12969 => '1',
		12970 => '1',
		12971 => '1',
		12972 => '1',
		12973 => '1',
		12974 => '1',
		12975 => '1',
		12976 => '1',
		12977 => '1',
		12978 => '1',
		12979 => '1',
		12980 => '1',
		12981 => '1',
		12982 => '1',
		12983 => '1',
		12984 => '1',
		12985 => '1',
		12986 => '1',
		12987 => '1',
		12988 => '1',
		12989 => '1',
		12990 => '1',
		12991 => '1',
		12992 => '1',
		12993 => '1',
		12994 => '1',
		12995 => '1',
		12996 => '1',
		12997 => '1',
		12998 => '1',
		12999 => '1',
		13000 => '1',
		13001 => '1',
		13002 => '1',
		13003 => '1',
		13004 => '1',
		13005 => '1',
		13006 => '1',
		13007 => '1',
		13008 => '0',
		13009 => '0',
		13010 => '0',
		13011 => '0',
		13012 => '0',
		13013 => '1',
		13014 => '1',
		13015 => '1',
		13016 => '1',
		13017 => '0',
		13018 => '0',
		13019 => '0',
		13020 => '0',
		13021 => '1',
		13022 => '1',
		13023 => '0',
		13024 => '0',
		13025 => '0',
		13026 => '0',
		13027 => '0',
		13028 => '0',
		13029 => '0',
		13030 => '0',
		13031 => '0',
		13032 => '0',
		13033 => '0',
		13034 => '0',
		13035 => '0',
		13036 => '0',
		13037 => '0',
		13038 => '0',
		13039 => '0',
		13040 => '0',
		13041 => '0',
		13042 => '0',
		13043 => '0',
		13044 => '0',
		13045 => '0',
		13046 => '0',
		13047 => '0',
		13056 => '0',
		13057 => '0',
		13058 => '0',
		13059 => '0',
		13060 => '0',
		13061 => '0',
		13062 => '0',
		13063 => '0',
		13064 => '0',
		13065 => '0',
		13066 => '0',
		13067 => '0',
		13068 => '0',
		13069 => '0',
		13070 => '0',
		13071 => '0',
		13072 => '0',
		13073 => '0',
		13074 => '0',
		13075 => '0',
		13076 => '0',
		13077 => '0',
		13078 => '0',
		13079 => '0',
		13080 => '0',
		13081 => '0',
		13082 => '0',
		13083 => '0',
		13084 => '0',
		13085 => '0',
		13086 => '0',
		13087 => '0',
		13088 => '0',
		13089 => '0',
		13090 => '0',
		13091 => '0',
		13092 => '1',
		13093 => '1',
		13094 => '1',
		13095 => '0',
		13096 => '0',
		13097 => '0',
		13098 => '1',
		13099 => '1',
		13100 => '1',
		13101 => '1',
		13102 => '1',
		13103 => '1',
		13104 => '1',
		13105 => '1',
		13106 => '1',
		13107 => '1',
		13108 => '1',
		13109 => '1',
		13110 => '1',
		13111 => '1',
		13112 => '1',
		13113 => '1',
		13114 => '1',
		13115 => '1',
		13116 => '1',
		13117 => '1',
		13118 => '1',
		13119 => '1',
		13120 => '1',
		13121 => '1',
		13122 => '1',
		13123 => '1',
		13124 => '1',
		13125 => '1',
		13126 => '1',
		13127 => '1',
		13128 => '1',
		13129 => '1',
		13130 => '1',
		13131 => '1',
		13132 => '1',
		13133 => '1',
		13134 => '0',
		13135 => '0',
		13136 => '0',
		13137 => '0',
		13138 => '0',
		13139 => '1',
		13140 => '1',
		13141 => '1',
		13142 => '1',
		13143 => '1',
		13144 => '0',
		13145 => '0',
		13146 => '0',
		13147 => '0',
		13148 => '1',
		13149 => '1',
		13150 => '0',
		13151 => '0',
		13152 => '0',
		13153 => '0',
		13154 => '0',
		13155 => '0',
		13156 => '0',
		13157 => '0',
		13158 => '0',
		13159 => '0',
		13160 => '0',
		13161 => '0',
		13162 => '0',
		13163 => '0',
		13164 => '0',
		13165 => '0',
		13166 => '0',
		13167 => '0',
		13168 => '0',
		13169 => '0',
		13170 => '0',
		13171 => '0',
		13172 => '0',
		13173 => '0',
		13174 => '0',
		13175 => '0',
		13184 => '0',
		13185 => '0',
		13186 => '0',
		13187 => '0',
		13188 => '0',
		13189 => '0',
		13190 => '0',
		13191 => '0',
		13192 => '0',
		13193 => '0',
		13194 => '0',
		13195 => '0',
		13196 => '0',
		13197 => '0',
		13198 => '0',
		13199 => '0',
		13200 => '0',
		13201 => '0',
		13202 => '0',
		13203 => '0',
		13204 => '0',
		13205 => '0',
		13206 => '0',
		13207 => '0',
		13208 => '0',
		13209 => '0',
		13210 => '0',
		13211 => '0',
		13212 => '0',
		13213 => '0',
		13214 => '0',
		13215 => '0',
		13216 => '0',
		13217 => '0',
		13218 => '0',
		13219 => '1',
		13220 => '0',
		13221 => '0',
		13222 => '1',
		13223 => '1',
		13224 => '1',
		13225 => '0',
		13226 => '0',
		13227 => '0',
		13228 => '1',
		13229 => '1',
		13230 => '1',
		13231 => '1',
		13232 => '1',
		13233 => '1',
		13234 => '1',
		13235 => '1',
		13236 => '1',
		13237 => '1',
		13238 => '1',
		13239 => '1',
		13240 => '1',
		13241 => '1',
		13242 => '1',
		13243 => '1',
		13244 => '1',
		13245 => '1',
		13246 => '1',
		13247 => '1',
		13248 => '1',
		13249 => '1',
		13250 => '1',
		13251 => '1',
		13252 => '1',
		13253 => '1',
		13254 => '1',
		13255 => '1',
		13256 => '1',
		13257 => '1',
		13258 => '1',
		13259 => '1',
		13260 => '0',
		13261 => '0',
		13262 => '0',
		13263 => '0',
		13264 => '0',
		13265 => '1',
		13266 => '1',
		13267 => '1',
		13268 => '1',
		13269 => '1',
		13270 => '0',
		13271 => '0',
		13272 => '0',
		13273 => '0',
		13274 => '1',
		13275 => '1',
		13276 => '1',
		13277 => '0',
		13278 => '0',
		13279 => '0',
		13280 => '0',
		13281 => '0',
		13282 => '0',
		13283 => '0',
		13284 => '0',
		13285 => '0',
		13286 => '0',
		13287 => '0',
		13288 => '0',
		13289 => '0',
		13290 => '0',
		13291 => '0',
		13292 => '0',
		13293 => '0',
		13294 => '0',
		13295 => '0',
		13296 => '0',
		13297 => '0',
		13298 => '0',
		13299 => '0',
		13300 => '0',
		13301 => '0',
		13302 => '0',
		13303 => '0',
		13312 => '0',
		13313 => '0',
		13314 => '0',
		13315 => '0',
		13316 => '0',
		13317 => '0',
		13318 => '0',
		13319 => '0',
		13320 => '0',
		13321 => '0',
		13322 => '0',
		13323 => '0',
		13324 => '0',
		13325 => '0',
		13326 => '0',
		13327 => '0',
		13328 => '0',
		13329 => '0',
		13330 => '0',
		13331 => '0',
		13332 => '0',
		13333 => '0',
		13334 => '0',
		13335 => '0',
		13336 => '0',
		13337 => '0',
		13338 => '0',
		13339 => '0',
		13340 => '0',
		13341 => '0',
		13342 => '0',
		13343 => '0',
		13344 => '0',
		13345 => '0',
		13346 => '0',
		13347 => '0',
		13348 => '0',
		13349 => '0',
		13350 => '0',
		13351 => '0',
		13352 => '1',
		13353 => '1',
		13354 => '1',
		13355 => '0',
		13356 => '0',
		13357 => '0',
		13358 => '0',
		13359 => '1',
		13360 => '1',
		13361 => '1',
		13362 => '1',
		13363 => '1',
		13364 => '1',
		13365 => '1',
		13366 => '1',
		13367 => '1',
		13368 => '1',
		13369 => '1',
		13370 => '1',
		13371 => '1',
		13372 => '1',
		13373 => '1',
		13374 => '1',
		13375 => '1',
		13376 => '1',
		13377 => '1',
		13378 => '1',
		13379 => '1',
		13380 => '1',
		13381 => '1',
		13382 => '1',
		13383 => '1',
		13384 => '1',
		13385 => '0',
		13386 => '0',
		13387 => '0',
		13388 => '0',
		13389 => '0',
		13390 => '0',
		13391 => '1',
		13392 => '1',
		13393 => '1',
		13394 => '1',
		13395 => '1',
		13396 => '0',
		13397 => '0',
		13398 => '0',
		13399 => '0',
		13400 => '0',
		13401 => '1',
		13402 => '1',
		13403 => '0',
		13404 => '0',
		13405 => '0',
		13406 => '0',
		13407 => '0',
		13408 => '0',
		13409 => '0',
		13410 => '0',
		13411 => '0',
		13412 => '0',
		13413 => '0',
		13414 => '0',
		13415 => '0',
		13416 => '0',
		13417 => '0',
		13418 => '0',
		13419 => '0',
		13420 => '0',
		13421 => '0',
		13422 => '0',
		13423 => '0',
		13424 => '0',
		13425 => '0',
		13426 => '0',
		13427 => '0',
		13428 => '0',
		13429 => '0',
		13430 => '0',
		13431 => '0',
		13440 => '0',
		13441 => '0',
		13442 => '0',
		13443 => '0',
		13444 => '0',
		13445 => '0',
		13446 => '0',
		13447 => '0',
		13448 => '0',
		13449 => '0',
		13450 => '0',
		13451 => '0',
		13452 => '0',
		13453 => '0',
		13454 => '0',
		13455 => '0',
		13456 => '0',
		13457 => '0',
		13458 => '0',
		13459 => '0',
		13460 => '0',
		13461 => '0',
		13462 => '0',
		13463 => '0',
		13464 => '0',
		13465 => '0',
		13466 => '0',
		13467 => '0',
		13468 => '0',
		13469 => '0',
		13470 => '0',
		13471 => '0',
		13472 => '0',
		13473 => '0',
		13474 => '0',
		13475 => '0',
		13476 => '0',
		13477 => '0',
		13478 => '1',
		13479 => '0',
		13480 => '0',
		13481 => '0',
		13482 => '1',
		13483 => '1',
		13484 => '1',
		13485 => '0',
		13486 => '0',
		13487 => '0',
		13488 => '0',
		13489 => '0',
		13490 => '0',
		13491 => '0',
		13492 => '1',
		13493 => '1',
		13494 => '1',
		13495 => '1',
		13496 => '1',
		13497 => '1',
		13498 => '1',
		13499 => '1',
		13500 => '1',
		13501 => '1',
		13502 => '1',
		13503 => '1',
		13504 => '1',
		13505 => '1',
		13506 => '1',
		13507 => '1',
		13508 => '0',
		13509 => '0',
		13510 => '0',
		13511 => '0',
		13512 => '0',
		13513 => '0',
		13514 => '0',
		13515 => '0',
		13516 => '0',
		13517 => '1',
		13518 => '1',
		13519 => '1',
		13520 => '1',
		13521 => '1',
		13522 => '0',
		13523 => '0',
		13524 => '0',
		13525 => '0',
		13526 => '0',
		13527 => '1',
		13528 => '1',
		13529 => '1',
		13530 => '0',
		13531 => '0',
		13532 => '0',
		13533 => '0',
		13534 => '0',
		13535 => '0',
		13536 => '0',
		13537 => '0',
		13538 => '0',
		13539 => '0',
		13540 => '0',
		13541 => '0',
		13542 => '0',
		13543 => '0',
		13544 => '0',
		13545 => '0',
		13546 => '0',
		13547 => '0',
		13548 => '0',
		13549 => '0',
		13550 => '0',
		13551 => '0',
		13552 => '0',
		13553 => '0',
		13554 => '0',
		13555 => '0',
		13556 => '0',
		13557 => '0',
		13558 => '0',
		13559 => '0',
		13568 => '0',
		13569 => '0',
		13570 => '0',
		13571 => '0',
		13572 => '0',
		13573 => '0',
		13574 => '0',
		13575 => '0',
		13576 => '0',
		13577 => '0',
		13578 => '0',
		13579 => '0',
		13580 => '0',
		13581 => '0',
		13582 => '0',
		13583 => '0',
		13584 => '0',
		13585 => '0',
		13586 => '0',
		13587 => '0',
		13588 => '0',
		13589 => '0',
		13590 => '0',
		13591 => '0',
		13592 => '0',
		13593 => '0',
		13594 => '0',
		13595 => '0',
		13596 => '0',
		13597 => '0',
		13598 => '0',
		13599 => '0',
		13600 => '0',
		13601 => '0',
		13602 => '0',
		13603 => '0',
		13604 => '0',
		13605 => '0',
		13606 => '0',
		13607 => '0',
		13608 => '1',
		13609 => '0',
		13610 => '0',
		13611 => '0',
		13612 => '1',
		13613 => '1',
		13614 => '1',
		13615 => '1',
		13616 => '0',
		13617 => '0',
		13618 => '0',
		13619 => '0',
		13620 => '0',
		13621 => '0',
		13622 => '0',
		13623 => '0',
		13624 => '0',
		13625 => '0',
		13626 => '0',
		13627 => '0',
		13628 => '0',
		13629 => '0',
		13630 => '0',
		13631 => '0',
		13632 => '0',
		13633 => '0',
		13634 => '0',
		13635 => '0',
		13636 => '0',
		13637 => '0',
		13638 => '0',
		13639 => '0',
		13640 => '0',
		13641 => '0',
		13642 => '1',
		13643 => '1',
		13644 => '1',
		13645 => '1',
		13646 => '1',
		13647 => '1',
		13648 => '0',
		13649 => '0',
		13650 => '0',
		13651 => '0',
		13652 => '0',
		13653 => '1',
		13654 => '1',
		13655 => '1',
		13656 => '0',
		13657 => '0',
		13658 => '0',
		13659 => '0',
		13660 => '0',
		13661 => '0',
		13662 => '0',
		13663 => '0',
		13664 => '0',
		13665 => '0',
		13666 => '0',
		13667 => '0',
		13668 => '0',
		13669 => '0',
		13670 => '0',
		13671 => '0',
		13672 => '0',
		13673 => '0',
		13674 => '0',
		13675 => '0',
		13676 => '0',
		13677 => '0',
		13678 => '0',
		13679 => '0',
		13680 => '0',
		13681 => '0',
		13682 => '0',
		13683 => '0',
		13684 => '0',
		13685 => '0',
		13686 => '0',
		13687 => '0',
		13696 => '0',
		13697 => '0',
		13698 => '0',
		13699 => '0',
		13700 => '0',
		13701 => '0',
		13702 => '0',
		13703 => '0',
		13704 => '0',
		13705 => '0',
		13706 => '0',
		13707 => '0',
		13708 => '0',
		13709 => '0',
		13710 => '0',
		13711 => '0',
		13712 => '0',
		13713 => '0',
		13714 => '0',
		13715 => '0',
		13716 => '0',
		13717 => '0',
		13718 => '0',
		13719 => '0',
		13720 => '0',
		13721 => '0',
		13722 => '0',
		13723 => '0',
		13724 => '0',
		13725 => '0',
		13726 => '0',
		13727 => '0',
		13728 => '0',
		13729 => '0',
		13730 => '0',
		13731 => '0',
		13732 => '0',
		13733 => '0',
		13734 => '0',
		13735 => '0',
		13736 => '0',
		13737 => '0',
		13738 => '1',
		13739 => '0',
		13740 => '0',
		13741 => '0',
		13742 => '1',
		13743 => '1',
		13744 => '1',
		13745 => '1',
		13746 => '1',
		13747 => '1',
		13748 => '1',
		13749 => '0',
		13750 => '0',
		13751 => '0',
		13752 => '0',
		13753 => '0',
		13754 => '0',
		13755 => '0',
		13756 => '0',
		13757 => '0',
		13758 => '0',
		13759 => '0',
		13760 => '0',
		13761 => '0',
		13762 => '0',
		13763 => '0',
		13764 => '0',
		13765 => '1',
		13766 => '1',
		13767 => '1',
		13768 => '1',
		13769 => '1',
		13770 => '1',
		13771 => '1',
		13772 => '1',
		13773 => '1',
		13774 => '0',
		13775 => '0',
		13776 => '0',
		13777 => '0',
		13778 => '0',
		13779 => '1',
		13780 => '1',
		13781 => '1',
		13782 => '0',
		13783 => '0',
		13784 => '0',
		13785 => '0',
		13786 => '0',
		13787 => '0',
		13788 => '0',
		13789 => '0',
		13790 => '0',
		13791 => '0',
		13792 => '0',
		13793 => '0',
		13794 => '0',
		13795 => '0',
		13796 => '0',
		13797 => '0',
		13798 => '0',
		13799 => '0',
		13800 => '0',
		13801 => '0',
		13802 => '0',
		13803 => '0',
		13804 => '0',
		13805 => '0',
		13806 => '0',
		13807 => '0',
		13808 => '0',
		13809 => '0',
		13810 => '0',
		13811 => '0',
		13812 => '0',
		13813 => '0',
		13814 => '0',
		13815 => '0',
		13824 => '0',
		13825 => '0',
		13826 => '0',
		13827 => '0',
		13828 => '0',
		13829 => '0',
		13830 => '0',
		13831 => '0',
		13832 => '0',
		13833 => '0',
		13834 => '0',
		13835 => '0',
		13836 => '0',
		13837 => '0',
		13838 => '0',
		13839 => '0',
		13840 => '0',
		13841 => '0',
		13842 => '0',
		13843 => '0',
		13844 => '0',
		13845 => '0',
		13846 => '0',
		13847 => '0',
		13848 => '0',
		13849 => '0',
		13850 => '0',
		13851 => '0',
		13852 => '0',
		13853 => '0',
		13854 => '0',
		13855 => '0',
		13856 => '0',
		13857 => '0',
		13858 => '0',
		13859 => '0',
		13860 => '0',
		13861 => '0',
		13862 => '0',
		13863 => '0',
		13864 => '0',
		13865 => '0',
		13866 => '0',
		13867 => '0',
		13868 => '1',
		13869 => '0',
		13870 => '0',
		13871 => '0',
		13872 => '0',
		13873 => '1',
		13874 => '1',
		13875 => '1',
		13876 => '1',
		13877 => '1',
		13878 => '1',
		13879 => '1',
		13880 => '1',
		13881 => '1',
		13882 => '1',
		13883 => '1',
		13884 => '1',
		13885 => '1',
		13886 => '1',
		13887 => '1',
		13888 => '1',
		13889 => '1',
		13890 => '1',
		13891 => '1',
		13892 => '1',
		13893 => '1',
		13894 => '1',
		13895 => '1',
		13896 => '1',
		13897 => '1',
		13898 => '1',
		13899 => '0',
		13900 => '0',
		13901 => '0',
		13902 => '0',
		13903 => '0',
		13904 => '0',
		13905 => '1',
		13906 => '1',
		13907 => '1',
		13908 => '0',
		13909 => '0',
		13910 => '0',
		13911 => '0',
		13912 => '0',
		13913 => '0',
		13914 => '0',
		13915 => '0',
		13916 => '0',
		13917 => '0',
		13918 => '0',
		13919 => '0',
		13920 => '0',
		13921 => '0',
		13922 => '0',
		13923 => '0',
		13924 => '0',
		13925 => '0',
		13926 => '0',
		13927 => '0',
		13928 => '0',
		13929 => '0',
		13930 => '0',
		13931 => '0',
		13932 => '0',
		13933 => '0',
		13934 => '0',
		13935 => '0',
		13936 => '0',
		13937 => '0',
		13938 => '0',
		13939 => '0',
		13940 => '0',
		13941 => '0',
		13942 => '0',
		13943 => '0',
		13952 => '0',
		13953 => '0',
		13954 => '0',
		13955 => '0',
		13956 => '0',
		13957 => '0',
		13958 => '0',
		13959 => '0',
		13960 => '0',
		13961 => '0',
		13962 => '0',
		13963 => '0',
		13964 => '0',
		13965 => '0',
		13966 => '0',
		13967 => '0',
		13968 => '0',
		13969 => '0',
		13970 => '0',
		13971 => '0',
		13972 => '0',
		13973 => '0',
		13974 => '0',
		13975 => '0',
		13976 => '0',
		13977 => '0',
		13978 => '0',
		13979 => '0',
		13980 => '0',
		13981 => '0',
		13982 => '0',
		13983 => '0',
		13984 => '0',
		13985 => '0',
		13986 => '0',
		13987 => '0',
		13988 => '0',
		13989 => '0',
		13990 => '0',
		13991 => '0',
		13992 => '0',
		13993 => '0',
		13994 => '0',
		13995 => '0',
		13996 => '0',
		13997 => '0',
		13998 => '1',
		13999 => '0',
		14000 => '0',
		14001 => '0',
		14002 => '0',
		14003 => '0',
		14004 => '0',
		14005 => '0',
		14006 => '1',
		14007 => '1',
		14008 => '1',
		14009 => '1',
		14010 => '1',
		14011 => '1',
		14012 => '1',
		14013 => '1',
		14014 => '1',
		14015 => '1',
		14016 => '1',
		14017 => '1',
		14018 => '1',
		14019 => '1',
		14020 => '1',
		14021 => '1',
		14022 => '0',
		14023 => '0',
		14024 => '0',
		14025 => '0',
		14026 => '0',
		14027 => '0',
		14028 => '0',
		14029 => '0',
		14030 => '0',
		14031 => '1',
		14032 => '1',
		14033 => '1',
		14034 => '0',
		14035 => '0',
		14036 => '0',
		14037 => '0',
		14038 => '0',
		14039 => '0',
		14040 => '0',
		14041 => '0',
		14042 => '0',
		14043 => '0',
		14044 => '0',
		14045 => '0',
		14046 => '0',
		14047 => '0',
		14048 => '0',
		14049 => '0',
		14050 => '0',
		14051 => '0',
		14052 => '0',
		14053 => '0',
		14054 => '0',
		14055 => '0',
		14056 => '0',
		14057 => '0',
		14058 => '0',
		14059 => '0',
		14060 => '0',
		14061 => '0',
		14062 => '0',
		14063 => '0',
		14064 => '0',
		14065 => '0',
		14066 => '0',
		14067 => '0',
		14068 => '0',
		14069 => '0',
		14070 => '0',
		14071 => '0',
		14080 => '0',
		14081 => '0',
		14082 => '0',
		14083 => '0',
		14084 => '0',
		14085 => '0',
		14086 => '0',
		14087 => '0',
		14088 => '0',
		14089 => '0',
		14090 => '0',
		14091 => '0',
		14092 => '0',
		14093 => '0',
		14094 => '0',
		14095 => '0',
		14096 => '0',
		14097 => '0',
		14098 => '0',
		14099 => '0',
		14100 => '0',
		14101 => '0',
		14102 => '0',
		14103 => '0',
		14104 => '0',
		14105 => '0',
		14106 => '0',
		14107 => '0',
		14108 => '0',
		14109 => '0',
		14110 => '0',
		14111 => '0',
		14112 => '0',
		14113 => '0',
		14114 => '0',
		14115 => '0',
		14116 => '0',
		14117 => '0',
		14118 => '0',
		14119 => '0',
		14120 => '0',
		14121 => '0',
		14122 => '0',
		14123 => '0',
		14124 => '0',
		14125 => '0',
		14126 => '0',
		14127 => '0',
		14128 => '1',
		14129 => '1',
		14130 => '0',
		14131 => '0',
		14132 => '0',
		14133 => '0',
		14134 => '0',
		14135 => '0',
		14136 => '0',
		14137 => '0',
		14138 => '0',
		14139 => '0',
		14140 => '0',
		14141 => '0',
		14142 => '0',
		14143 => '0',
		14144 => '0',
		14145 => '0',
		14146 => '0',
		14147 => '0',
		14148 => '0',
		14149 => '0',
		14150 => '0',
		14151 => '0',
		14152 => '0',
		14153 => '0',
		14154 => '0',
		14155 => '0',
		14156 => '1',
		14157 => '1',
		14158 => '1',
		14159 => '1',
		14160 => '0',
		14161 => '0',
		14162 => '0',
		14163 => '0',
		14164 => '0',
		14165 => '0',
		14166 => '0',
		14167 => '0',
		14168 => '0',
		14169 => '0',
		14170 => '0',
		14171 => '0',
		14172 => '0',
		14173 => '0',
		14174 => '0',
		14175 => '0',
		14176 => '0',
		14177 => '0',
		14178 => '0',
		14179 => '0',
		14180 => '0',
		14181 => '0',
		14182 => '0',
		14183 => '0',
		14184 => '0',
		14185 => '0',
		14186 => '0',
		14187 => '0',
		14188 => '0',
		14189 => '0',
		14190 => '0',
		14191 => '0',
		14192 => '0',
		14193 => '0',
		14194 => '0',
		14195 => '0',
		14196 => '0',
		14197 => '0',
		14198 => '0',
		14199 => '0',
		14208 => '0',
		14209 => '0',
		14210 => '0',
		14211 => '0',
		14212 => '0',
		14213 => '0',
		14214 => '0',
		14215 => '0',
		14216 => '0',
		14217 => '0',
		14218 => '0',
		14219 => '0',
		14220 => '0',
		14221 => '0',
		14222 => '0',
		14223 => '0',
		14224 => '0',
		14225 => '0',
		14226 => '0',
		14227 => '0',
		14228 => '0',
		14229 => '0',
		14230 => '0',
		14231 => '0',
		14232 => '0',
		14233 => '0',
		14234 => '0',
		14235 => '0',
		14236 => '0',
		14237 => '0',
		14238 => '0',
		14239 => '0',
		14240 => '0',
		14241 => '0',
		14242 => '0',
		14243 => '0',
		14244 => '0',
		14245 => '0',
		14246 => '0',
		14247 => '0',
		14248 => '0',
		14249 => '0',
		14250 => '0',
		14251 => '0',
		14252 => '0',
		14253 => '0',
		14254 => '0',
		14255 => '0',
		14256 => '0',
		14257 => '0',
		14258 => '0',
		14259 => '1',
		14260 => '1',
		14261 => '1',
		14262 => '1',
		14263 => '0',
		14264 => '0',
		14265 => '0',
		14266 => '0',
		14267 => '0',
		14268 => '0',
		14269 => '0',
		14270 => '0',
		14271 => '0',
		14272 => '0',
		14273 => '0',
		14274 => '0',
		14275 => '0',
		14276 => '0',
		14277 => '0',
		14278 => '0',
		14279 => '1',
		14280 => '1',
		14281 => '1',
		14282 => '1',
		14283 => '1',
		14284 => '1',
		14285 => '0',
		14286 => '0',
		14287 => '0',
		14288 => '0',
		14289 => '0',
		14290 => '0',
		14291 => '0',
		14292 => '0',
		14293 => '0',
		14294 => '0',
		14295 => '0',
		14296 => '0',
		14297 => '0',
		14298 => '0',
		14299 => '0',
		14300 => '0',
		14301 => '0',
		14302 => '0',
		14303 => '0',
		14304 => '0',
		14305 => '0',
		14306 => '0',
		14307 => '0',
		14308 => '0',
		14309 => '0',
		14310 => '0',
		14311 => '0',
		14312 => '0',
		14313 => '0',
		14314 => '0',
		14315 => '0',
		14316 => '0',
		14317 => '0',
		14318 => '0',
		14319 => '0',
		14320 => '0',
		14321 => '0',
		14322 => '0',
		14323 => '0',
		14324 => '0',
		14325 => '0',
		14326 => '0',
		14327 => '0',
		14336 => '0',
		14337 => '0',
		14338 => '0',
		14339 => '0',
		14340 => '0',
		14341 => '0',
		14342 => '0',
		14343 => '0',
		14344 => '0',
		14345 => '0',
		14346 => '0',
		14347 => '0',
		14348 => '0',
		14349 => '0',
		14350 => '0',
		14351 => '0',
		14352 => '0',
		14353 => '0',
		14354 => '0',
		14355 => '0',
		14356 => '0',
		14357 => '0',
		14358 => '0',
		14359 => '0',
		14360 => '0',
		14361 => '0',
		14362 => '0',
		14363 => '0',
		14364 => '0',
		14365 => '0',
		14366 => '0',
		14367 => '0',
		14368 => '0',
		14369 => '0',
		14370 => '0',
		14371 => '0',
		14372 => '0',
		14373 => '0',
		14374 => '0',
		14375 => '0',
		14376 => '0',
		14377 => '0',
		14378 => '0',
		14379 => '0',
		14380 => '0',
		14381 => '0',
		14382 => '0',
		14383 => '0',
		14384 => '0',
		14385 => '0',
		14386 => '0',
		14387 => '0',
		14388 => '0',
		14389 => '0',
		14390 => '0',
		14391 => '0',
		14392 => '1',
		14393 => '1',
		14394 => '1',
		14395 => '1',
		14396 => '1',
		14397 => '1',
		14398 => '1',
		14399 => '1',
		14400 => '1',
		14401 => '1',
		14402 => '1',
		14403 => '1',
		14404 => '1',
		14405 => '1',
		14406 => '1',
		14407 => '1',
		14408 => '0',
		14409 => '0',
		14410 => '0',
		14411 => '0',
		14412 => '0',
		14413 => '0',
		14414 => '0',
		14415 => '0',
		14416 => '0',
		14417 => '0',
		14418 => '0',
		14419 => '0',
		14420 => '0',
		14421 => '0',
		14422 => '0',
		14423 => '0',
		14424 => '0',
		14425 => '0',
		14426 => '0',
		14427 => '0',
		14428 => '0',
		14429 => '0',
		14430 => '0',
		14431 => '0',
		14432 => '0',
		14433 => '0',
		14434 => '0',
		14435 => '0',
		14436 => '0',
		14437 => '0',
		14438 => '0',
		14439 => '0',
		14440 => '0',
		14441 => '0',
		14442 => '0',
		14443 => '0',
		14444 => '0',
		14445 => '0',
		14446 => '0',
		14447 => '0',
		14448 => '0',
		14449 => '0',
		14450 => '0',
		14451 => '0',
		14452 => '0',
		14453 => '0',
		14454 => '0',
		14455 => '0',
		14464 => '0',
		14465 => '0',
		14466 => '0',
		14467 => '0',
		14468 => '0',
		14469 => '0',
		14470 => '0',
		14471 => '0',
		14472 => '0',
		14473 => '0',
		14474 => '0',
		14475 => '0',
		14476 => '0',
		14477 => '0',
		14478 => '0',
		14479 => '0',
		14480 => '0',
		14481 => '0',
		14482 => '0',
		14483 => '0',
		14484 => '0',
		14485 => '0',
		14486 => '0',
		14487 => '0',
		14488 => '0',
		14489 => '0',
		14490 => '0',
		14491 => '0',
		14492 => '0',
		14493 => '0',
		14494 => '0',
		14495 => '0',
		14496 => '0',
		14497 => '0',
		14498 => '0',
		14499 => '0',
		14500 => '0',
		14501 => '0',
		14502 => '0',
		14503 => '0',
		14504 => '0',
		14505 => '0',
		14506 => '0',
		14507 => '0',
		14508 => '0',
		14509 => '0',
		14510 => '0',
		14511 => '0',
		14512 => '0',
		14513 => '0',
		14514 => '0',
		14515 => '0',
		14516 => '0',
		14517 => '0',
		14518 => '0',
		14519 => '0',
		14520 => '0',
		14521 => '0',
		14522 => '0',
		14523 => '0',
		14524 => '0',
		14525 => '0',
		14526 => '0',
		14527 => '0',
		14528 => '0',
		14529 => '0',
		14530 => '0',
		14531 => '0',
		14532 => '0',
		14533 => '0',
		14534 => '0',
		14535 => '0',
		14536 => '0',
		14537 => '0',
		14538 => '0',
		14539 => '0',
		14540 => '0',
		14541 => '0',
		14542 => '0',
		14543 => '0',
		14544 => '0',
		14545 => '0',
		14546 => '0',
		14547 => '0',
		14548 => '0',
		14549 => '0',
		14550 => '0',
		14551 => '0',
		14552 => '0',
		14553 => '0',
		14554 => '0',
		14555 => '0',
		14556 => '0',
		14557 => '0',
		14558 => '0',
		14559 => '0',
		14560 => '0',
		14561 => '0',
		14562 => '0',
		14563 => '0',
		14564 => '0',
		14565 => '0',
		14566 => '0',
		14567 => '0',
		14568 => '0',
		14569 => '0',
		14570 => '0',
		14571 => '0',
		14572 => '0',
		14573 => '0',
		14574 => '0',
		14575 => '0',
		14576 => '0',
		14577 => '0',
		14578 => '0',
		14579 => '0',
		14580 => '0',
		14581 => '0',
		14582 => '0',
		14583 => '0',
		14592 => '0',
		14593 => '0',
		14594 => '0',
		14595 => '0',
		14596 => '0',
		14597 => '0',
		14598 => '0',
		14599 => '0',
		14600 => '0',
		14601 => '0',
		14602 => '0',
		14603 => '0',
		14604 => '0',
		14605 => '0',
		14606 => '0',
		14607 => '0',
		14608 => '0',
		14609 => '0',
		14610 => '0',
		14611 => '0',
		14612 => '0',
		14613 => '0',
		14614 => '0',
		14615 => '0',
		14616 => '0',
		14617 => '0',
		14618 => '0',
		14619 => '0',
		14620 => '0',
		14621 => '0',
		14622 => '0',
		14623 => '0',
		14624 => '0',
		14625 => '0',
		14626 => '0',
		14627 => '0',
		14628 => '0',
		14629 => '0',
		14630 => '0',
		14631 => '0',
		14632 => '0',
		14633 => '0',
		14634 => '0',
		14635 => '0',
		14636 => '0',
		14637 => '0',
		14638 => '0',
		14639 => '0',
		14640 => '0',
		14641 => '0',
		14642 => '0',
		14643 => '0',
		14644 => '0',
		14645 => '0',
		14646 => '0',
		14647 => '0',
		14648 => '0',
		14649 => '0',
		14650 => '0',
		14651 => '0',
		14652 => '0',
		14653 => '0',
		14654 => '0',
		14655 => '0',
		14656 => '0',
		14657 => '0',
		14658 => '0',
		14659 => '0',
		14660 => '0',
		14661 => '0',
		14662 => '0',
		14663 => '0',
		14664 => '0',
		14665 => '0',
		14666 => '0',
		14667 => '0',
		14668 => '0',
		14669 => '0',
		14670 => '0',
		14671 => '0',
		14672 => '0',
		14673 => '0',
		14674 => '0',
		14675 => '0',
		14676 => '0',
		14677 => '0',
		14678 => '0',
		14679 => '0',
		14680 => '0',
		14681 => '0',
		14682 => '0',
		14683 => '0',
		14684 => '0',
		14685 => '0',
		14686 => '0',
		14687 => '0',
		14688 => '0',
		14689 => '0',
		14690 => '0',
		14691 => '0',
		14692 => '0',
		14693 => '0',
		14694 => '0',
		14695 => '0',
		14696 => '0',
		14697 => '0',
		14698 => '0',
		14699 => '0',
		14700 => '0',
		14701 => '0',
		14702 => '0',
		14703 => '0',
		14704 => '0',
		14705 => '0',
		14706 => '0',
		14707 => '0',
		14708 => '0',
		14709 => '0',
		14710 => '0',
		14711 => '0',
		14720 => '0',
		14721 => '0',
		14722 => '0',
		14723 => '0',
		14724 => '0',
		14725 => '0',
		14726 => '0',
		14727 => '0',
		14728 => '0',
		14729 => '0',
		14730 => '0',
		14731 => '0',
		14732 => '0',
		14733 => '0',
		14734 => '0',
		14735 => '0',
		14736 => '0',
		14737 => '0',
		14738 => '0',
		14739 => '0',
		14740 => '0',
		14741 => '0',
		14742 => '0',
		14743 => '0',
		14744 => '0',
		14745 => '0',
		14746 => '0',
		14747 => '0',
		14748 => '0',
		14749 => '0',
		14750 => '0',
		14751 => '0',
		14752 => '0',
		14753 => '0',
		14754 => '0',
		14755 => '0',
		14756 => '0',
		14757 => '0',
		14758 => '0',
		14759 => '0',
		14760 => '0',
		14761 => '0',
		14762 => '0',
		14763 => '0',
		14764 => '0',
		14765 => '0',
		14766 => '0',
		14767 => '0',
		14768 => '0',
		14769 => '0',
		14770 => '0',
		14771 => '0',
		14772 => '0',
		14773 => '0',
		14774 => '0',
		14775 => '0',
		14776 => '0',
		14777 => '0',
		14778 => '0',
		14779 => '0',
		14780 => '0',
		14781 => '0',
		14782 => '0',
		14783 => '0',
		14784 => '0',
		14785 => '0',
		14786 => '0',
		14787 => '0',
		14788 => '0',
		14789 => '0',
		14790 => '0',
		14791 => '0',
		14792 => '0',
		14793 => '0',
		14794 => '0',
		14795 => '0',
		14796 => '0',
		14797 => '0',
		14798 => '0',
		14799 => '0',
		14800 => '0',
		14801 => '0',
		14802 => '0',
		14803 => '0',
		14804 => '0',
		14805 => '0',
		14806 => '0',
		14807 => '0',
		14808 => '0',
		14809 => '0',
		14810 => '0',
		14811 => '0',
		14812 => '0',
		14813 => '0',
		14814 => '0',
		14815 => '0',
		14816 => '0',
		14817 => '0',
		14818 => '0',
		14819 => '0',
		14820 => '0',
		14821 => '0',
		14822 => '0',
		14823 => '0',
		14824 => '0',
		14825 => '0',
		14826 => '0',
		14827 => '0',
		14828 => '0',
		14829 => '0',
		14830 => '0',
		14831 => '0',
		14832 => '0',
		14833 => '0',
		14834 => '0',
		14835 => '0',
		14836 => '0',
		14837 => '0',
		14838 => '0',
		14839 => '0',
		14848 => '0',
		14849 => '0',
		14850 => '0',
		14851 => '0',
		14852 => '0',
		14853 => '0',
		14854 => '0',
		14855 => '0',
		14856 => '0',
		14857 => '0',
		14858 => '0',
		14859 => '0',
		14860 => '0',
		14861 => '0',
		14862 => '0',
		14863 => '0',
		14864 => '0',
		14865 => '0',
		14866 => '0',
		14867 => '0',
		14868 => '0',
		14869 => '0',
		14870 => '0',
		14871 => '0',
		14872 => '0',
		14873 => '0',
		14874 => '0',
		14875 => '0',
		14876 => '0',
		14877 => '0',
		14878 => '0',
		14879 => '0',
		14880 => '0',
		14881 => '0',
		14882 => '0',
		14883 => '0',
		14884 => '0',
		14885 => '0',
		14886 => '0',
		14887 => '0',
		14888 => '0',
		14889 => '0',
		14890 => '0',
		14891 => '0',
		14892 => '0',
		14893 => '0',
		14894 => '0',
		14895 => '0',
		14896 => '0',
		14897 => '0',
		14898 => '0',
		14899 => '0',
		14900 => '0',
		14901 => '0',
		14902 => '0',
		14903 => '0',
		14904 => '0',
		14905 => '0',
		14906 => '0',
		14907 => '0',
		14908 => '0',
		14909 => '0',
		14910 => '0',
		14911 => '0',
		14912 => '0',
		14913 => '0',
		14914 => '0',
		14915 => '0',
		14916 => '0',
		14917 => '0',
		14918 => '0',
		14919 => '0',
		14920 => '0',
		14921 => '0',
		14922 => '0',
		14923 => '0',
		14924 => '0',
		14925 => '0',
		14926 => '0',
		14927 => '0',
		14928 => '0',
		14929 => '0',
		14930 => '0',
		14931 => '0',
		14932 => '0',
		14933 => '0',
		14934 => '0',
		14935 => '0',
		14936 => '0',
		14937 => '0',
		14938 => '0',
		14939 => '0',
		14940 => '0',
		14941 => '0',
		14942 => '0',
		14943 => '0',
		14944 => '0',
		14945 => '0',
		14946 => '0',
		14947 => '0',
		14948 => '0',
		14949 => '0',
		14950 => '0',
		14951 => '0',
		14952 => '0',
		14953 => '0',
		14954 => '0',
		14955 => '0',
		14956 => '0',
		14957 => '0',
		14958 => '0',
		14959 => '0',
		14960 => '0',
		14961 => '0',
		14962 => '0',
		14963 => '0',
		14964 => '0',
		14965 => '0',
		14966 => '0',
		14967 => '0',
		14976 => '0',
		14977 => '0',
		14978 => '0',
		14979 => '0',
		14980 => '0',
		14981 => '0',
		14982 => '0',
		14983 => '0',
		14984 => '0',
		14985 => '0',
		14986 => '0',
		14987 => '0',
		14988 => '0',
		14989 => '0',
		14990 => '0',
		14991 => '0',
		14992 => '0',
		14993 => '0',
		14994 => '0',
		14995 => '0',
		14996 => '0',
		14997 => '0',
		14998 => '0',
		14999 => '0',
		15000 => '0',
		15001 => '0',
		15002 => '0',
		15003 => '0',
		15004 => '0',
		15005 => '0',
		15006 => '0',
		15007 => '0',
		15008 => '0',
		15009 => '0',
		15010 => '0',
		15011 => '0',
		15012 => '0',
		15013 => '0',
		15014 => '0',
		15015 => '0',
		15016 => '0',
		15017 => '0',
		15018 => '0',
		15019 => '0',
		15020 => '0',
		15021 => '0',
		15022 => '0',
		15023 => '0',
		15024 => '0',
		15025 => '0',
		15026 => '0',
		15027 => '0',
		15028 => '0',
		15029 => '0',
		15030 => '0',
		15031 => '0',
		15032 => '0',
		15033 => '0',
		15034 => '0',
		15035 => '0',
		15036 => '0',
		15037 => '0',
		15038 => '0',
		15039 => '0',
		15040 => '0',
		15041 => '0',
		15042 => '0',
		15043 => '0',
		15044 => '0',
		15045 => '0',
		15046 => '0',
		15047 => '0',
		15048 => '0',
		15049 => '0',
		15050 => '0',
		15051 => '0',
		15052 => '0',
		15053 => '0',
		15054 => '0',
		15055 => '0',
		15056 => '0',
		15057 => '0',
		15058 => '0',
		15059 => '0',
		15060 => '0',
		15061 => '0',
		15062 => '0',
		15063 => '0',
		15064 => '0',
		15065 => '0',
		15066 => '0',
		15067 => '0',
		15068 => '0',
		15069 => '0',
		15070 => '0',
		15071 => '0',
		15072 => '0',
		15073 => '0',
		15074 => '0',
		15075 => '0',
		15076 => '0',
		15077 => '0',
		15078 => '0',
		15079 => '0',
		15080 => '0',
		15081 => '0',
		15082 => '0',
		15083 => '0',
		15084 => '0',
		15085 => '0',
		15086 => '0',
		15087 => '0',
		15088 => '0',
		15089 => '0',
		15090 => '0',
		15091 => '0',
		15092 => '0',
		15093 => '0',
		15094 => '0',
		15095 => '0',
		15104 => '0',
		15105 => '0',
		15106 => '0',
		15107 => '0',
		15108 => '0',
		15109 => '0',
		15110 => '0',
		15111 => '0',
		15112 => '0',
		15113 => '0',
		15114 => '0',
		15115 => '0',
		15116 => '0',
		15117 => '0',
		15118 => '0',
		15119 => '0',
		15120 => '0',
		15121 => '0',
		15122 => '0',
		15123 => '0',
		15124 => '0',
		15125 => '0',
		15126 => '0',
		15127 => '0',
		15128 => '0',
		15129 => '0',
		15130 => '0',
		15131 => '0',
		15132 => '0',
		15133 => '0',
		15134 => '0',
		15135 => '0',
		15136 => '0',
		15137 => '0',
		15138 => '0',
		15139 => '0',
		15140 => '0',
		15141 => '0',
		15142 => '0',
		15143 => '0',
		15144 => '0',
		15145 => '0',
		15146 => '0',
		15147 => '0',
		15148 => '0',
		15149 => '0',
		15150 => '0',
		15151 => '0',
		15152 => '0',
		15153 => '0',
		15154 => '0',
		15155 => '0',
		15156 => '0',
		15157 => '0',
		15158 => '0',
		15159 => '0',
		15160 => '0',
		15161 => '0',
		15162 => '0',
		15163 => '0',
		15164 => '0',
		15165 => '0',
		15166 => '0',
		15167 => '0',
		15168 => '0',
		15169 => '0',
		15170 => '0',
		15171 => '0',
		15172 => '0',
		15173 => '0',
		15174 => '0',
		15175 => '0',
		15176 => '0',
		15177 => '0',
		15178 => '0',
		15179 => '0',
		15180 => '0',
		15181 => '0',
		15182 => '0',
		15183 => '0',
		15184 => '0',
		15185 => '0',
		15186 => '0',
		15187 => '0',
		15188 => '0',
		15189 => '0',
		15190 => '0',
		15191 => '0',
		15192 => '0',
		15193 => '0',
		15194 => '0',
		15195 => '0',
		15196 => '0',
		15197 => '0',
		15198 => '0',
		15199 => '0',
		15200 => '0',
		15201 => '0',
		15202 => '0',
		15203 => '0',
		15204 => '0',
		15205 => '0',
		15206 => '0',
		15207 => '0',
		15208 => '0',
		15209 => '0',
		15210 => '0',
		15211 => '0',
		15212 => '0',
		15213 => '0',
		15214 => '0',
		15215 => '0',
		15216 => '0',
		15217 => '0',
		15218 => '0',
		15219 => '0',
		15220 => '0',
		15221 => '0',
		15222 => '0',
		15223 => '0',
		15232 => '0',
		15233 => '0',
		15234 => '0',
		15235 => '0',
		15236 => '0',
		15237 => '0',
		15238 => '0',
		15239 => '0',
		15240 => '0',
		15241 => '0',
		15242 => '0',
		15243 => '0',
		15244 => '0',
		15245 => '0',
		15246 => '0',
		15247 => '0',
		15248 => '0',
		15249 => '0',
		15250 => '0',
		15251 => '0',
		15252 => '0',
		15253 => '0',
		15254 => '0',
		15255 => '0',
		15256 => '0',
		15257 => '0',
		15258 => '0',
		15259 => '0',
		15260 => '0',
		15261 => '0',
		15262 => '0',
		15263 => '0',
		15264 => '0',
		15265 => '0',
		15266 => '0',
		15267 => '0',
		15268 => '0',
		15269 => '0',
		15270 => '0',
		15271 => '0',
		15272 => '0',
		15273 => '0',
		15274 => '0',
		15275 => '0',
		15276 => '0',
		15277 => '0',
		15278 => '0',
		15279 => '0',
		15280 => '0',
		15281 => '0',
		15282 => '0',
		15283 => '0',
		15284 => '0',
		15285 => '0',
		15286 => '0',
		15287 => '0',
		15288 => '0',
		15289 => '0',
		15290 => '0',
		15291 => '0',
		15292 => '0',
		15293 => '0',
		15294 => '0',
		15295 => '0',
		15296 => '0',
		15297 => '0',
		15298 => '0',
		15299 => '0',
		15300 => '0',
		15301 => '0',
		15302 => '0',
		15303 => '0',
		15304 => '0',
		15305 => '0',
		15306 => '0',
		15307 => '0',
		15308 => '0',
		15309 => '0',
		15310 => '0',
		15311 => '0',
		15312 => '0',
		15313 => '0',
		15314 => '0',
		15315 => '0',
		15316 => '0',
		15317 => '0',
		15318 => '0',
		15319 => '0',
		15320 => '0',
		15321 => '0',
		15322 => '0',
		15323 => '0',
		15324 => '0',
		15325 => '0',
		15326 => '0',
		15327 => '0',
		15328 => '0',
		15329 => '0',
		15330 => '0',
		15331 => '0',
		15332 => '0',
		15333 => '0',
		15334 => '0',
		15335 => '0',
		15336 => '0',
		15337 => '0',
		15338 => '0',
		15339 => '0',
		15340 => '0',
		15341 => '0',
		15342 => '0',
		15343 => '0',
		15344 => '0',
		15345 => '0',
		15346 => '0',
		15347 => '0',
		15348 => '0',
		15349 => '0',
		15350 => '0',
		15351 => '0',

	others => '0'
);

begin
	
	-- process ROM
	process (CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (EN = '1') then
				DATA <= ROM(to_integer(unsigned(ADDR)));
			end if;
		end if;
	end process;
	
end Behavioral;

